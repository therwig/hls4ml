
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This doocument may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_vld_v1 (idat, ivld, dat, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             ivld;
  input  [width-1:0] dat;
  input              vld;

  wire   [width-1:0] idat;
  wire               ivld;

  assign idat = dat;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_vld_v1 (dat, vld, idat, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             vld;
  input  [width-1:0] idat;
  input              ivld;

  wire   [width-1:0] dat;
  wire               vld;

  assign dat = idat;
  assign vld = ivld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Mar  8 19:20:36 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module econ_4x4_d10_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for econ_4x4_d10_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : econ_4x4_d10_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_staller
// ------------------------------------------------------------------


module econ_4x4_d10_core_staller (
  clk, rst, core_wen, core_wten, input_1_rsci_wen_comp, w2_rsci_wen_comp, b2_rsci_wen_comp,
      w4_rsci_wen_comp, b4_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_1_rsci_wen_comp;
  input w2_rsci_wen_comp;
  input b2_rsci_wen_comp;
  input w4_rsci_wen_comp;
  input b4_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_1_rsci_wen_comp & w2_rsci_wen_comp & b2_rsci_wen_comp &
      w4_rsci_wen_comp & b4_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl (
  core_wten, b4_rsc_triosy_obj_iswt0, b4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;
  output b4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b4_rsc_triosy_obj_ld_core_sct = b4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl (
  core_wten, w4_rsc_triosy_obj_iswt0, w4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;
  output w4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w4_rsc_triosy_obj_ld_core_sct = w4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl (
  core_wten, b2_rsc_triosy_obj_iswt0, b2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;
  output b2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b2_rsc_triosy_obj_ld_core_sct = b2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl (
  core_wten, w2_rsc_triosy_obj_iswt0, w2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;
  output w2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w2_rsc_triosy_obj_ld_core_sct = w2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_out_1_rsc_triosy_obj_iswt0, const_size_out_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;
  output const_size_out_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsc_triosy_obj_ld_core_sct = const_size_out_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_in_1_rsc_triosy_obj_iswt0, const_size_in_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;
  output const_size_in_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsc_triosy_obj_ld_core_sct = const_size_in_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
    (
  core_wten, layer5_out_rsc_triosy_obj_iswt0, layer5_out_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;
  output layer5_out_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsc_triosy_obj_ld_core_sct = layer5_out_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl (
  core_wten, input_1_rsc_triosy_obj_iswt0, input_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;
  output input_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsc_triosy_obj_ld_core_sct = input_1_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsci (
  b4_rsc_dat, b4_rsc_vld, b4_rsci_oswt, b4_rsci_wen_comp, b4_rsci_idat_mxwt
);
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [79:0] b4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b4_rsci_ivld;
  wire [79:0] b4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd8),
  .width(32'sd80)) b4_rsci (
      .vld(b4_rsc_vld),
      .dat(b4_rsc_dat),
      .ivld(b4_rsci_ivld),
      .idat(b4_rsci_idat)
    );
  assign b4_rsci_idat_mxwt = b4_rsci_idat;
  assign b4_rsci_wen_comp = (~ b4_rsci_oswt) | b4_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsci (
  w4_rsc_dat, w4_rsc_vld, w4_rsci_oswt, w4_rsci_wen_comp, w4_rsci_idat_mxwt
);
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [10239:0] w4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w4_rsci_ivld;
  wire [10239:0] w4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd7),
  .width(32'sd10240)) w4_rsci (
      .vld(w4_rsc_vld),
      .dat(w4_rsc_dat),
      .ivld(w4_rsci_ivld),
      .idat(w4_rsci_idat)
    );
  assign w4_rsci_idat_mxwt = w4_rsci_idat;
  assign w4_rsci_wen_comp = (~ w4_rsci_oswt) | w4_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsci (
  b2_rsc_dat, b2_rsc_vld, b2_rsci_oswt, b2_rsci_wen_comp, b2_rsci_idat_mxwt
);
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [63:0] b2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b2_rsci_ivld;
  wire [63:0] b2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd6),
  .width(32'sd64)) b2_rsci (
      .vld(b2_rsc_vld),
      .dat(b2_rsc_dat),
      .ivld(b2_rsci_ivld),
      .idat(b2_rsci_idat)
    );
  assign b2_rsci_idat_mxwt = b2_rsci_idat;
  assign b2_rsci_wen_comp = (~ b2_rsci_oswt) | b2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsci (
  w2_rsc_dat, w2_rsc_vld, w2_rsci_oswt, w2_rsci_wen_comp, w2_rsci_idat_mxwt
);
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [1727:0] w2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w2_rsci_ivld;
  wire [1727:0] w2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd5),
  .width(32'sd1728)) w2_rsci (
      .vld(w2_rsc_vld),
      .dat(w2_rsc_dat),
      .ivld(w2_rsci_ivld),
      .idat(w2_rsci_idat)
    );
  assign w2_rsci_idat_mxwt = w2_rsci_idat;
  assign w2_rsci_wen_comp = (~ w2_rsci_oswt) | w2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wten, const_size_out_1_rsci_iswt0, const_size_out_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_out_1_rsci_iswt0;
  output const_size_out_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wten, const_size_in_1_rsci_iswt0, const_size_in_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_in_1_rsci_iswt0;
  output const_size_in_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl (
  core_wten, layer5_out_rsci_iswt0, layer5_out_rsci_ivld_core_sct
);
  input core_wten;
  input layer5_out_rsci_iswt0;
  output layer5_out_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_ivld_core_sct = layer5_out_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsci (
  input_1_rsc_dat, input_1_rsc_vld, input_1_rsci_oswt, input_1_rsci_wen_comp, input_1_rsci_idat_mxwt
);
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [1055:0] input_1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_1_rsci_ivld;
  wire [1055:0] input_1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd1),
  .width(32'sd1056)) input_1_rsci (
      .vld(input_1_rsc_vld),
      .dat(input_1_rsc_dat),
      .ivld(input_1_rsci_ivld),
      .idat(input_1_rsci_idat)
    );
  assign input_1_rsci_idat_mxwt = input_1_rsci_idat;
  assign input_1_rsci_wen_comp = (~ input_1_rsci_oswt) | input_1_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj (
  b4_rsc_triosy_lz, core_wten, b4_rsc_triosy_obj_iswt0
);
  output b4_rsc_triosy_lz;
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b4_rsc_triosy_obj (
      .ld(b4_rsc_triosy_obj_ld_core_sct),
      .lz(b4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(b4_rsc_triosy_obj_iswt0),
      .b4_rsc_triosy_obj_ld_core_sct(b4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj (
  w4_rsc_triosy_lz, core_wten, w4_rsc_triosy_obj_iswt0
);
  output w4_rsc_triosy_lz;
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w4_rsc_triosy_obj (
      .ld(w4_rsc_triosy_obj_ld_core_sct),
      .lz(w4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(w4_rsc_triosy_obj_iswt0),
      .w4_rsc_triosy_obj_ld_core_sct(w4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj (
  b2_rsc_triosy_lz, core_wten, b2_rsc_triosy_obj_iswt0
);
  output b2_rsc_triosy_lz;
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b2_rsc_triosy_obj (
      .ld(b2_rsc_triosy_obj_ld_core_sct),
      .lz(b2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(b2_rsc_triosy_obj_iswt0),
      .b2_rsc_triosy_obj_ld_core_sct(b2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj (
  w2_rsc_triosy_lz, core_wten, w2_rsc_triosy_obj_iswt0
);
  output w2_rsc_triosy_lz;
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w2_rsc_triosy_obj (
      .ld(w2_rsc_triosy_obj_ld_core_sct),
      .lz(w2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(w2_rsc_triosy_obj_iswt0),
      .w2_rsc_triosy_obj_ld_core_sct(w2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj (
  const_size_out_1_rsc_triosy_lz, core_wten, const_size_out_1_rsc_triosy_obj_iswt0
);
  output const_size_out_1_rsc_triosy_lz;
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_out_1_rsc_triosy_obj (
      .ld(const_size_out_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_out_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(const_size_out_1_rsc_triosy_obj_iswt0),
      .const_size_out_1_rsc_triosy_obj_ld_core_sct(const_size_out_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj (
  const_size_in_1_rsc_triosy_lz, core_wten, const_size_in_1_rsc_triosy_obj_iswt0
);
  output const_size_in_1_rsc_triosy_lz;
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_in_1_rsc_triosy_obj (
      .ld(const_size_in_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_in_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(const_size_in_1_rsc_triosy_obj_iswt0),
      .const_size_in_1_rsc_triosy_obj_ld_core_sct(const_size_in_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj (
  layer5_out_rsc_triosy_lz, core_wten, layer5_out_rsc_triosy_obj_iswt0
);
  output layer5_out_rsc_triosy_lz;
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire layer5_out_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) layer5_out_rsc_triosy_obj (
      .ld(layer5_out_rsc_triosy_obj_ld_core_sct),
      .lz(layer5_out_rsc_triosy_lz)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(layer5_out_rsc_triosy_obj_iswt0),
      .layer5_out_rsc_triosy_obj_ld_core_sct(layer5_out_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj (
  input_1_rsc_triosy_lz, core_wten, input_1_rsc_triosy_obj_iswt0
);
  output input_1_rsc_triosy_lz;
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire input_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) input_1_rsc_triosy_obj (
      .ld(input_1_rsc_triosy_obj_ld_core_sct),
      .lz(input_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(input_1_rsc_triosy_obj_iswt0),
      .input_1_rsc_triosy_obj_ld_core_sct(input_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci (
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, core_wten, const_size_out_1_rsci_iswt0
);
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input core_wten;
  input const_size_out_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd4),
  .width(32'sd16)) const_size_out_1_rsci (
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000001010),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(const_size_out_1_rsci_iswt0),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci (
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, core_wten, const_size_in_1_rsci_iswt0
);
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input core_wten;
  input const_size_in_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd3),
  .width(32'sd16)) const_size_in_1_rsci (
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000110000),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(const_size_in_1_rsci_iswt0),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci (
  layer5_out_rsc_dat, layer5_out_rsc_vld, core_wten, layer5_out_rsci_iswt0, layer5_out_rsci_idat
);
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input core_wten;
  input layer5_out_rsci_iswt0;
  input [219:0] layer5_out_rsci_idat;


  // Interconnect Declarations
  wire layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [219:0] nl_layer5_out_rsci_idat;
  assign nl_layer5_out_rsci_idat = {1'b0 , (layer5_out_rsci_idat[218:198]) , 1'b0
      , (layer5_out_rsci_idat[196:176]) , 1'b0 , (layer5_out_rsci_idat[174:154])
      , 1'b0 , (layer5_out_rsci_idat[152:132]) , 1'b0 , (layer5_out_rsci_idat[130:110])
      , 1'b0 , (layer5_out_rsci_idat[108:88]) , 1'b0 , (layer5_out_rsci_idat[86:66])
      , 1'b0 , (layer5_out_rsci_idat[64:44]) , 1'b0 , (layer5_out_rsci_idat[42:22])
      , 1'b0 , (layer5_out_rsci_idat[20:0])};
  ccs_out_vld_v1 #(.rscid(32'sd2),
  .width(32'sd220)) layer5_out_rsci (
      .ivld(layer5_out_rsci_ivld_core_sct),
      .idat(nl_layer5_out_rsci_idat[219:0]),
      .vld(layer5_out_rsc_vld),
      .dat(layer5_out_rsc_dat)
    );
  econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer5_out_rsci_iswt0(layer5_out_rsci_iswt0),
      .layer5_out_rsci_ivld_core_sct(layer5_out_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core
// ------------------------------------------------------------------


module econ_4x4_d10_core (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_triosy_lz, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_triosy_lz, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld, w2_rsc_triosy_lz, b2_rsc_dat,
      b2_rsc_vld, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_triosy_lz, b4_rsc_dat,
      b4_rsc_vld, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_triosy_lz;
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_triosy_lz;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_1_rsci_wen_comp;
  wire [1055:0] input_1_rsci_idat_mxwt;
  wire w2_rsci_wen_comp;
  wire [1727:0] w2_rsci_idat_mxwt;
  wire b2_rsci_wen_comp;
  wire [63:0] b2_rsci_idat_mxwt;
  wire w4_rsci_wen_comp;
  wire [10239:0] w4_rsci_idat_mxwt;
  wire b4_rsci_wen_comp;
  wire [79:0] b4_rsci_idat_mxwt;
  reg [20:0] layer5_out_rsci_idat_196_176;
  reg [20:0] layer5_out_rsci_idat_174_154;
  reg [20:0] layer5_out_rsci_idat_152_132;
  reg [20:0] layer5_out_rsci_idat_130_110;
  reg [20:0] layer5_out_rsci_idat_108_88;
  reg [20:0] layer5_out_rsci_idat_86_66;
  reg [20:0] layer5_out_rsci_idat_64_44;
  reg [20:0] layer5_out_rsci_idat_42_22;
  reg [20:0] layer5_out_rsci_idat_20_0;
  reg [20:0] layer5_out_rsci_idat_218_198;
  wire [1:0] fsm_output;
  reg main_stage_0_2;
  wire [21:0] MultLoop_1280_MultLoop_acc_3_ncse_sva_1;
  wire [22:0] nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1;
  wire [21:0] layer4_out_0_sva_1;
  wire [22:0] nl_layer4_out_0_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1;
  wire [21:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1;
  wire [22:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [23:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [24:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1;
  wire [24:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1;
  wire [23:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1;
  wire layer5_out_and_cse;
  reg reg_b4_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse;
  reg [21:0] MultLoop_acc_130_itm_1;
  wire [22:0] nl_MultLoop_acc_130_itm_1;
  reg [21:0] MultLoop_acc_121_itm_1;
  wire [23:0] nl_MultLoop_acc_121_itm_1;
  reg [21:0] MultLoop_acc_120_itm_1;
  wire [23:0] nl_MultLoop_acc_120_itm_1;
  reg [21:0] MultLoop_acc_119_itm_1;
  wire [23:0] nl_MultLoop_acc_119_itm_1;
  reg [21:0] MultLoop_acc_118_itm_1;
  wire [23:0] nl_MultLoop_acc_118_itm_1;
  reg [21:0] MultLoop_acc_117_itm_1;
  wire [23:0] nl_MultLoop_acc_117_itm_1;
  reg [21:0] MultLoop_acc_116_itm_1;
  wire [23:0] nl_MultLoop_acc_116_itm_1;
  reg [21:0] MultLoop_acc_115_itm_1;
  wire [23:0] nl_MultLoop_acc_115_itm_1;
  reg [21:0] MultLoop_acc_114_itm_1;
  wire [23:0] nl_MultLoop_acc_114_itm_1;
  reg [21:0] MultLoop_acc_113_itm_1;
  wire [23:0] nl_MultLoop_acc_113_itm_1;
  reg [21:0] MultLoop_acc_112_itm_1;
  wire [23:0] nl_MultLoop_acc_112_itm_1;
  reg [21:0] MultLoop_acc_111_itm_1;
  wire [23:0] nl_MultLoop_acc_111_itm_1;
  reg [21:0] MultLoop_acc_110_itm_1;
  wire [23:0] nl_MultLoop_acc_110_itm_1;
  reg [21:0] MultLoop_acc_109_itm_1;
  wire [23:0] nl_MultLoop_acc_109_itm_1;
  reg [21:0] MultLoop_acc_108_itm_1;
  wire [23:0] nl_MultLoop_acc_108_itm_1;
  reg [21:0] MultLoop_acc_107_itm_1;
  wire [23:0] nl_MultLoop_acc_107_itm_1;
  reg [21:0] MultLoop_acc_249_itm_1;
  wire [22:0] nl_MultLoop_acc_249_itm_1;
  reg [21:0] MultLoop_acc_248_itm_1;
  wire [23:0] nl_MultLoop_acc_248_itm_1;
  reg [21:0] MultLoop_acc_247_itm_1;
  wire [23:0] nl_MultLoop_acc_247_itm_1;
  reg [21:0] MultLoop_acc_246_itm_1;
  wire [23:0] nl_MultLoop_acc_246_itm_1;
  reg [21:0] MultLoop_acc_245_itm_1;
  wire [23:0] nl_MultLoop_acc_245_itm_1;
  reg [21:0] MultLoop_acc_244_itm_1;
  wire [23:0] nl_MultLoop_acc_244_itm_1;
  reg [21:0] MultLoop_acc_243_itm_1;
  wire [23:0] nl_MultLoop_acc_243_itm_1;
  reg [21:0] MultLoop_acc_242_itm_1;
  wire [23:0] nl_MultLoop_acc_242_itm_1;
  reg [21:0] MultLoop_acc_241_itm_1;
  wire [23:0] nl_MultLoop_acc_241_itm_1;
  reg [21:0] MultLoop_acc_240_itm_1;
  wire [23:0] nl_MultLoop_acc_240_itm_1;
  reg [21:0] MultLoop_acc_239_itm_1;
  wire [23:0] nl_MultLoop_acc_239_itm_1;
  reg [21:0] MultLoop_acc_238_itm_1;
  wire [23:0] nl_MultLoop_acc_238_itm_1;
  reg [21:0] MultLoop_acc_237_itm_1;
  wire [23:0] nl_MultLoop_acc_237_itm_1;
  reg [21:0] MultLoop_acc_236_itm_1;
  wire [23:0] nl_MultLoop_acc_236_itm_1;
  reg [21:0] MultLoop_acc_235_itm_1;
  wire [23:0] nl_MultLoop_acc_235_itm_1;
  reg [21:0] MultLoop_acc_234_itm_1;
  wire [23:0] nl_MultLoop_acc_234_itm_1;
  reg [21:0] MultLoop_acc_376_itm_1;
  wire [22:0] nl_MultLoop_acc_376_itm_1;
  reg [21:0] MultLoop_acc_375_itm_1;
  wire [23:0] nl_MultLoop_acc_375_itm_1;
  reg [21:0] MultLoop_acc_374_itm_1;
  wire [23:0] nl_MultLoop_acc_374_itm_1;
  reg [21:0] MultLoop_acc_373_itm_1;
  wire [23:0] nl_MultLoop_acc_373_itm_1;
  reg [21:0] MultLoop_acc_372_itm_1;
  wire [23:0] nl_MultLoop_acc_372_itm_1;
  reg [21:0] MultLoop_acc_371_itm_1;
  wire [23:0] nl_MultLoop_acc_371_itm_1;
  reg [21:0] MultLoop_acc_370_itm_1;
  wire [23:0] nl_MultLoop_acc_370_itm_1;
  reg [21:0] MultLoop_acc_369_itm_1;
  wire [23:0] nl_MultLoop_acc_369_itm_1;
  reg [21:0] MultLoop_acc_368_itm_1;
  wire [23:0] nl_MultLoop_acc_368_itm_1;
  reg [21:0] MultLoop_acc_367_itm_1;
  wire [23:0] nl_MultLoop_acc_367_itm_1;
  reg [21:0] MultLoop_acc_366_itm_1;
  wire [23:0] nl_MultLoop_acc_366_itm_1;
  reg [21:0] MultLoop_acc_365_itm_1;
  wire [23:0] nl_MultLoop_acc_365_itm_1;
  reg [21:0] MultLoop_acc_364_itm_1;
  wire [23:0] nl_MultLoop_acc_364_itm_1;
  reg [21:0] MultLoop_acc_363_itm_1;
  wire [23:0] nl_MultLoop_acc_363_itm_1;
  reg [21:0] MultLoop_acc_362_itm_1;
  wire [23:0] nl_MultLoop_acc_362_itm_1;
  reg [21:0] MultLoop_acc_361_itm_1;
  wire [23:0] nl_MultLoop_acc_361_itm_1;
  reg [21:0] MultLoop_acc_503_itm_1;
  wire [22:0] nl_MultLoop_acc_503_itm_1;
  reg [21:0] MultLoop_acc_502_itm_1;
  wire [23:0] nl_MultLoop_acc_502_itm_1;
  reg [21:0] MultLoop_acc_501_itm_1;
  wire [23:0] nl_MultLoop_acc_501_itm_1;
  reg [21:0] MultLoop_acc_500_itm_1;
  wire [23:0] nl_MultLoop_acc_500_itm_1;
  reg [21:0] MultLoop_acc_499_itm_1;
  wire [23:0] nl_MultLoop_acc_499_itm_1;
  reg [21:0] MultLoop_acc_498_itm_1;
  wire [23:0] nl_MultLoop_acc_498_itm_1;
  reg [21:0] MultLoop_acc_497_itm_1;
  wire [23:0] nl_MultLoop_acc_497_itm_1;
  reg [21:0] MultLoop_acc_496_itm_1;
  wire [23:0] nl_MultLoop_acc_496_itm_1;
  reg [21:0] MultLoop_acc_495_itm_1;
  wire [23:0] nl_MultLoop_acc_495_itm_1;
  reg [21:0] MultLoop_acc_494_itm_1;
  wire [23:0] nl_MultLoop_acc_494_itm_1;
  reg [21:0] MultLoop_acc_493_itm_1;
  wire [23:0] nl_MultLoop_acc_493_itm_1;
  reg [21:0] MultLoop_acc_492_itm_1;
  wire [23:0] nl_MultLoop_acc_492_itm_1;
  reg [21:0] MultLoop_acc_491_itm_1;
  wire [23:0] nl_MultLoop_acc_491_itm_1;
  reg [21:0] MultLoop_acc_490_itm_1;
  wire [23:0] nl_MultLoop_acc_490_itm_1;
  reg [21:0] MultLoop_acc_489_itm_1;
  wire [23:0] nl_MultLoop_acc_489_itm_1;
  reg [21:0] MultLoop_acc_488_itm_1;
  wire [23:0] nl_MultLoop_acc_488_itm_1;
  reg [21:0] MultLoop_acc_630_itm_1;
  wire [22:0] nl_MultLoop_acc_630_itm_1;
  reg [21:0] MultLoop_acc_629_itm_1;
  wire [23:0] nl_MultLoop_acc_629_itm_1;
  reg [21:0] MultLoop_acc_628_itm_1;
  wire [23:0] nl_MultLoop_acc_628_itm_1;
  reg [21:0] MultLoop_acc_627_itm_1;
  wire [23:0] nl_MultLoop_acc_627_itm_1;
  reg [21:0] MultLoop_acc_626_itm_1;
  wire [23:0] nl_MultLoop_acc_626_itm_1;
  reg [21:0] MultLoop_acc_625_itm_1;
  wire [23:0] nl_MultLoop_acc_625_itm_1;
  reg [21:0] MultLoop_acc_624_itm_1;
  wire [23:0] nl_MultLoop_acc_624_itm_1;
  reg [21:0] MultLoop_acc_623_itm_1;
  wire [23:0] nl_MultLoop_acc_623_itm_1;
  reg [21:0] MultLoop_acc_622_itm_1;
  wire [23:0] nl_MultLoop_acc_622_itm_1;
  reg [21:0] MultLoop_acc_621_itm_1;
  wire [23:0] nl_MultLoop_acc_621_itm_1;
  reg [21:0] MultLoop_acc_620_itm_1;
  wire [23:0] nl_MultLoop_acc_620_itm_1;
  reg [21:0] MultLoop_acc_619_itm_1;
  wire [23:0] nl_MultLoop_acc_619_itm_1;
  reg [21:0] MultLoop_acc_618_itm_1;
  wire [23:0] nl_MultLoop_acc_618_itm_1;
  reg [21:0] MultLoop_acc_617_itm_1;
  wire [23:0] nl_MultLoop_acc_617_itm_1;
  reg [21:0] MultLoop_acc_616_itm_1;
  wire [23:0] nl_MultLoop_acc_616_itm_1;
  reg [21:0] MultLoop_acc_615_itm_1;
  wire [23:0] nl_MultLoop_acc_615_itm_1;
  reg [21:0] MultLoop_acc_757_itm_1;
  wire [22:0] nl_MultLoop_acc_757_itm_1;
  reg [21:0] MultLoop_acc_756_itm_1;
  wire [23:0] nl_MultLoop_acc_756_itm_1;
  reg [21:0] MultLoop_acc_755_itm_1;
  wire [23:0] nl_MultLoop_acc_755_itm_1;
  reg [21:0] MultLoop_acc_754_itm_1;
  wire [23:0] nl_MultLoop_acc_754_itm_1;
  reg [21:0] MultLoop_acc_753_itm_1;
  wire [23:0] nl_MultLoop_acc_753_itm_1;
  reg [21:0] MultLoop_acc_752_itm_1;
  wire [23:0] nl_MultLoop_acc_752_itm_1;
  reg [21:0] MultLoop_acc_751_itm_1;
  wire [23:0] nl_MultLoop_acc_751_itm_1;
  reg [21:0] MultLoop_acc_750_itm_1;
  wire [23:0] nl_MultLoop_acc_750_itm_1;
  reg [21:0] MultLoop_acc_749_itm_1;
  wire [23:0] nl_MultLoop_acc_749_itm_1;
  reg [21:0] MultLoop_acc_748_itm_1;
  wire [23:0] nl_MultLoop_acc_748_itm_1;
  reg [21:0] MultLoop_acc_747_itm_1;
  wire [23:0] nl_MultLoop_acc_747_itm_1;
  reg [21:0] MultLoop_acc_746_itm_1;
  wire [23:0] nl_MultLoop_acc_746_itm_1;
  reg [21:0] MultLoop_acc_745_itm_1;
  wire [23:0] nl_MultLoop_acc_745_itm_1;
  reg [21:0] MultLoop_acc_744_itm_1;
  wire [23:0] nl_MultLoop_acc_744_itm_1;
  reg [21:0] MultLoop_acc_743_itm_1;
  wire [23:0] nl_MultLoop_acc_743_itm_1;
  reg [21:0] MultLoop_acc_742_itm_1;
  wire [23:0] nl_MultLoop_acc_742_itm_1;
  reg [21:0] MultLoop_acc_884_itm_1;
  wire [22:0] nl_MultLoop_acc_884_itm_1;
  reg [21:0] MultLoop_acc_883_itm_1;
  wire [23:0] nl_MultLoop_acc_883_itm_1;
  reg [21:0] MultLoop_acc_882_itm_1;
  wire [23:0] nl_MultLoop_acc_882_itm_1;
  reg [21:0] MultLoop_acc_881_itm_1;
  wire [23:0] nl_MultLoop_acc_881_itm_1;
  reg [21:0] MultLoop_acc_880_itm_1;
  wire [23:0] nl_MultLoop_acc_880_itm_1;
  reg [21:0] MultLoop_acc_879_itm_1;
  wire [23:0] nl_MultLoop_acc_879_itm_1;
  reg [21:0] MultLoop_acc_878_itm_1;
  wire [23:0] nl_MultLoop_acc_878_itm_1;
  reg [21:0] MultLoop_acc_877_itm_1;
  wire [23:0] nl_MultLoop_acc_877_itm_1;
  reg [21:0] MultLoop_acc_876_itm_1;
  wire [23:0] nl_MultLoop_acc_876_itm_1;
  reg [21:0] MultLoop_acc_875_itm_1;
  wire [23:0] nl_MultLoop_acc_875_itm_1;
  reg [21:0] MultLoop_acc_874_itm_1;
  wire [23:0] nl_MultLoop_acc_874_itm_1;
  reg [21:0] MultLoop_acc_873_itm_1;
  wire [23:0] nl_MultLoop_acc_873_itm_1;
  reg [21:0] MultLoop_acc_872_itm_1;
  wire [23:0] nl_MultLoop_acc_872_itm_1;
  reg [21:0] MultLoop_acc_871_itm_1;
  wire [23:0] nl_MultLoop_acc_871_itm_1;
  reg [21:0] MultLoop_acc_870_itm_1;
  wire [23:0] nl_MultLoop_acc_870_itm_1;
  reg [21:0] MultLoop_acc_869_itm_1;
  wire [23:0] nl_MultLoop_acc_869_itm_1;
  reg [21:0] MultLoop_acc_1011_itm_1;
  wire [22:0] nl_MultLoop_acc_1011_itm_1;
  reg [21:0] MultLoop_acc_1010_itm_1;
  wire [23:0] nl_MultLoop_acc_1010_itm_1;
  reg [21:0] MultLoop_acc_1009_itm_1;
  wire [23:0] nl_MultLoop_acc_1009_itm_1;
  reg [21:0] MultLoop_acc_1008_itm_1;
  wire [23:0] nl_MultLoop_acc_1008_itm_1;
  reg [21:0] MultLoop_acc_1007_itm_1;
  wire [23:0] nl_MultLoop_acc_1007_itm_1;
  reg [21:0] MultLoop_acc_1006_itm_1;
  wire [23:0] nl_MultLoop_acc_1006_itm_1;
  reg [21:0] MultLoop_acc_1005_itm_1;
  wire [23:0] nl_MultLoop_acc_1005_itm_1;
  reg [21:0] MultLoop_acc_1004_itm_1;
  wire [23:0] nl_MultLoop_acc_1004_itm_1;
  reg [21:0] MultLoop_acc_1003_itm_1;
  wire [23:0] nl_MultLoop_acc_1003_itm_1;
  reg [21:0] MultLoop_acc_1002_itm_1;
  wire [23:0] nl_MultLoop_acc_1002_itm_1;
  reg [21:0] MultLoop_acc_1001_itm_1;
  wire [23:0] nl_MultLoop_acc_1001_itm_1;
  reg [21:0] MultLoop_acc_1000_itm_1;
  wire [23:0] nl_MultLoop_acc_1000_itm_1;
  reg [21:0] MultLoop_acc_999_itm_1;
  wire [23:0] nl_MultLoop_acc_999_itm_1;
  reg [21:0] MultLoop_acc_998_itm_1;
  wire [23:0] nl_MultLoop_acc_998_itm_1;
  reg [21:0] MultLoop_acc_997_itm_1;
  wire [23:0] nl_MultLoop_acc_997_itm_1;
  reg [21:0] MultLoop_acc_996_itm_1;
  wire [23:0] nl_MultLoop_acc_996_itm_1;
  reg [21:0] MultLoop_acc_1138_itm_1;
  wire [22:0] nl_MultLoop_acc_1138_itm_1;
  reg [21:0] MultLoop_acc_1137_itm_1;
  wire [23:0] nl_MultLoop_acc_1137_itm_1;
  reg [21:0] MultLoop_acc_1136_itm_1;
  wire [23:0] nl_MultLoop_acc_1136_itm_1;
  reg [21:0] MultLoop_acc_1135_itm_1;
  wire [23:0] nl_MultLoop_acc_1135_itm_1;
  reg [21:0] MultLoop_acc_1134_itm_1;
  wire [23:0] nl_MultLoop_acc_1134_itm_1;
  reg [21:0] MultLoop_acc_1133_itm_1;
  wire [23:0] nl_MultLoop_acc_1133_itm_1;
  reg [21:0] MultLoop_acc_1132_itm_1;
  wire [23:0] nl_MultLoop_acc_1132_itm_1;
  reg [21:0] MultLoop_acc_1131_itm_1;
  wire [23:0] nl_MultLoop_acc_1131_itm_1;
  reg [21:0] MultLoop_acc_1130_itm_1;
  wire [23:0] nl_MultLoop_acc_1130_itm_1;
  reg [21:0] MultLoop_acc_1129_itm_1;
  wire [23:0] nl_MultLoop_acc_1129_itm_1;
  reg [21:0] MultLoop_acc_1128_itm_1;
  wire [23:0] nl_MultLoop_acc_1128_itm_1;
  reg [21:0] MultLoop_acc_1127_itm_1;
  wire [23:0] nl_MultLoop_acc_1127_itm_1;
  reg [21:0] MultLoop_acc_1126_itm_1;
  wire [23:0] nl_MultLoop_acc_1126_itm_1;
  reg [21:0] MultLoop_acc_1125_itm_1;
  wire [23:0] nl_MultLoop_acc_1125_itm_1;
  reg [21:0] MultLoop_acc_1124_itm_1;
  wire [23:0] nl_MultLoop_acc_1124_itm_1;
  reg [21:0] MultLoop_acc_1123_itm_1;
  wire [23:0] nl_MultLoop_acc_1123_itm_1;
  reg [21:0] MultLoop_acc_1265_itm_1;
  wire [22:0] nl_MultLoop_acc_1265_itm_1;
  reg [21:0] MultLoop_acc_1264_itm_1;
  wire [23:0] nl_MultLoop_acc_1264_itm_1;
  reg [21:0] MultLoop_acc_1263_itm_1;
  wire [23:0] nl_MultLoop_acc_1263_itm_1;
  reg [21:0] MultLoop_acc_1262_itm_1;
  wire [23:0] nl_MultLoop_acc_1262_itm_1;
  reg [21:0] MultLoop_acc_1261_itm_1;
  wire [23:0] nl_MultLoop_acc_1261_itm_1;
  reg [21:0] MultLoop_acc_1260_itm_1;
  wire [23:0] nl_MultLoop_acc_1260_itm_1;
  reg [21:0] MultLoop_acc_1259_itm_1;
  wire [23:0] nl_MultLoop_acc_1259_itm_1;
  reg [21:0] MultLoop_acc_1258_itm_1;
  wire [23:0] nl_MultLoop_acc_1258_itm_1;
  reg [21:0] MultLoop_acc_1257_itm_1;
  wire [23:0] nl_MultLoop_acc_1257_itm_1;
  reg [21:0] MultLoop_acc_1256_itm_1;
  wire [23:0] nl_MultLoop_acc_1256_itm_1;
  reg [21:0] MultLoop_acc_1255_itm_1;
  wire [23:0] nl_MultLoop_acc_1255_itm_1;
  reg [21:0] MultLoop_acc_1254_itm_1;
  wire [23:0] nl_MultLoop_acc_1254_itm_1;
  reg [21:0] MultLoop_acc_1253_itm_1;
  wire [23:0] nl_MultLoop_acc_1253_itm_1;
  reg [21:0] MultLoop_acc_1252_itm_1;
  wire [23:0] nl_MultLoop_acc_1252_itm_1;
  reg [21:0] MultLoop_acc_1251_itm_1;
  wire [23:0] nl_MultLoop_acc_1251_itm_1;
  reg [21:0] MultLoop_acc_1250_itm_1;
  wire [23:0] nl_MultLoop_acc_1250_itm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289;
  wire [21:0] MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [21:0] MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;
  wire [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9;

  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[21:0] MultLoop_acc_1249_nl;
  wire[22:0] nl_MultLoop_acc_1249_nl;
  wire[21:0] MultLoop_acc_1217_nl;
  wire[22:0] nl_MultLoop_acc_1217_nl;
  wire[10:0] MultLoop_acc_1289_nl;
  wire[11:0] nl_MultLoop_acc_1289_nl;
  wire[28:0] MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1216_nl;
  wire[22:0] nl_MultLoop_acc_1216_nl;
  wire[28:0] MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1248_nl;
  wire[22:0] nl_MultLoop_acc_1248_nl;
  wire[21:0] MultLoop_acc_1215_nl;
  wire[22:0] nl_MultLoop_acc_1215_nl;
  wire[28:0] MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1214_nl;
  wire[22:0] nl_MultLoop_acc_1214_nl;
  wire[28:0] MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1213_nl;
  wire[22:0] nl_MultLoop_acc_1213_nl;
  wire[28:0] MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1212_nl;
  wire[22:0] nl_MultLoop_acc_1212_nl;
  wire[28:0] MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1211_nl;
  wire[22:0] nl_MultLoop_acc_1211_nl;
  wire[28:0] MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1210_nl;
  wire[22:0] nl_MultLoop_acc_1210_nl;
  wire[28:0] MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1209_nl;
  wire[22:0] nl_MultLoop_acc_1209_nl;
  wire[28:0] MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1208_nl;
  wire[22:0] nl_MultLoop_acc_1208_nl;
  wire[28:0] MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1207_nl;
  wire[22:0] nl_MultLoop_acc_1207_nl;
  wire[28:0] MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1206_nl;
  wire[22:0] nl_MultLoop_acc_1206_nl;
  wire[28:0] MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1205_nl;
  wire[22:0] nl_MultLoop_acc_1205_nl;
  wire[28:0] MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1204_nl;
  wire[22:0] nl_MultLoop_acc_1204_nl;
  wire[28:0] MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1203_nl;
  wire[22:0] nl_MultLoop_acc_1203_nl;
  wire[28:0] MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1202_nl;
  wire[22:0] nl_MultLoop_acc_1202_nl;
  wire[28:0] MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1201_nl;
  wire[22:0] nl_MultLoop_acc_1201_nl;
  wire[28:0] MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1200_nl;
  wire[22:0] nl_MultLoop_acc_1200_nl;
  wire[28:0] MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1199_nl;
  wire[22:0] nl_MultLoop_acc_1199_nl;
  wire[28:0] MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1198_nl;
  wire[22:0] nl_MultLoop_acc_1198_nl;
  wire[28:0] MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1197_nl;
  wire[22:0] nl_MultLoop_acc_1197_nl;
  wire[28:0] MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1196_nl;
  wire[22:0] nl_MultLoop_acc_1196_nl;
  wire[28:0] MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1195_nl;
  wire[22:0] nl_MultLoop_acc_1195_nl;
  wire[28:0] MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1194_nl;
  wire[22:0] nl_MultLoop_acc_1194_nl;
  wire[28:0] MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1193_nl;
  wire[22:0] nl_MultLoop_acc_1193_nl;
  wire[28:0] MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1192_nl;
  wire[22:0] nl_MultLoop_acc_1192_nl;
  wire[28:0] MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1191_nl;
  wire[22:0] nl_MultLoop_acc_1191_nl;
  wire[28:0] MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1190_nl;
  wire[22:0] nl_MultLoop_acc_1190_nl;
  wire[28:0] MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1189_nl;
  wire[22:0] nl_MultLoop_acc_1189_nl;
  wire[28:0] MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1188_nl;
  wire[22:0] nl_MultLoop_acc_1188_nl;
  wire[28:0] MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1187_nl;
  wire[22:0] nl_MultLoop_acc_1187_nl;
  wire[28:0] MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1186_nl;
  wire[22:0] nl_MultLoop_acc_1186_nl;
  wire[28:0] MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1185_nl;
  wire[22:0] nl_MultLoop_acc_1185_nl;
  wire[28:0] MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1184_nl;
  wire[22:0] nl_MultLoop_acc_1184_nl;
  wire[28:0] MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1183_nl;
  wire[22:0] nl_MultLoop_acc_1183_nl;
  wire[28:0] MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1182_nl;
  wire[22:0] nl_MultLoop_acc_1182_nl;
  wire[28:0] MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1181_nl;
  wire[22:0] nl_MultLoop_acc_1181_nl;
  wire[28:0] MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1180_nl;
  wire[22:0] nl_MultLoop_acc_1180_nl;
  wire[28:0] MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1179_nl;
  wire[22:0] nl_MultLoop_acc_1179_nl;
  wire[28:0] MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1178_nl;
  wire[22:0] nl_MultLoop_acc_1178_nl;
  wire[28:0] MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1177_nl;
  wire[22:0] nl_MultLoop_acc_1177_nl;
  wire[28:0] MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1176_nl;
  wire[22:0] nl_MultLoop_acc_1176_nl;
  wire[28:0] MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1175_nl;
  wire[22:0] nl_MultLoop_acc_1175_nl;
  wire[28:0] MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1174_nl;
  wire[22:0] nl_MultLoop_acc_1174_nl;
  wire[28:0] MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1173_nl;
  wire[22:0] nl_MultLoop_acc_1173_nl;
  wire[28:0] MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1172_nl;
  wire[22:0] nl_MultLoop_acc_1172_nl;
  wire[28:0] MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1171_nl;
  wire[22:0] nl_MultLoop_acc_1171_nl;
  wire[28:0] MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1170_nl;
  wire[22:0] nl_MultLoop_acc_1170_nl;
  wire[28:0] MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1169_nl;
  wire[22:0] nl_MultLoop_acc_1169_nl;
  wire[28:0] MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1168_nl;
  wire[22:0] nl_MultLoop_acc_1168_nl;
  wire[28:0] MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1167_nl;
  wire[22:0] nl_MultLoop_acc_1167_nl;
  wire[28:0] MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1166_nl;
  wire[22:0] nl_MultLoop_acc_1166_nl;
  wire[28:0] MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1165_nl;
  wire[22:0] nl_MultLoop_acc_1165_nl;
  wire[28:0] MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1164_nl;
  wire[22:0] nl_MultLoop_acc_1164_nl;
  wire[28:0] MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1163_nl;
  wire[22:0] nl_MultLoop_acc_1163_nl;
  wire[28:0] MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1162_nl;
  wire[22:0] nl_MultLoop_acc_1162_nl;
  wire[28:0] MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1161_nl;
  wire[22:0] nl_MultLoop_acc_1161_nl;
  wire[28:0] MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1160_nl;
  wire[22:0] nl_MultLoop_acc_1160_nl;
  wire[28:0] MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1159_nl;
  wire[22:0] nl_MultLoop_acc_1159_nl;
  wire[28:0] MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1158_nl;
  wire[22:0] nl_MultLoop_acc_1158_nl;
  wire[28:0] MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1157_nl;
  wire[22:0] nl_MultLoop_acc_1157_nl;
  wire[28:0] MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1156_nl;
  wire[22:0] nl_MultLoop_acc_1156_nl;
  wire[28:0] MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1155_nl;
  wire[22:0] nl_MultLoop_acc_1155_nl;
  wire[28:0] MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1154_nl;
  wire[22:0] nl_MultLoop_acc_1154_nl;
  wire[28:0] MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1122_nl;
  wire[22:0] nl_MultLoop_acc_1122_nl;
  wire[21:0] MultLoop_acc_1090_nl;
  wire[22:0] nl_MultLoop_acc_1090_nl;
  wire[10:0] MultLoop_acc_1288_nl;
  wire[11:0] nl_MultLoop_acc_1288_nl;
  wire[28:0] MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1089_nl;
  wire[22:0] nl_MultLoop_acc_1089_nl;
  wire[28:0] MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1121_nl;
  wire[22:0] nl_MultLoop_acc_1121_nl;
  wire[21:0] MultLoop_acc_1088_nl;
  wire[22:0] nl_MultLoop_acc_1088_nl;
  wire[28:0] MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1087_nl;
  wire[22:0] nl_MultLoop_acc_1087_nl;
  wire[28:0] MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1086_nl;
  wire[22:0] nl_MultLoop_acc_1086_nl;
  wire[28:0] MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1085_nl;
  wire[22:0] nl_MultLoop_acc_1085_nl;
  wire[28:0] MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1084_nl;
  wire[22:0] nl_MultLoop_acc_1084_nl;
  wire[28:0] MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1083_nl;
  wire[22:0] nl_MultLoop_acc_1083_nl;
  wire[28:0] MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1082_nl;
  wire[22:0] nl_MultLoop_acc_1082_nl;
  wire[28:0] MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1081_nl;
  wire[22:0] nl_MultLoop_acc_1081_nl;
  wire[28:0] MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1080_nl;
  wire[22:0] nl_MultLoop_acc_1080_nl;
  wire[28:0] MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1079_nl;
  wire[22:0] nl_MultLoop_acc_1079_nl;
  wire[28:0] MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1078_nl;
  wire[22:0] nl_MultLoop_acc_1078_nl;
  wire[28:0] MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1077_nl;
  wire[22:0] nl_MultLoop_acc_1077_nl;
  wire[28:0] MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1076_nl;
  wire[22:0] nl_MultLoop_acc_1076_nl;
  wire[28:0] MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1075_nl;
  wire[22:0] nl_MultLoop_acc_1075_nl;
  wire[28:0] MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1074_nl;
  wire[22:0] nl_MultLoop_acc_1074_nl;
  wire[28:0] MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1073_nl;
  wire[22:0] nl_MultLoop_acc_1073_nl;
  wire[28:0] MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1072_nl;
  wire[22:0] nl_MultLoop_acc_1072_nl;
  wire[28:0] MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1071_nl;
  wire[22:0] nl_MultLoop_acc_1071_nl;
  wire[28:0] MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1070_nl;
  wire[22:0] nl_MultLoop_acc_1070_nl;
  wire[28:0] MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1069_nl;
  wire[22:0] nl_MultLoop_acc_1069_nl;
  wire[28:0] MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1068_nl;
  wire[22:0] nl_MultLoop_acc_1068_nl;
  wire[28:0] MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1067_nl;
  wire[22:0] nl_MultLoop_acc_1067_nl;
  wire[28:0] MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1066_nl;
  wire[22:0] nl_MultLoop_acc_1066_nl;
  wire[28:0] MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1065_nl;
  wire[22:0] nl_MultLoop_acc_1065_nl;
  wire[28:0] MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1064_nl;
  wire[22:0] nl_MultLoop_acc_1064_nl;
  wire[28:0] MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1063_nl;
  wire[22:0] nl_MultLoop_acc_1063_nl;
  wire[28:0] MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1062_nl;
  wire[22:0] nl_MultLoop_acc_1062_nl;
  wire[28:0] MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1061_nl;
  wire[22:0] nl_MultLoop_acc_1061_nl;
  wire[28:0] MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1060_nl;
  wire[22:0] nl_MultLoop_acc_1060_nl;
  wire[28:0] MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1059_nl;
  wire[22:0] nl_MultLoop_acc_1059_nl;
  wire[28:0] MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1058_nl;
  wire[22:0] nl_MultLoop_acc_1058_nl;
  wire[28:0] MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1057_nl;
  wire[22:0] nl_MultLoop_acc_1057_nl;
  wire[28:0] MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1056_nl;
  wire[22:0] nl_MultLoop_acc_1056_nl;
  wire[28:0] MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1055_nl;
  wire[22:0] nl_MultLoop_acc_1055_nl;
  wire[28:0] MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1054_nl;
  wire[22:0] nl_MultLoop_acc_1054_nl;
  wire[28:0] MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1053_nl;
  wire[22:0] nl_MultLoop_acc_1053_nl;
  wire[28:0] MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1052_nl;
  wire[22:0] nl_MultLoop_acc_1052_nl;
  wire[28:0] MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1051_nl;
  wire[22:0] nl_MultLoop_acc_1051_nl;
  wire[28:0] MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1050_nl;
  wire[22:0] nl_MultLoop_acc_1050_nl;
  wire[28:0] MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1049_nl;
  wire[22:0] nl_MultLoop_acc_1049_nl;
  wire[28:0] MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1048_nl;
  wire[22:0] nl_MultLoop_acc_1048_nl;
  wire[28:0] MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1047_nl;
  wire[22:0] nl_MultLoop_acc_1047_nl;
  wire[28:0] MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1046_nl;
  wire[22:0] nl_MultLoop_acc_1046_nl;
  wire[28:0] MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1045_nl;
  wire[22:0] nl_MultLoop_acc_1045_nl;
  wire[28:0] MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1044_nl;
  wire[22:0] nl_MultLoop_acc_1044_nl;
  wire[28:0] MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1043_nl;
  wire[22:0] nl_MultLoop_acc_1043_nl;
  wire[28:0] MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1042_nl;
  wire[22:0] nl_MultLoop_acc_1042_nl;
  wire[28:0] MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1041_nl;
  wire[22:0] nl_MultLoop_acc_1041_nl;
  wire[28:0] MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1040_nl;
  wire[22:0] nl_MultLoop_acc_1040_nl;
  wire[28:0] MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1039_nl;
  wire[22:0] nl_MultLoop_acc_1039_nl;
  wire[28:0] MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1038_nl;
  wire[22:0] nl_MultLoop_acc_1038_nl;
  wire[28:0] MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1037_nl;
  wire[22:0] nl_MultLoop_acc_1037_nl;
  wire[28:0] MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1036_nl;
  wire[22:0] nl_MultLoop_acc_1036_nl;
  wire[28:0] MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1035_nl;
  wire[22:0] nl_MultLoop_acc_1035_nl;
  wire[28:0] MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1034_nl;
  wire[22:0] nl_MultLoop_acc_1034_nl;
  wire[28:0] MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1033_nl;
  wire[22:0] nl_MultLoop_acc_1033_nl;
  wire[28:0] MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1032_nl;
  wire[22:0] nl_MultLoop_acc_1032_nl;
  wire[28:0] MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1031_nl;
  wire[22:0] nl_MultLoop_acc_1031_nl;
  wire[28:0] MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1030_nl;
  wire[22:0] nl_MultLoop_acc_1030_nl;
  wire[28:0] MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1029_nl;
  wire[22:0] nl_MultLoop_acc_1029_nl;
  wire[28:0] MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1028_nl;
  wire[22:0] nl_MultLoop_acc_1028_nl;
  wire[28:0] MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1027_nl;
  wire[22:0] nl_MultLoop_acc_1027_nl;
  wire[28:0] MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_995_nl;
  wire[22:0] nl_MultLoop_acc_995_nl;
  wire[21:0] MultLoop_acc_963_nl;
  wire[22:0] nl_MultLoop_acc_963_nl;
  wire[10:0] MultLoop_acc_1287_nl;
  wire[11:0] nl_MultLoop_acc_1287_nl;
  wire[28:0] MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_962_nl;
  wire[22:0] nl_MultLoop_acc_962_nl;
  wire[28:0] MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_994_nl;
  wire[22:0] nl_MultLoop_acc_994_nl;
  wire[21:0] MultLoop_acc_961_nl;
  wire[22:0] nl_MultLoop_acc_961_nl;
  wire[28:0] MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_960_nl;
  wire[22:0] nl_MultLoop_acc_960_nl;
  wire[28:0] MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_959_nl;
  wire[22:0] nl_MultLoop_acc_959_nl;
  wire[28:0] MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_958_nl;
  wire[22:0] nl_MultLoop_acc_958_nl;
  wire[28:0] MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_957_nl;
  wire[22:0] nl_MultLoop_acc_957_nl;
  wire[28:0] MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_956_nl;
  wire[22:0] nl_MultLoop_acc_956_nl;
  wire[28:0] MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_955_nl;
  wire[22:0] nl_MultLoop_acc_955_nl;
  wire[28:0] MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_954_nl;
  wire[22:0] nl_MultLoop_acc_954_nl;
  wire[28:0] MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_953_nl;
  wire[22:0] nl_MultLoop_acc_953_nl;
  wire[28:0] MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_952_nl;
  wire[22:0] nl_MultLoop_acc_952_nl;
  wire[28:0] MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_951_nl;
  wire[22:0] nl_MultLoop_acc_951_nl;
  wire[28:0] MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_950_nl;
  wire[22:0] nl_MultLoop_acc_950_nl;
  wire[28:0] MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_949_nl;
  wire[22:0] nl_MultLoop_acc_949_nl;
  wire[28:0] MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_948_nl;
  wire[22:0] nl_MultLoop_acc_948_nl;
  wire[28:0] MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_947_nl;
  wire[22:0] nl_MultLoop_acc_947_nl;
  wire[28:0] MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_946_nl;
  wire[22:0] nl_MultLoop_acc_946_nl;
  wire[28:0] MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_945_nl;
  wire[22:0] nl_MultLoop_acc_945_nl;
  wire[28:0] MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_944_nl;
  wire[22:0] nl_MultLoop_acc_944_nl;
  wire[28:0] MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_943_nl;
  wire[22:0] nl_MultLoop_acc_943_nl;
  wire[28:0] MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_942_nl;
  wire[22:0] nl_MultLoop_acc_942_nl;
  wire[28:0] MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_941_nl;
  wire[22:0] nl_MultLoop_acc_941_nl;
  wire[28:0] MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_940_nl;
  wire[22:0] nl_MultLoop_acc_940_nl;
  wire[28:0] MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_939_nl;
  wire[22:0] nl_MultLoop_acc_939_nl;
  wire[28:0] MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_938_nl;
  wire[22:0] nl_MultLoop_acc_938_nl;
  wire[28:0] MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_937_nl;
  wire[22:0] nl_MultLoop_acc_937_nl;
  wire[28:0] MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_936_nl;
  wire[22:0] nl_MultLoop_acc_936_nl;
  wire[28:0] MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_935_nl;
  wire[22:0] nl_MultLoop_acc_935_nl;
  wire[28:0] MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_934_nl;
  wire[22:0] nl_MultLoop_acc_934_nl;
  wire[28:0] MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_933_nl;
  wire[22:0] nl_MultLoop_acc_933_nl;
  wire[28:0] MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_932_nl;
  wire[22:0] nl_MultLoop_acc_932_nl;
  wire[28:0] MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_931_nl;
  wire[22:0] nl_MultLoop_acc_931_nl;
  wire[28:0] MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_930_nl;
  wire[22:0] nl_MultLoop_acc_930_nl;
  wire[28:0] MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_929_nl;
  wire[22:0] nl_MultLoop_acc_929_nl;
  wire[28:0] MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_928_nl;
  wire[22:0] nl_MultLoop_acc_928_nl;
  wire[28:0] MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_927_nl;
  wire[22:0] nl_MultLoop_acc_927_nl;
  wire[28:0] MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_926_nl;
  wire[22:0] nl_MultLoop_acc_926_nl;
  wire[28:0] MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_925_nl;
  wire[22:0] nl_MultLoop_acc_925_nl;
  wire[28:0] MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_924_nl;
  wire[22:0] nl_MultLoop_acc_924_nl;
  wire[28:0] MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_923_nl;
  wire[22:0] nl_MultLoop_acc_923_nl;
  wire[28:0] MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_922_nl;
  wire[22:0] nl_MultLoop_acc_922_nl;
  wire[28:0] MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_921_nl;
  wire[22:0] nl_MultLoop_acc_921_nl;
  wire[28:0] MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_920_nl;
  wire[22:0] nl_MultLoop_acc_920_nl;
  wire[28:0] MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_919_nl;
  wire[22:0] nl_MultLoop_acc_919_nl;
  wire[28:0] MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_918_nl;
  wire[22:0] nl_MultLoop_acc_918_nl;
  wire[28:0] MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_917_nl;
  wire[22:0] nl_MultLoop_acc_917_nl;
  wire[28:0] MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_916_nl;
  wire[22:0] nl_MultLoop_acc_916_nl;
  wire[28:0] MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_915_nl;
  wire[22:0] nl_MultLoop_acc_915_nl;
  wire[28:0] MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_914_nl;
  wire[22:0] nl_MultLoop_acc_914_nl;
  wire[28:0] MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_913_nl;
  wire[22:0] nl_MultLoop_acc_913_nl;
  wire[28:0] MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_912_nl;
  wire[22:0] nl_MultLoop_acc_912_nl;
  wire[28:0] MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_911_nl;
  wire[22:0] nl_MultLoop_acc_911_nl;
  wire[28:0] MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_910_nl;
  wire[22:0] nl_MultLoop_acc_910_nl;
  wire[28:0] MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_909_nl;
  wire[22:0] nl_MultLoop_acc_909_nl;
  wire[28:0] MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_908_nl;
  wire[22:0] nl_MultLoop_acc_908_nl;
  wire[28:0] MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_907_nl;
  wire[22:0] nl_MultLoop_acc_907_nl;
  wire[28:0] MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_906_nl;
  wire[22:0] nl_MultLoop_acc_906_nl;
  wire[28:0] MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_905_nl;
  wire[22:0] nl_MultLoop_acc_905_nl;
  wire[28:0] MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_904_nl;
  wire[22:0] nl_MultLoop_acc_904_nl;
  wire[28:0] MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_903_nl;
  wire[22:0] nl_MultLoop_acc_903_nl;
  wire[28:0] MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_902_nl;
  wire[22:0] nl_MultLoop_acc_902_nl;
  wire[28:0] MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_901_nl;
  wire[22:0] nl_MultLoop_acc_901_nl;
  wire[28:0] MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_900_nl;
  wire[22:0] nl_MultLoop_acc_900_nl;
  wire[28:0] MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_868_nl;
  wire[22:0] nl_MultLoop_acc_868_nl;
  wire[21:0] MultLoop_acc_836_nl;
  wire[22:0] nl_MultLoop_acc_836_nl;
  wire[10:0] MultLoop_acc_1286_nl;
  wire[11:0] nl_MultLoop_acc_1286_nl;
  wire[28:0] MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_835_nl;
  wire[22:0] nl_MultLoop_acc_835_nl;
  wire[28:0] MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_867_nl;
  wire[22:0] nl_MultLoop_acc_867_nl;
  wire[21:0] MultLoop_acc_834_nl;
  wire[22:0] nl_MultLoop_acc_834_nl;
  wire[28:0] MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_833_nl;
  wire[22:0] nl_MultLoop_acc_833_nl;
  wire[28:0] MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_832_nl;
  wire[22:0] nl_MultLoop_acc_832_nl;
  wire[28:0] MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_831_nl;
  wire[22:0] nl_MultLoop_acc_831_nl;
  wire[28:0] MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_830_nl;
  wire[22:0] nl_MultLoop_acc_830_nl;
  wire[28:0] MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_829_nl;
  wire[22:0] nl_MultLoop_acc_829_nl;
  wire[28:0] MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_828_nl;
  wire[22:0] nl_MultLoop_acc_828_nl;
  wire[28:0] MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_827_nl;
  wire[22:0] nl_MultLoop_acc_827_nl;
  wire[28:0] MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_826_nl;
  wire[22:0] nl_MultLoop_acc_826_nl;
  wire[28:0] MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_825_nl;
  wire[22:0] nl_MultLoop_acc_825_nl;
  wire[28:0] MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_824_nl;
  wire[22:0] nl_MultLoop_acc_824_nl;
  wire[28:0] MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_823_nl;
  wire[22:0] nl_MultLoop_acc_823_nl;
  wire[28:0] MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_822_nl;
  wire[22:0] nl_MultLoop_acc_822_nl;
  wire[28:0] MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_821_nl;
  wire[22:0] nl_MultLoop_acc_821_nl;
  wire[28:0] MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_820_nl;
  wire[22:0] nl_MultLoop_acc_820_nl;
  wire[28:0] MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_819_nl;
  wire[22:0] nl_MultLoop_acc_819_nl;
  wire[28:0] MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_818_nl;
  wire[22:0] nl_MultLoop_acc_818_nl;
  wire[28:0] MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_817_nl;
  wire[22:0] nl_MultLoop_acc_817_nl;
  wire[28:0] MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_816_nl;
  wire[22:0] nl_MultLoop_acc_816_nl;
  wire[28:0] MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_815_nl;
  wire[22:0] nl_MultLoop_acc_815_nl;
  wire[28:0] MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_814_nl;
  wire[22:0] nl_MultLoop_acc_814_nl;
  wire[28:0] MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_813_nl;
  wire[22:0] nl_MultLoop_acc_813_nl;
  wire[28:0] MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_812_nl;
  wire[22:0] nl_MultLoop_acc_812_nl;
  wire[28:0] MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_811_nl;
  wire[22:0] nl_MultLoop_acc_811_nl;
  wire[28:0] MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_810_nl;
  wire[22:0] nl_MultLoop_acc_810_nl;
  wire[28:0] MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_809_nl;
  wire[22:0] nl_MultLoop_acc_809_nl;
  wire[28:0] MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_808_nl;
  wire[22:0] nl_MultLoop_acc_808_nl;
  wire[28:0] MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_807_nl;
  wire[22:0] nl_MultLoop_acc_807_nl;
  wire[28:0] MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_806_nl;
  wire[22:0] nl_MultLoop_acc_806_nl;
  wire[28:0] MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_805_nl;
  wire[22:0] nl_MultLoop_acc_805_nl;
  wire[28:0] MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_804_nl;
  wire[22:0] nl_MultLoop_acc_804_nl;
  wire[28:0] MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_803_nl;
  wire[22:0] nl_MultLoop_acc_803_nl;
  wire[28:0] MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_802_nl;
  wire[22:0] nl_MultLoop_acc_802_nl;
  wire[28:0] MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_801_nl;
  wire[22:0] nl_MultLoop_acc_801_nl;
  wire[28:0] MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_800_nl;
  wire[22:0] nl_MultLoop_acc_800_nl;
  wire[28:0] MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_799_nl;
  wire[22:0] nl_MultLoop_acc_799_nl;
  wire[28:0] MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_798_nl;
  wire[22:0] nl_MultLoop_acc_798_nl;
  wire[28:0] MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_797_nl;
  wire[22:0] nl_MultLoop_acc_797_nl;
  wire[28:0] MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_796_nl;
  wire[22:0] nl_MultLoop_acc_796_nl;
  wire[28:0] MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_795_nl;
  wire[22:0] nl_MultLoop_acc_795_nl;
  wire[28:0] MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_794_nl;
  wire[22:0] nl_MultLoop_acc_794_nl;
  wire[28:0] MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_793_nl;
  wire[22:0] nl_MultLoop_acc_793_nl;
  wire[28:0] MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_792_nl;
  wire[22:0] nl_MultLoop_acc_792_nl;
  wire[28:0] MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_791_nl;
  wire[22:0] nl_MultLoop_acc_791_nl;
  wire[28:0] MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_790_nl;
  wire[22:0] nl_MultLoop_acc_790_nl;
  wire[28:0] MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_789_nl;
  wire[22:0] nl_MultLoop_acc_789_nl;
  wire[28:0] MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_788_nl;
  wire[22:0] nl_MultLoop_acc_788_nl;
  wire[28:0] MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_787_nl;
  wire[22:0] nl_MultLoop_acc_787_nl;
  wire[28:0] MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_786_nl;
  wire[22:0] nl_MultLoop_acc_786_nl;
  wire[28:0] MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_785_nl;
  wire[22:0] nl_MultLoop_acc_785_nl;
  wire[28:0] MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_784_nl;
  wire[22:0] nl_MultLoop_acc_784_nl;
  wire[28:0] MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_783_nl;
  wire[22:0] nl_MultLoop_acc_783_nl;
  wire[28:0] MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_782_nl;
  wire[22:0] nl_MultLoop_acc_782_nl;
  wire[28:0] MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_781_nl;
  wire[22:0] nl_MultLoop_acc_781_nl;
  wire[28:0] MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_780_nl;
  wire[22:0] nl_MultLoop_acc_780_nl;
  wire[28:0] MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_779_nl;
  wire[22:0] nl_MultLoop_acc_779_nl;
  wire[28:0] MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_778_nl;
  wire[22:0] nl_MultLoop_acc_778_nl;
  wire[28:0] MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_777_nl;
  wire[22:0] nl_MultLoop_acc_777_nl;
  wire[28:0] MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_776_nl;
  wire[22:0] nl_MultLoop_acc_776_nl;
  wire[28:0] MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_775_nl;
  wire[22:0] nl_MultLoop_acc_775_nl;
  wire[28:0] MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_774_nl;
  wire[22:0] nl_MultLoop_acc_774_nl;
  wire[28:0] MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_773_nl;
  wire[22:0] nl_MultLoop_acc_773_nl;
  wire[28:0] MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_741_nl;
  wire[22:0] nl_MultLoop_acc_741_nl;
  wire[21:0] MultLoop_acc_709_nl;
  wire[22:0] nl_MultLoop_acc_709_nl;
  wire[10:0] MultLoop_acc_1285_nl;
  wire[11:0] nl_MultLoop_acc_1285_nl;
  wire[28:0] MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_708_nl;
  wire[22:0] nl_MultLoop_acc_708_nl;
  wire[28:0] MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_740_nl;
  wire[22:0] nl_MultLoop_acc_740_nl;
  wire[21:0] MultLoop_acc_707_nl;
  wire[22:0] nl_MultLoop_acc_707_nl;
  wire[28:0] MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_706_nl;
  wire[22:0] nl_MultLoop_acc_706_nl;
  wire[28:0] MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_705_nl;
  wire[22:0] nl_MultLoop_acc_705_nl;
  wire[28:0] MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_704_nl;
  wire[22:0] nl_MultLoop_acc_704_nl;
  wire[28:0] MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_703_nl;
  wire[22:0] nl_MultLoop_acc_703_nl;
  wire[28:0] MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_702_nl;
  wire[22:0] nl_MultLoop_acc_702_nl;
  wire[28:0] MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_701_nl;
  wire[22:0] nl_MultLoop_acc_701_nl;
  wire[28:0] MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_700_nl;
  wire[22:0] nl_MultLoop_acc_700_nl;
  wire[28:0] MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_699_nl;
  wire[22:0] nl_MultLoop_acc_699_nl;
  wire[28:0] MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_698_nl;
  wire[22:0] nl_MultLoop_acc_698_nl;
  wire[28:0] MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_697_nl;
  wire[22:0] nl_MultLoop_acc_697_nl;
  wire[28:0] MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_696_nl;
  wire[22:0] nl_MultLoop_acc_696_nl;
  wire[28:0] MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_695_nl;
  wire[22:0] nl_MultLoop_acc_695_nl;
  wire[28:0] MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_694_nl;
  wire[22:0] nl_MultLoop_acc_694_nl;
  wire[28:0] MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_693_nl;
  wire[22:0] nl_MultLoop_acc_693_nl;
  wire[28:0] MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_692_nl;
  wire[22:0] nl_MultLoop_acc_692_nl;
  wire[28:0] MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_691_nl;
  wire[22:0] nl_MultLoop_acc_691_nl;
  wire[28:0] MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_690_nl;
  wire[22:0] nl_MultLoop_acc_690_nl;
  wire[28:0] MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_689_nl;
  wire[22:0] nl_MultLoop_acc_689_nl;
  wire[28:0] MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_688_nl;
  wire[22:0] nl_MultLoop_acc_688_nl;
  wire[28:0] MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_687_nl;
  wire[22:0] nl_MultLoop_acc_687_nl;
  wire[28:0] MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_686_nl;
  wire[22:0] nl_MultLoop_acc_686_nl;
  wire[28:0] MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_685_nl;
  wire[22:0] nl_MultLoop_acc_685_nl;
  wire[28:0] MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_684_nl;
  wire[22:0] nl_MultLoop_acc_684_nl;
  wire[28:0] MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_683_nl;
  wire[22:0] nl_MultLoop_acc_683_nl;
  wire[28:0] MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_682_nl;
  wire[22:0] nl_MultLoop_acc_682_nl;
  wire[28:0] MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_681_nl;
  wire[22:0] nl_MultLoop_acc_681_nl;
  wire[28:0] MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_680_nl;
  wire[22:0] nl_MultLoop_acc_680_nl;
  wire[28:0] MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_679_nl;
  wire[22:0] nl_MultLoop_acc_679_nl;
  wire[28:0] MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_678_nl;
  wire[22:0] nl_MultLoop_acc_678_nl;
  wire[28:0] MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_677_nl;
  wire[22:0] nl_MultLoop_acc_677_nl;
  wire[28:0] MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_676_nl;
  wire[22:0] nl_MultLoop_acc_676_nl;
  wire[28:0] MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_675_nl;
  wire[22:0] nl_MultLoop_acc_675_nl;
  wire[28:0] MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_674_nl;
  wire[22:0] nl_MultLoop_acc_674_nl;
  wire[28:0] MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_673_nl;
  wire[22:0] nl_MultLoop_acc_673_nl;
  wire[28:0] MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_672_nl;
  wire[22:0] nl_MultLoop_acc_672_nl;
  wire[28:0] MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_671_nl;
  wire[22:0] nl_MultLoop_acc_671_nl;
  wire[28:0] MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_670_nl;
  wire[22:0] nl_MultLoop_acc_670_nl;
  wire[28:0] MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_669_nl;
  wire[22:0] nl_MultLoop_acc_669_nl;
  wire[28:0] MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_668_nl;
  wire[22:0] nl_MultLoop_acc_668_nl;
  wire[28:0] MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_667_nl;
  wire[22:0] nl_MultLoop_acc_667_nl;
  wire[28:0] MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_666_nl;
  wire[22:0] nl_MultLoop_acc_666_nl;
  wire[28:0] MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_665_nl;
  wire[22:0] nl_MultLoop_acc_665_nl;
  wire[28:0] MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_664_nl;
  wire[22:0] nl_MultLoop_acc_664_nl;
  wire[28:0] MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_663_nl;
  wire[22:0] nl_MultLoop_acc_663_nl;
  wire[28:0] MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_662_nl;
  wire[22:0] nl_MultLoop_acc_662_nl;
  wire[28:0] MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_661_nl;
  wire[22:0] nl_MultLoop_acc_661_nl;
  wire[28:0] MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_660_nl;
  wire[22:0] nl_MultLoop_acc_660_nl;
  wire[28:0] MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_659_nl;
  wire[22:0] nl_MultLoop_acc_659_nl;
  wire[28:0] MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_658_nl;
  wire[22:0] nl_MultLoop_acc_658_nl;
  wire[28:0] MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_657_nl;
  wire[22:0] nl_MultLoop_acc_657_nl;
  wire[28:0] MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_656_nl;
  wire[22:0] nl_MultLoop_acc_656_nl;
  wire[28:0] MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_655_nl;
  wire[22:0] nl_MultLoop_acc_655_nl;
  wire[28:0] MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_654_nl;
  wire[22:0] nl_MultLoop_acc_654_nl;
  wire[28:0] MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_653_nl;
  wire[22:0] nl_MultLoop_acc_653_nl;
  wire[28:0] MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_652_nl;
  wire[22:0] nl_MultLoop_acc_652_nl;
  wire[28:0] MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_651_nl;
  wire[22:0] nl_MultLoop_acc_651_nl;
  wire[28:0] MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_650_nl;
  wire[22:0] nl_MultLoop_acc_650_nl;
  wire[28:0] MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_649_nl;
  wire[22:0] nl_MultLoop_acc_649_nl;
  wire[28:0] MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_648_nl;
  wire[22:0] nl_MultLoop_acc_648_nl;
  wire[28:0] MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_647_nl;
  wire[22:0] nl_MultLoop_acc_647_nl;
  wire[28:0] MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_646_nl;
  wire[22:0] nl_MultLoop_acc_646_nl;
  wire[28:0] MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_614_nl;
  wire[22:0] nl_MultLoop_acc_614_nl;
  wire[21:0] MultLoop_acc_582_nl;
  wire[22:0] nl_MultLoop_acc_582_nl;
  wire[10:0] MultLoop_acc_1284_nl;
  wire[11:0] nl_MultLoop_acc_1284_nl;
  wire[28:0] MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_581_nl;
  wire[22:0] nl_MultLoop_acc_581_nl;
  wire[28:0] MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_613_nl;
  wire[22:0] nl_MultLoop_acc_613_nl;
  wire[21:0] MultLoop_acc_580_nl;
  wire[22:0] nl_MultLoop_acc_580_nl;
  wire[28:0] MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_579_nl;
  wire[22:0] nl_MultLoop_acc_579_nl;
  wire[28:0] MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_578_nl;
  wire[22:0] nl_MultLoop_acc_578_nl;
  wire[28:0] MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_577_nl;
  wire[22:0] nl_MultLoop_acc_577_nl;
  wire[28:0] MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_576_nl;
  wire[22:0] nl_MultLoop_acc_576_nl;
  wire[28:0] MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_575_nl;
  wire[22:0] nl_MultLoop_acc_575_nl;
  wire[28:0] MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_574_nl;
  wire[22:0] nl_MultLoop_acc_574_nl;
  wire[28:0] MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_573_nl;
  wire[22:0] nl_MultLoop_acc_573_nl;
  wire[28:0] MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_572_nl;
  wire[22:0] nl_MultLoop_acc_572_nl;
  wire[28:0] MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_571_nl;
  wire[22:0] nl_MultLoop_acc_571_nl;
  wire[28:0] MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_570_nl;
  wire[22:0] nl_MultLoop_acc_570_nl;
  wire[28:0] MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_569_nl;
  wire[22:0] nl_MultLoop_acc_569_nl;
  wire[28:0] MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_568_nl;
  wire[22:0] nl_MultLoop_acc_568_nl;
  wire[28:0] MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_567_nl;
  wire[22:0] nl_MultLoop_acc_567_nl;
  wire[28:0] MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_566_nl;
  wire[22:0] nl_MultLoop_acc_566_nl;
  wire[28:0] MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_565_nl;
  wire[22:0] nl_MultLoop_acc_565_nl;
  wire[28:0] MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_564_nl;
  wire[22:0] nl_MultLoop_acc_564_nl;
  wire[28:0] MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_563_nl;
  wire[22:0] nl_MultLoop_acc_563_nl;
  wire[28:0] MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_562_nl;
  wire[22:0] nl_MultLoop_acc_562_nl;
  wire[28:0] MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_561_nl;
  wire[22:0] nl_MultLoop_acc_561_nl;
  wire[28:0] MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_560_nl;
  wire[22:0] nl_MultLoop_acc_560_nl;
  wire[28:0] MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_559_nl;
  wire[22:0] nl_MultLoop_acc_559_nl;
  wire[28:0] MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_558_nl;
  wire[22:0] nl_MultLoop_acc_558_nl;
  wire[28:0] MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_557_nl;
  wire[22:0] nl_MultLoop_acc_557_nl;
  wire[28:0] MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_556_nl;
  wire[22:0] nl_MultLoop_acc_556_nl;
  wire[28:0] MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_555_nl;
  wire[22:0] nl_MultLoop_acc_555_nl;
  wire[28:0] MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_554_nl;
  wire[22:0] nl_MultLoop_acc_554_nl;
  wire[28:0] MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_553_nl;
  wire[22:0] nl_MultLoop_acc_553_nl;
  wire[28:0] MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_552_nl;
  wire[22:0] nl_MultLoop_acc_552_nl;
  wire[28:0] MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_551_nl;
  wire[22:0] nl_MultLoop_acc_551_nl;
  wire[28:0] MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_550_nl;
  wire[22:0] nl_MultLoop_acc_550_nl;
  wire[28:0] MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_549_nl;
  wire[22:0] nl_MultLoop_acc_549_nl;
  wire[28:0] MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_548_nl;
  wire[22:0] nl_MultLoop_acc_548_nl;
  wire[28:0] MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_547_nl;
  wire[22:0] nl_MultLoop_acc_547_nl;
  wire[28:0] MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_546_nl;
  wire[22:0] nl_MultLoop_acc_546_nl;
  wire[28:0] MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_545_nl;
  wire[22:0] nl_MultLoop_acc_545_nl;
  wire[28:0] MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_544_nl;
  wire[22:0] nl_MultLoop_acc_544_nl;
  wire[28:0] MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_543_nl;
  wire[22:0] nl_MultLoop_acc_543_nl;
  wire[28:0] MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_542_nl;
  wire[22:0] nl_MultLoop_acc_542_nl;
  wire[28:0] MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_541_nl;
  wire[22:0] nl_MultLoop_acc_541_nl;
  wire[28:0] MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_540_nl;
  wire[22:0] nl_MultLoop_acc_540_nl;
  wire[28:0] MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_539_nl;
  wire[22:0] nl_MultLoop_acc_539_nl;
  wire[28:0] MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_538_nl;
  wire[22:0] nl_MultLoop_acc_538_nl;
  wire[28:0] MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_537_nl;
  wire[22:0] nl_MultLoop_acc_537_nl;
  wire[28:0] MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_536_nl;
  wire[22:0] nl_MultLoop_acc_536_nl;
  wire[28:0] MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_535_nl;
  wire[22:0] nl_MultLoop_acc_535_nl;
  wire[28:0] MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_534_nl;
  wire[22:0] nl_MultLoop_acc_534_nl;
  wire[28:0] MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_533_nl;
  wire[22:0] nl_MultLoop_acc_533_nl;
  wire[28:0] MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_532_nl;
  wire[22:0] nl_MultLoop_acc_532_nl;
  wire[28:0] MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_531_nl;
  wire[22:0] nl_MultLoop_acc_531_nl;
  wire[28:0] MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_530_nl;
  wire[22:0] nl_MultLoop_acc_530_nl;
  wire[28:0] MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_529_nl;
  wire[22:0] nl_MultLoop_acc_529_nl;
  wire[28:0] MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_528_nl;
  wire[22:0] nl_MultLoop_acc_528_nl;
  wire[28:0] MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_527_nl;
  wire[22:0] nl_MultLoop_acc_527_nl;
  wire[28:0] MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_526_nl;
  wire[22:0] nl_MultLoop_acc_526_nl;
  wire[28:0] MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_525_nl;
  wire[22:0] nl_MultLoop_acc_525_nl;
  wire[28:0] MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_524_nl;
  wire[22:0] nl_MultLoop_acc_524_nl;
  wire[28:0] MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_523_nl;
  wire[22:0] nl_MultLoop_acc_523_nl;
  wire[28:0] MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_522_nl;
  wire[22:0] nl_MultLoop_acc_522_nl;
  wire[28:0] MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_521_nl;
  wire[22:0] nl_MultLoop_acc_521_nl;
  wire[28:0] MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_520_nl;
  wire[22:0] nl_MultLoop_acc_520_nl;
  wire[28:0] MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_519_nl;
  wire[22:0] nl_MultLoop_acc_519_nl;
  wire[28:0] MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_487_nl;
  wire[22:0] nl_MultLoop_acc_487_nl;
  wire[21:0] MultLoop_acc_455_nl;
  wire[22:0] nl_MultLoop_acc_455_nl;
  wire[10:0] MultLoop_acc_1283_nl;
  wire[11:0] nl_MultLoop_acc_1283_nl;
  wire[28:0] MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_454_nl;
  wire[22:0] nl_MultLoop_acc_454_nl;
  wire[28:0] MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_486_nl;
  wire[22:0] nl_MultLoop_acc_486_nl;
  wire[21:0] MultLoop_acc_453_nl;
  wire[22:0] nl_MultLoop_acc_453_nl;
  wire[28:0] MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_452_nl;
  wire[22:0] nl_MultLoop_acc_452_nl;
  wire[28:0] MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_451_nl;
  wire[22:0] nl_MultLoop_acc_451_nl;
  wire[28:0] MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_450_nl;
  wire[22:0] nl_MultLoop_acc_450_nl;
  wire[28:0] MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_449_nl;
  wire[22:0] nl_MultLoop_acc_449_nl;
  wire[28:0] MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_448_nl;
  wire[22:0] nl_MultLoop_acc_448_nl;
  wire[28:0] MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_447_nl;
  wire[22:0] nl_MultLoop_acc_447_nl;
  wire[28:0] MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_446_nl;
  wire[22:0] nl_MultLoop_acc_446_nl;
  wire[28:0] MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_445_nl;
  wire[22:0] nl_MultLoop_acc_445_nl;
  wire[28:0] MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_444_nl;
  wire[22:0] nl_MultLoop_acc_444_nl;
  wire[28:0] MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_443_nl;
  wire[22:0] nl_MultLoop_acc_443_nl;
  wire[28:0] MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_442_nl;
  wire[22:0] nl_MultLoop_acc_442_nl;
  wire[28:0] MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_441_nl;
  wire[22:0] nl_MultLoop_acc_441_nl;
  wire[28:0] MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_440_nl;
  wire[22:0] nl_MultLoop_acc_440_nl;
  wire[28:0] MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_439_nl;
  wire[22:0] nl_MultLoop_acc_439_nl;
  wire[28:0] MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_438_nl;
  wire[22:0] nl_MultLoop_acc_438_nl;
  wire[28:0] MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_437_nl;
  wire[22:0] nl_MultLoop_acc_437_nl;
  wire[28:0] MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_436_nl;
  wire[22:0] nl_MultLoop_acc_436_nl;
  wire[28:0] MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_435_nl;
  wire[22:0] nl_MultLoop_acc_435_nl;
  wire[28:0] MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_434_nl;
  wire[22:0] nl_MultLoop_acc_434_nl;
  wire[28:0] MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_433_nl;
  wire[22:0] nl_MultLoop_acc_433_nl;
  wire[28:0] MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_432_nl;
  wire[22:0] nl_MultLoop_acc_432_nl;
  wire[28:0] MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_431_nl;
  wire[22:0] nl_MultLoop_acc_431_nl;
  wire[28:0] MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_430_nl;
  wire[22:0] nl_MultLoop_acc_430_nl;
  wire[28:0] MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_429_nl;
  wire[22:0] nl_MultLoop_acc_429_nl;
  wire[28:0] MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_428_nl;
  wire[22:0] nl_MultLoop_acc_428_nl;
  wire[28:0] MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_427_nl;
  wire[22:0] nl_MultLoop_acc_427_nl;
  wire[28:0] MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_426_nl;
  wire[22:0] nl_MultLoop_acc_426_nl;
  wire[28:0] MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_425_nl;
  wire[22:0] nl_MultLoop_acc_425_nl;
  wire[28:0] MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_424_nl;
  wire[22:0] nl_MultLoop_acc_424_nl;
  wire[28:0] MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_423_nl;
  wire[22:0] nl_MultLoop_acc_423_nl;
  wire[28:0] MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_422_nl;
  wire[22:0] nl_MultLoop_acc_422_nl;
  wire[28:0] MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_421_nl;
  wire[22:0] nl_MultLoop_acc_421_nl;
  wire[28:0] MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_420_nl;
  wire[22:0] nl_MultLoop_acc_420_nl;
  wire[28:0] MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_419_nl;
  wire[22:0] nl_MultLoop_acc_419_nl;
  wire[28:0] MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_418_nl;
  wire[22:0] nl_MultLoop_acc_418_nl;
  wire[28:0] MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_417_nl;
  wire[22:0] nl_MultLoop_acc_417_nl;
  wire[28:0] MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_416_nl;
  wire[22:0] nl_MultLoop_acc_416_nl;
  wire[28:0] MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_415_nl;
  wire[22:0] nl_MultLoop_acc_415_nl;
  wire[28:0] MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_414_nl;
  wire[22:0] nl_MultLoop_acc_414_nl;
  wire[28:0] MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_413_nl;
  wire[22:0] nl_MultLoop_acc_413_nl;
  wire[28:0] MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_412_nl;
  wire[22:0] nl_MultLoop_acc_412_nl;
  wire[28:0] MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_411_nl;
  wire[22:0] nl_MultLoop_acc_411_nl;
  wire[28:0] MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_410_nl;
  wire[22:0] nl_MultLoop_acc_410_nl;
  wire[28:0] MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_409_nl;
  wire[22:0] nl_MultLoop_acc_409_nl;
  wire[28:0] MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_408_nl;
  wire[22:0] nl_MultLoop_acc_408_nl;
  wire[28:0] MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_407_nl;
  wire[22:0] nl_MultLoop_acc_407_nl;
  wire[28:0] MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_406_nl;
  wire[22:0] nl_MultLoop_acc_406_nl;
  wire[28:0] MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_405_nl;
  wire[22:0] nl_MultLoop_acc_405_nl;
  wire[28:0] MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_404_nl;
  wire[22:0] nl_MultLoop_acc_404_nl;
  wire[28:0] MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_403_nl;
  wire[22:0] nl_MultLoop_acc_403_nl;
  wire[28:0] MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_402_nl;
  wire[22:0] nl_MultLoop_acc_402_nl;
  wire[28:0] MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_401_nl;
  wire[22:0] nl_MultLoop_acc_401_nl;
  wire[28:0] MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_400_nl;
  wire[22:0] nl_MultLoop_acc_400_nl;
  wire[28:0] MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_399_nl;
  wire[22:0] nl_MultLoop_acc_399_nl;
  wire[28:0] MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_398_nl;
  wire[22:0] nl_MultLoop_acc_398_nl;
  wire[28:0] MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_397_nl;
  wire[22:0] nl_MultLoop_acc_397_nl;
  wire[28:0] MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_396_nl;
  wire[22:0] nl_MultLoop_acc_396_nl;
  wire[28:0] MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_395_nl;
  wire[22:0] nl_MultLoop_acc_395_nl;
  wire[28:0] MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_394_nl;
  wire[22:0] nl_MultLoop_acc_394_nl;
  wire[28:0] MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_393_nl;
  wire[22:0] nl_MultLoop_acc_393_nl;
  wire[28:0] MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_392_nl;
  wire[22:0] nl_MultLoop_acc_392_nl;
  wire[28:0] MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_360_nl;
  wire[22:0] nl_MultLoop_acc_360_nl;
  wire[21:0] MultLoop_acc_328_nl;
  wire[22:0] nl_MultLoop_acc_328_nl;
  wire[10:0] MultLoop_acc_1282_nl;
  wire[11:0] nl_MultLoop_acc_1282_nl;
  wire[28:0] MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_327_nl;
  wire[22:0] nl_MultLoop_acc_327_nl;
  wire[28:0] MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_359_nl;
  wire[22:0] nl_MultLoop_acc_359_nl;
  wire[21:0] MultLoop_acc_326_nl;
  wire[22:0] nl_MultLoop_acc_326_nl;
  wire[28:0] MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_325_nl;
  wire[22:0] nl_MultLoop_acc_325_nl;
  wire[28:0] MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_324_nl;
  wire[22:0] nl_MultLoop_acc_324_nl;
  wire[28:0] MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_323_nl;
  wire[22:0] nl_MultLoop_acc_323_nl;
  wire[28:0] MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_322_nl;
  wire[22:0] nl_MultLoop_acc_322_nl;
  wire[28:0] MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_321_nl;
  wire[22:0] nl_MultLoop_acc_321_nl;
  wire[28:0] MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_320_nl;
  wire[22:0] nl_MultLoop_acc_320_nl;
  wire[28:0] MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_319_nl;
  wire[22:0] nl_MultLoop_acc_319_nl;
  wire[28:0] MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_318_nl;
  wire[22:0] nl_MultLoop_acc_318_nl;
  wire[28:0] MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_317_nl;
  wire[22:0] nl_MultLoop_acc_317_nl;
  wire[28:0] MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_316_nl;
  wire[22:0] nl_MultLoop_acc_316_nl;
  wire[28:0] MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_315_nl;
  wire[22:0] nl_MultLoop_acc_315_nl;
  wire[28:0] MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_314_nl;
  wire[22:0] nl_MultLoop_acc_314_nl;
  wire[28:0] MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_313_nl;
  wire[22:0] nl_MultLoop_acc_313_nl;
  wire[28:0] MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_312_nl;
  wire[22:0] nl_MultLoop_acc_312_nl;
  wire[28:0] MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_311_nl;
  wire[22:0] nl_MultLoop_acc_311_nl;
  wire[28:0] MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_310_nl;
  wire[22:0] nl_MultLoop_acc_310_nl;
  wire[28:0] MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_309_nl;
  wire[22:0] nl_MultLoop_acc_309_nl;
  wire[28:0] MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_308_nl;
  wire[22:0] nl_MultLoop_acc_308_nl;
  wire[28:0] MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_307_nl;
  wire[22:0] nl_MultLoop_acc_307_nl;
  wire[28:0] MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_306_nl;
  wire[22:0] nl_MultLoop_acc_306_nl;
  wire[28:0] MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_305_nl;
  wire[22:0] nl_MultLoop_acc_305_nl;
  wire[28:0] MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_304_nl;
  wire[22:0] nl_MultLoop_acc_304_nl;
  wire[28:0] MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_303_nl;
  wire[22:0] nl_MultLoop_acc_303_nl;
  wire[28:0] MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_302_nl;
  wire[22:0] nl_MultLoop_acc_302_nl;
  wire[28:0] MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_301_nl;
  wire[22:0] nl_MultLoop_acc_301_nl;
  wire[28:0] MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_300_nl;
  wire[22:0] nl_MultLoop_acc_300_nl;
  wire[28:0] MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_299_nl;
  wire[22:0] nl_MultLoop_acc_299_nl;
  wire[28:0] MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_298_nl;
  wire[22:0] nl_MultLoop_acc_298_nl;
  wire[28:0] MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_297_nl;
  wire[22:0] nl_MultLoop_acc_297_nl;
  wire[28:0] MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_296_nl;
  wire[22:0] nl_MultLoop_acc_296_nl;
  wire[28:0] MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_295_nl;
  wire[22:0] nl_MultLoop_acc_295_nl;
  wire[28:0] MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_294_nl;
  wire[22:0] nl_MultLoop_acc_294_nl;
  wire[28:0] MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_293_nl;
  wire[22:0] nl_MultLoop_acc_293_nl;
  wire[28:0] MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_292_nl;
  wire[22:0] nl_MultLoop_acc_292_nl;
  wire[28:0] MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_291_nl;
  wire[22:0] nl_MultLoop_acc_291_nl;
  wire[28:0] MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_290_nl;
  wire[22:0] nl_MultLoop_acc_290_nl;
  wire[28:0] MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_289_nl;
  wire[22:0] nl_MultLoop_acc_289_nl;
  wire[28:0] MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_288_nl;
  wire[22:0] nl_MultLoop_acc_288_nl;
  wire[28:0] MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_287_nl;
  wire[22:0] nl_MultLoop_acc_287_nl;
  wire[28:0] MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_286_nl;
  wire[22:0] nl_MultLoop_acc_286_nl;
  wire[28:0] MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_285_nl;
  wire[22:0] nl_MultLoop_acc_285_nl;
  wire[28:0] MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_284_nl;
  wire[22:0] nl_MultLoop_acc_284_nl;
  wire[28:0] MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_283_nl;
  wire[22:0] nl_MultLoop_acc_283_nl;
  wire[28:0] MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_282_nl;
  wire[22:0] nl_MultLoop_acc_282_nl;
  wire[28:0] MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_281_nl;
  wire[22:0] nl_MultLoop_acc_281_nl;
  wire[28:0] MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_280_nl;
  wire[22:0] nl_MultLoop_acc_280_nl;
  wire[28:0] MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_279_nl;
  wire[22:0] nl_MultLoop_acc_279_nl;
  wire[28:0] MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_278_nl;
  wire[22:0] nl_MultLoop_acc_278_nl;
  wire[28:0] MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_277_nl;
  wire[22:0] nl_MultLoop_acc_277_nl;
  wire[28:0] MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_276_nl;
  wire[22:0] nl_MultLoop_acc_276_nl;
  wire[28:0] MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_275_nl;
  wire[22:0] nl_MultLoop_acc_275_nl;
  wire[28:0] MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_274_nl;
  wire[22:0] nl_MultLoop_acc_274_nl;
  wire[28:0] MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_273_nl;
  wire[22:0] nl_MultLoop_acc_273_nl;
  wire[28:0] MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_272_nl;
  wire[22:0] nl_MultLoop_acc_272_nl;
  wire[28:0] MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_271_nl;
  wire[22:0] nl_MultLoop_acc_271_nl;
  wire[28:0] MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_270_nl;
  wire[22:0] nl_MultLoop_acc_270_nl;
  wire[28:0] MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_269_nl;
  wire[22:0] nl_MultLoop_acc_269_nl;
  wire[28:0] MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_268_nl;
  wire[22:0] nl_MultLoop_acc_268_nl;
  wire[28:0] MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_267_nl;
  wire[22:0] nl_MultLoop_acc_267_nl;
  wire[28:0] MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_266_nl;
  wire[22:0] nl_MultLoop_acc_266_nl;
  wire[28:0] MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_265_nl;
  wire[22:0] nl_MultLoop_acc_265_nl;
  wire[28:0] MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_233_nl;
  wire[22:0] nl_MultLoop_acc_233_nl;
  wire[21:0] MultLoop_acc_201_nl;
  wire[22:0] nl_MultLoop_acc_201_nl;
  wire[10:0] MultLoop_acc_1281_nl;
  wire[11:0] nl_MultLoop_acc_1281_nl;
  wire[28:0] MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_200_nl;
  wire[22:0] nl_MultLoop_acc_200_nl;
  wire[28:0] MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_232_nl;
  wire[22:0] nl_MultLoop_acc_232_nl;
  wire[21:0] MultLoop_acc_199_nl;
  wire[22:0] nl_MultLoop_acc_199_nl;
  wire[28:0] MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_198_nl;
  wire[22:0] nl_MultLoop_acc_198_nl;
  wire[28:0] MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_197_nl;
  wire[22:0] nl_MultLoop_acc_197_nl;
  wire[28:0] MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_196_nl;
  wire[22:0] nl_MultLoop_acc_196_nl;
  wire[28:0] MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_195_nl;
  wire[22:0] nl_MultLoop_acc_195_nl;
  wire[28:0] MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_194_nl;
  wire[22:0] nl_MultLoop_acc_194_nl;
  wire[28:0] MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_193_nl;
  wire[22:0] nl_MultLoop_acc_193_nl;
  wire[28:0] MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_192_nl;
  wire[22:0] nl_MultLoop_acc_192_nl;
  wire[28:0] MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_191_nl;
  wire[22:0] nl_MultLoop_acc_191_nl;
  wire[28:0] MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_190_nl;
  wire[22:0] nl_MultLoop_acc_190_nl;
  wire[28:0] MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_189_nl;
  wire[22:0] nl_MultLoop_acc_189_nl;
  wire[28:0] MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_188_nl;
  wire[22:0] nl_MultLoop_acc_188_nl;
  wire[28:0] MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_187_nl;
  wire[22:0] nl_MultLoop_acc_187_nl;
  wire[28:0] MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_186_nl;
  wire[22:0] nl_MultLoop_acc_186_nl;
  wire[28:0] MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_185_nl;
  wire[22:0] nl_MultLoop_acc_185_nl;
  wire[28:0] MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_184_nl;
  wire[22:0] nl_MultLoop_acc_184_nl;
  wire[28:0] MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_183_nl;
  wire[22:0] nl_MultLoop_acc_183_nl;
  wire[28:0] MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_182_nl;
  wire[22:0] nl_MultLoop_acc_182_nl;
  wire[28:0] MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_181_nl;
  wire[22:0] nl_MultLoop_acc_181_nl;
  wire[28:0] MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_180_nl;
  wire[22:0] nl_MultLoop_acc_180_nl;
  wire[28:0] MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_179_nl;
  wire[22:0] nl_MultLoop_acc_179_nl;
  wire[28:0] MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_178_nl;
  wire[22:0] nl_MultLoop_acc_178_nl;
  wire[28:0] MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_177_nl;
  wire[22:0] nl_MultLoop_acc_177_nl;
  wire[28:0] MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_176_nl;
  wire[22:0] nl_MultLoop_acc_176_nl;
  wire[28:0] MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_175_nl;
  wire[22:0] nl_MultLoop_acc_175_nl;
  wire[28:0] MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_174_nl;
  wire[22:0] nl_MultLoop_acc_174_nl;
  wire[28:0] MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_173_nl;
  wire[22:0] nl_MultLoop_acc_173_nl;
  wire[28:0] MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_172_nl;
  wire[22:0] nl_MultLoop_acc_172_nl;
  wire[28:0] MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_171_nl;
  wire[22:0] nl_MultLoop_acc_171_nl;
  wire[28:0] MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_170_nl;
  wire[22:0] nl_MultLoop_acc_170_nl;
  wire[28:0] MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_169_nl;
  wire[22:0] nl_MultLoop_acc_169_nl;
  wire[28:0] MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_168_nl;
  wire[22:0] nl_MultLoop_acc_168_nl;
  wire[28:0] MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_167_nl;
  wire[22:0] nl_MultLoop_acc_167_nl;
  wire[28:0] MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_166_nl;
  wire[22:0] nl_MultLoop_acc_166_nl;
  wire[28:0] MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_165_nl;
  wire[22:0] nl_MultLoop_acc_165_nl;
  wire[28:0] MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_164_nl;
  wire[22:0] nl_MultLoop_acc_164_nl;
  wire[28:0] MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_163_nl;
  wire[22:0] nl_MultLoop_acc_163_nl;
  wire[28:0] MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_162_nl;
  wire[22:0] nl_MultLoop_acc_162_nl;
  wire[28:0] MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_161_nl;
  wire[22:0] nl_MultLoop_acc_161_nl;
  wire[28:0] MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_160_nl;
  wire[22:0] nl_MultLoop_acc_160_nl;
  wire[28:0] MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_159_nl;
  wire[22:0] nl_MultLoop_acc_159_nl;
  wire[28:0] MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_158_nl;
  wire[22:0] nl_MultLoop_acc_158_nl;
  wire[28:0] MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_157_nl;
  wire[22:0] nl_MultLoop_acc_157_nl;
  wire[28:0] MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_156_nl;
  wire[22:0] nl_MultLoop_acc_156_nl;
  wire[28:0] MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_155_nl;
  wire[22:0] nl_MultLoop_acc_155_nl;
  wire[28:0] MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_154_nl;
  wire[22:0] nl_MultLoop_acc_154_nl;
  wire[28:0] MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_153_nl;
  wire[22:0] nl_MultLoop_acc_153_nl;
  wire[28:0] MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_152_nl;
  wire[22:0] nl_MultLoop_acc_152_nl;
  wire[28:0] MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_151_nl;
  wire[22:0] nl_MultLoop_acc_151_nl;
  wire[28:0] MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_150_nl;
  wire[22:0] nl_MultLoop_acc_150_nl;
  wire[28:0] MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_149_nl;
  wire[22:0] nl_MultLoop_acc_149_nl;
  wire[28:0] MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_148_nl;
  wire[22:0] nl_MultLoop_acc_148_nl;
  wire[28:0] MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_147_nl;
  wire[22:0] nl_MultLoop_acc_147_nl;
  wire[28:0] MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_146_nl;
  wire[22:0] nl_MultLoop_acc_146_nl;
  wire[28:0] MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_145_nl;
  wire[22:0] nl_MultLoop_acc_145_nl;
  wire[28:0] MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_144_nl;
  wire[22:0] nl_MultLoop_acc_144_nl;
  wire[28:0] MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_143_nl;
  wire[22:0] nl_MultLoop_acc_143_nl;
  wire[28:0] MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_142_nl;
  wire[22:0] nl_MultLoop_acc_142_nl;
  wire[28:0] MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_141_nl;
  wire[22:0] nl_MultLoop_acc_141_nl;
  wire[28:0] MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_140_nl;
  wire[22:0] nl_MultLoop_acc_140_nl;
  wire[28:0] MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_139_nl;
  wire[22:0] nl_MultLoop_acc_139_nl;
  wire[28:0] MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_138_nl;
  wire[22:0] nl_MultLoop_acc_138_nl;
  wire[28:0] MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_122_nl;
  wire[22:0] nl_MultLoop_acc_122_nl;
  wire[21:0] MultLoop_acc_106_nl;
  wire[22:0] nl_MultLoop_acc_106_nl;
  wire[10:0] MultLoop_acc_1280_nl;
  wire[11:0] nl_MultLoop_acc_1280_nl;
  wire[28:0] MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_73_nl;
  wire[22:0] nl_MultLoop_acc_73_nl;
  wire[28:0] MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_105_nl;
  wire[22:0] nl_MultLoop_acc_105_nl;
  wire[21:0] MultLoop_acc_72_nl;
  wire[22:0] nl_MultLoop_acc_72_nl;
  wire[28:0] MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_71_nl;
  wire[22:0] nl_MultLoop_acc_71_nl;
  wire[28:0] MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_70_nl;
  wire[22:0] nl_MultLoop_acc_70_nl;
  wire[28:0] MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_69_nl;
  wire[22:0] nl_MultLoop_acc_69_nl;
  wire[28:0] MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_68_nl;
  wire[22:0] nl_MultLoop_acc_68_nl;
  wire[28:0] MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_67_nl;
  wire[22:0] nl_MultLoop_acc_67_nl;
  wire[28:0] MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_66_nl;
  wire[22:0] nl_MultLoop_acc_66_nl;
  wire[28:0] MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_65_nl;
  wire[22:0] nl_MultLoop_acc_65_nl;
  wire[28:0] MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_64_nl;
  wire[22:0] nl_MultLoop_acc_64_nl;
  wire[28:0] MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_63_nl;
  wire[22:0] nl_MultLoop_acc_63_nl;
  wire[28:0] MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_62_nl;
  wire[22:0] nl_MultLoop_acc_62_nl;
  wire[28:0] MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_61_nl;
  wire[22:0] nl_MultLoop_acc_61_nl;
  wire[28:0] MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_60_nl;
  wire[22:0] nl_MultLoop_acc_60_nl;
  wire[28:0] MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_59_nl;
  wire[22:0] nl_MultLoop_acc_59_nl;
  wire[28:0] MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_58_nl;
  wire[22:0] nl_MultLoop_acc_58_nl;
  wire[28:0] MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_57_nl;
  wire[22:0] nl_MultLoop_acc_57_nl;
  wire[28:0] MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_56_nl;
  wire[22:0] nl_MultLoop_acc_56_nl;
  wire[28:0] MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_55_nl;
  wire[22:0] nl_MultLoop_acc_55_nl;
  wire[28:0] MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_54_nl;
  wire[22:0] nl_MultLoop_acc_54_nl;
  wire[28:0] MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_53_nl;
  wire[22:0] nl_MultLoop_acc_53_nl;
  wire[28:0] MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_52_nl;
  wire[22:0] nl_MultLoop_acc_52_nl;
  wire[28:0] MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_51_nl;
  wire[22:0] nl_MultLoop_acc_51_nl;
  wire[28:0] MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_50_nl;
  wire[22:0] nl_MultLoop_acc_50_nl;
  wire[28:0] MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_49_nl;
  wire[22:0] nl_MultLoop_acc_49_nl;
  wire[28:0] MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_48_nl;
  wire[22:0] nl_MultLoop_acc_48_nl;
  wire[28:0] MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_47_nl;
  wire[22:0] nl_MultLoop_acc_47_nl;
  wire[28:0] MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_46_nl;
  wire[22:0] nl_MultLoop_acc_46_nl;
  wire[28:0] MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_45_nl;
  wire[22:0] nl_MultLoop_acc_45_nl;
  wire[28:0] MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_44_nl;
  wire[22:0] nl_MultLoop_acc_44_nl;
  wire[28:0] MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_43_nl;
  wire[22:0] nl_MultLoop_acc_43_nl;
  wire[28:0] MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_42_nl;
  wire[22:0] nl_MultLoop_acc_42_nl;
  wire[28:0] MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_41_nl;
  wire[22:0] nl_MultLoop_acc_41_nl;
  wire[28:0] MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_40_nl;
  wire[22:0] nl_MultLoop_acc_40_nl;
  wire[28:0] MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_39_nl;
  wire[22:0] nl_MultLoop_acc_39_nl;
  wire[28:0] MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_38_nl;
  wire[22:0] nl_MultLoop_acc_38_nl;
  wire[28:0] MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_37_nl;
  wire[22:0] nl_MultLoop_acc_37_nl;
  wire[28:0] MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_36_nl;
  wire[22:0] nl_MultLoop_acc_36_nl;
  wire[28:0] MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_35_nl;
  wire[22:0] nl_MultLoop_acc_35_nl;
  wire[28:0] MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_34_nl;
  wire[22:0] nl_MultLoop_acc_34_nl;
  wire[28:0] MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_33_nl;
  wire[22:0] nl_MultLoop_acc_33_nl;
  wire[28:0] MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_32_nl;
  wire[22:0] nl_MultLoop_acc_32_nl;
  wire[28:0] MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_31_nl;
  wire[22:0] nl_MultLoop_acc_31_nl;
  wire[28:0] MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_30_nl;
  wire[22:0] nl_MultLoop_acc_30_nl;
  wire[28:0] MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_29_nl;
  wire[22:0] nl_MultLoop_acc_29_nl;
  wire[28:0] MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_28_nl;
  wire[22:0] nl_MultLoop_acc_28_nl;
  wire[28:0] MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_27_nl;
  wire[22:0] nl_MultLoop_acc_27_nl;
  wire[28:0] MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_26_nl;
  wire[22:0] nl_MultLoop_acc_26_nl;
  wire[28:0] MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_25_nl;
  wire[22:0] nl_MultLoop_acc_25_nl;
  wire[28:0] MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_24_nl;
  wire[22:0] nl_MultLoop_acc_24_nl;
  wire[28:0] MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_23_nl;
  wire[22:0] nl_MultLoop_acc_23_nl;
  wire[28:0] MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_22_nl;
  wire[22:0] nl_MultLoop_acc_22_nl;
  wire[28:0] MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_21_nl;
  wire[22:0] nl_MultLoop_acc_21_nl;
  wire[28:0] MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_20_nl;
  wire[22:0] nl_MultLoop_acc_20_nl;
  wire[28:0] MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_19_nl;
  wire[22:0] nl_MultLoop_acc_19_nl;
  wire[28:0] MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_18_nl;
  wire[22:0] nl_MultLoop_acc_18_nl;
  wire[28:0] MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_17_nl;
  wire[22:0] nl_MultLoop_acc_17_nl;
  wire[28:0] MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_16_nl;
  wire[22:0] nl_MultLoop_acc_16_nl;
  wire[28:0] MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_15_nl;
  wire[22:0] nl_MultLoop_acc_15_nl;
  wire[28:0] MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_14_nl;
  wire[22:0] nl_MultLoop_acc_14_nl;
  wire[28:0] MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_13_nl;
  wire[22:0] nl_MultLoop_acc_13_nl;
  wire[28:0] MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_12_nl;
  wire[22:0] nl_MultLoop_acc_12_nl;
  wire[28:0] MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_11_nl;
  wire[22:0] nl_MultLoop_acc_11_nl;
  wire[28:0] MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[21:0] MultLoop_acc_1152_nl;
  wire[22:0] nl_MultLoop_acc_1152_nl;
  wire[21:0] MultLoop_acc_1150_nl;
  wire[22:0] nl_MultLoop_acc_1150_nl;
  wire[21:0] MultLoop_acc_1146_nl;
  wire[22:0] nl_MultLoop_acc_1146_nl;
  wire[21:0] MultLoop_acc_1145_nl;
  wire[22:0] nl_MultLoop_acc_1145_nl;
  wire[21:0] MultLoop_acc_1149_nl;
  wire[23:0] nl_MultLoop_acc_1149_nl;
  wire[21:0] MultLoop_acc_1151_nl;
  wire[24:0] nl_MultLoop_acc_1151_nl;
  wire[21:0] MultLoop_acc_1279_nl;
  wire[22:0] nl_MultLoop_acc_1279_nl;
  wire[21:0] MultLoop_acc_1277_nl;
  wire[22:0] nl_MultLoop_acc_1277_nl;
  wire[21:0] MultLoop_acc_1273_nl;
  wire[22:0] nl_MultLoop_acc_1273_nl;
  wire[21:0] MultLoop_acc_1272_nl;
  wire[22:0] nl_MultLoop_acc_1272_nl;
  wire[21:0] MultLoop_acc_1276_nl;
  wire[23:0] nl_MultLoop_acc_1276_nl;
  wire[21:0] MultLoop_acc_1278_nl;
  wire[24:0] nl_MultLoop_acc_1278_nl;
  wire[21:0] MultLoop_acc_1025_nl;
  wire[22:0] nl_MultLoop_acc_1025_nl;
  wire[21:0] MultLoop_acc_1023_nl;
  wire[22:0] nl_MultLoop_acc_1023_nl;
  wire[21:0] MultLoop_acc_1019_nl;
  wire[22:0] nl_MultLoop_acc_1019_nl;
  wire[21:0] MultLoop_acc_1018_nl;
  wire[22:0] nl_MultLoop_acc_1018_nl;
  wire[21:0] MultLoop_acc_1022_nl;
  wire[23:0] nl_MultLoop_acc_1022_nl;
  wire[21:0] MultLoop_acc_1024_nl;
  wire[24:0] nl_MultLoop_acc_1024_nl;
  wire[21:0] MultLoop_acc_nl;
  wire[22:0] nl_MultLoop_acc_nl;
  wire[21:0] MultLoop_acc_136_nl;
  wire[22:0] nl_MultLoop_acc_136_nl;
  wire[21:0] MultLoop_acc_134_nl;
  wire[22:0] nl_MultLoop_acc_134_nl;
  wire[21:0] MultLoop_acc_129_nl;
  wire[22:0] nl_MultLoop_acc_129_nl;
  wire[21:0] MultLoop_acc_133_nl;
  wire[23:0] nl_MultLoop_acc_133_nl;
  wire[21:0] MultLoop_acc_135_nl;
  wire[24:0] nl_MultLoop_acc_135_nl;
  wire[21:0] MultLoop_acc_898_nl;
  wire[22:0] nl_MultLoop_acc_898_nl;
  wire[21:0] MultLoop_acc_896_nl;
  wire[22:0] nl_MultLoop_acc_896_nl;
  wire[21:0] MultLoop_acc_892_nl;
  wire[22:0] nl_MultLoop_acc_892_nl;
  wire[21:0] MultLoop_acc_891_nl;
  wire[22:0] nl_MultLoop_acc_891_nl;
  wire[21:0] MultLoop_acc_895_nl;
  wire[23:0] nl_MultLoop_acc_895_nl;
  wire[21:0] MultLoop_acc_897_nl;
  wire[24:0] nl_MultLoop_acc_897_nl;
  wire[21:0] MultLoop_acc_263_nl;
  wire[22:0] nl_MultLoop_acc_263_nl;
  wire[21:0] MultLoop_acc_261_nl;
  wire[22:0] nl_MultLoop_acc_261_nl;
  wire[21:0] MultLoop_acc_257_nl;
  wire[22:0] nl_MultLoop_acc_257_nl;
  wire[21:0] MultLoop_acc_256_nl;
  wire[22:0] nl_MultLoop_acc_256_nl;
  wire[21:0] MultLoop_acc_260_nl;
  wire[23:0] nl_MultLoop_acc_260_nl;
  wire[21:0] MultLoop_acc_262_nl;
  wire[24:0] nl_MultLoop_acc_262_nl;
  wire[21:0] MultLoop_acc_771_nl;
  wire[22:0] nl_MultLoop_acc_771_nl;
  wire[21:0] MultLoop_acc_769_nl;
  wire[22:0] nl_MultLoop_acc_769_nl;
  wire[21:0] MultLoop_acc_765_nl;
  wire[22:0] nl_MultLoop_acc_765_nl;
  wire[21:0] MultLoop_acc_764_nl;
  wire[22:0] nl_MultLoop_acc_764_nl;
  wire[21:0] MultLoop_acc_768_nl;
  wire[23:0] nl_MultLoop_acc_768_nl;
  wire[21:0] MultLoop_acc_770_nl;
  wire[24:0] nl_MultLoop_acc_770_nl;
  wire[21:0] MultLoop_acc_390_nl;
  wire[22:0] nl_MultLoop_acc_390_nl;
  wire[21:0] MultLoop_acc_388_nl;
  wire[22:0] nl_MultLoop_acc_388_nl;
  wire[21:0] MultLoop_acc_384_nl;
  wire[22:0] nl_MultLoop_acc_384_nl;
  wire[21:0] MultLoop_acc_383_nl;
  wire[22:0] nl_MultLoop_acc_383_nl;
  wire[21:0] MultLoop_acc_387_nl;
  wire[23:0] nl_MultLoop_acc_387_nl;
  wire[21:0] MultLoop_acc_389_nl;
  wire[24:0] nl_MultLoop_acc_389_nl;
  wire[21:0] MultLoop_acc_644_nl;
  wire[22:0] nl_MultLoop_acc_644_nl;
  wire[21:0] MultLoop_acc_642_nl;
  wire[22:0] nl_MultLoop_acc_642_nl;
  wire[21:0] MultLoop_acc_638_nl;
  wire[22:0] nl_MultLoop_acc_638_nl;
  wire[21:0] MultLoop_acc_637_nl;
  wire[22:0] nl_MultLoop_acc_637_nl;
  wire[21:0] MultLoop_acc_641_nl;
  wire[23:0] nl_MultLoop_acc_641_nl;
  wire[21:0] MultLoop_acc_643_nl;
  wire[24:0] nl_MultLoop_acc_643_nl;
  wire[21:0] MultLoop_acc_517_nl;
  wire[22:0] nl_MultLoop_acc_517_nl;
  wire[21:0] MultLoop_acc_515_nl;
  wire[22:0] nl_MultLoop_acc_515_nl;
  wire[21:0] MultLoop_acc_511_nl;
  wire[22:0] nl_MultLoop_acc_511_nl;
  wire[21:0] MultLoop_acc_510_nl;
  wire[22:0] nl_MultLoop_acc_510_nl;
  wire[21:0] MultLoop_acc_514_nl;
  wire[23:0] nl_MultLoop_acc_514_nl;
  wire[21:0] MultLoop_acc_516_nl;
  wire[24:0] nl_MultLoop_acc_516_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[28:0] MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[28:0] MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[21:0] AccumDotWidth_acc_2271_nl;
  wire[23:0] nl_AccumDotWidth_acc_2271_nl;
  wire[9:0] AccumDotWidth_acc_2400_nl;
  wire[10:0] nl_AccumDotWidth_acc_2400_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2270_nl;
  wire[23:0] nl_AccumDotWidth_acc_2270_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2269_nl;
  wire[23:0] nl_AccumDotWidth_acc_2269_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2260_nl;
  wire[23:0] nl_AccumDotWidth_acc_2260_nl;
  wire[9:0] AccumDotWidth_acc_2399_nl;
  wire[10:0] nl_AccumDotWidth_acc_2399_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2259_nl;
  wire[23:0] nl_AccumDotWidth_acc_2259_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2258_nl;
  wire[23:0] nl_AccumDotWidth_acc_2258_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2249_nl;
  wire[23:0] nl_AccumDotWidth_acc_2249_nl;
  wire[9:0] AccumDotWidth_acc_2398_nl;
  wire[10:0] nl_AccumDotWidth_acc_2398_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2248_nl;
  wire[23:0] nl_AccumDotWidth_acc_2248_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2247_nl;
  wire[23:0] nl_AccumDotWidth_acc_2247_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2238_nl;
  wire[23:0] nl_AccumDotWidth_acc_2238_nl;
  wire[9:0] AccumDotWidth_acc_2397_nl;
  wire[10:0] nl_AccumDotWidth_acc_2397_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2237_nl;
  wire[23:0] nl_AccumDotWidth_acc_2237_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2236_nl;
  wire[23:0] nl_AccumDotWidth_acc_2236_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2227_nl;
  wire[23:0] nl_AccumDotWidth_acc_2227_nl;
  wire[9:0] AccumDotWidth_acc_2396_nl;
  wire[10:0] nl_AccumDotWidth_acc_2396_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2226_nl;
  wire[23:0] nl_AccumDotWidth_acc_2226_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2225_nl;
  wire[23:0] nl_AccumDotWidth_acc_2225_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2216_nl;
  wire[23:0] nl_AccumDotWidth_acc_2216_nl;
  wire[9:0] AccumDotWidth_acc_2395_nl;
  wire[10:0] nl_AccumDotWidth_acc_2395_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2215_nl;
  wire[23:0] nl_AccumDotWidth_acc_2215_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2214_nl;
  wire[23:0] nl_AccumDotWidth_acc_2214_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2205_nl;
  wire[23:0] nl_AccumDotWidth_acc_2205_nl;
  wire[9:0] AccumDotWidth_acc_2394_nl;
  wire[10:0] nl_AccumDotWidth_acc_2394_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2204_nl;
  wire[23:0] nl_AccumDotWidth_acc_2204_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2203_nl;
  wire[23:0] nl_AccumDotWidth_acc_2203_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2194_nl;
  wire[23:0] nl_AccumDotWidth_acc_2194_nl;
  wire[9:0] AccumDotWidth_acc_2393_nl;
  wire[10:0] nl_AccumDotWidth_acc_2393_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2193_nl;
  wire[23:0] nl_AccumDotWidth_acc_2193_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2192_nl;
  wire[23:0] nl_AccumDotWidth_acc_2192_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2182_nl;
  wire[24:0] nl_AccumDotWidth_acc_2182_nl;
  wire[9:0] AccumDotWidth_acc_2392_nl;
  wire[10:0] nl_AccumDotWidth_acc_2392_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2181_nl;
  wire[23:0] nl_AccumDotWidth_acc_2181_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2179_nl;
  wire[23:0] nl_AccumDotWidth_acc_2179_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2165_nl;
  wire[24:0] nl_AccumDotWidth_acc_2165_nl;
  wire[9:0] AccumDotWidth_acc_2391_nl;
  wire[10:0] nl_AccumDotWidth_acc_2391_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2164_nl;
  wire[23:0] nl_AccumDotWidth_acc_2164_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2162_nl;
  wire[23:0] nl_AccumDotWidth_acc_2162_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2148_nl;
  wire[24:0] nl_AccumDotWidth_acc_2148_nl;
  wire[9:0] AccumDotWidth_acc_2390_nl;
  wire[10:0] nl_AccumDotWidth_acc_2390_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2147_nl;
  wire[23:0] nl_AccumDotWidth_acc_2147_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2145_nl;
  wire[23:0] nl_AccumDotWidth_acc_2145_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2131_nl;
  wire[24:0] nl_AccumDotWidth_acc_2131_nl;
  wire[9:0] AccumDotWidth_acc_2389_nl;
  wire[10:0] nl_AccumDotWidth_acc_2389_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2130_nl;
  wire[23:0] nl_AccumDotWidth_acc_2130_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2128_nl;
  wire[23:0] nl_AccumDotWidth_acc_2128_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2114_nl;
  wire[24:0] nl_AccumDotWidth_acc_2114_nl;
  wire[9:0] AccumDotWidth_acc_2388_nl;
  wire[10:0] nl_AccumDotWidth_acc_2388_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2113_nl;
  wire[23:0] nl_AccumDotWidth_acc_2113_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2111_nl;
  wire[23:0] nl_AccumDotWidth_acc_2111_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2097_nl;
  wire[24:0] nl_AccumDotWidth_acc_2097_nl;
  wire[9:0] AccumDotWidth_acc_2387_nl;
  wire[10:0] nl_AccumDotWidth_acc_2387_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2096_nl;
  wire[23:0] nl_AccumDotWidth_acc_2096_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2094_nl;
  wire[23:0] nl_AccumDotWidth_acc_2094_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2080_nl;
  wire[24:0] nl_AccumDotWidth_acc_2080_nl;
  wire[9:0] AccumDotWidth_acc_2386_nl;
  wire[10:0] nl_AccumDotWidth_acc_2386_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2079_nl;
  wire[23:0] nl_AccumDotWidth_acc_2079_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2077_nl;
  wire[23:0] nl_AccumDotWidth_acc_2077_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2063_nl;
  wire[24:0] nl_AccumDotWidth_acc_2063_nl;
  wire[9:0] AccumDotWidth_acc_2385_nl;
  wire[10:0] nl_AccumDotWidth_acc_2385_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2062_nl;
  wire[23:0] nl_AccumDotWidth_acc_2062_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2060_nl;
  wire[23:0] nl_AccumDotWidth_acc_2060_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2046_nl;
  wire[24:0] nl_AccumDotWidth_acc_2046_nl;
  wire[9:0] AccumDotWidth_acc_2384_nl;
  wire[10:0] nl_AccumDotWidth_acc_2384_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2045_nl;
  wire[23:0] nl_AccumDotWidth_acc_2045_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2043_nl;
  wire[23:0] nl_AccumDotWidth_acc_2043_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2029_nl;
  wire[24:0] nl_AccumDotWidth_acc_2029_nl;
  wire[9:0] AccumDotWidth_acc_2383_nl;
  wire[10:0] nl_AccumDotWidth_acc_2383_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2028_nl;
  wire[23:0] nl_AccumDotWidth_acc_2028_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2026_nl;
  wire[23:0] nl_AccumDotWidth_acc_2026_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2012_nl;
  wire[24:0] nl_AccumDotWidth_acc_2012_nl;
  wire[9:0] AccumDotWidth_acc_2382_nl;
  wire[10:0] nl_AccumDotWidth_acc_2382_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2011_nl;
  wire[23:0] nl_AccumDotWidth_acc_2011_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_2009_nl;
  wire[23:0] nl_AccumDotWidth_acc_2009_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1995_nl;
  wire[24:0] nl_AccumDotWidth_acc_1995_nl;
  wire[9:0] AccumDotWidth_acc_2381_nl;
  wire[10:0] nl_AccumDotWidth_acc_2381_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1994_nl;
  wire[23:0] nl_AccumDotWidth_acc_1994_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1992_nl;
  wire[23:0] nl_AccumDotWidth_acc_1992_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1978_nl;
  wire[24:0] nl_AccumDotWidth_acc_1978_nl;
  wire[9:0] AccumDotWidth_acc_2380_nl;
  wire[10:0] nl_AccumDotWidth_acc_2380_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1977_nl;
  wire[23:0] nl_AccumDotWidth_acc_1977_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1975_nl;
  wire[23:0] nl_AccumDotWidth_acc_1975_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1961_nl;
  wire[24:0] nl_AccumDotWidth_acc_1961_nl;
  wire[9:0] AccumDotWidth_acc_2379_nl;
  wire[10:0] nl_AccumDotWidth_acc_2379_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1960_nl;
  wire[23:0] nl_AccumDotWidth_acc_1960_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1958_nl;
  wire[23:0] nl_AccumDotWidth_acc_1958_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1944_nl;
  wire[24:0] nl_AccumDotWidth_acc_1944_nl;
  wire[9:0] AccumDotWidth_acc_2378_nl;
  wire[10:0] nl_AccumDotWidth_acc_2378_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1943_nl;
  wire[23:0] nl_AccumDotWidth_acc_1943_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1941_nl;
  wire[23:0] nl_AccumDotWidth_acc_1941_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1927_nl;
  wire[24:0] nl_AccumDotWidth_acc_1927_nl;
  wire[9:0] AccumDotWidth_acc_2377_nl;
  wire[10:0] nl_AccumDotWidth_acc_2377_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1926_nl;
  wire[23:0] nl_AccumDotWidth_acc_1926_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1924_nl;
  wire[23:0] nl_AccumDotWidth_acc_1924_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1911_nl;
  wire[23:0] nl_AccumDotWidth_acc_1911_nl;
  wire[9:0] AccumDotWidth_acc_2376_nl;
  wire[10:0] nl_AccumDotWidth_acc_2376_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1910_nl;
  wire[23:0] nl_AccumDotWidth_acc_1910_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1909_nl;
  wire[23:0] nl_AccumDotWidth_acc_1909_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1900_nl;
  wire[23:0] nl_AccumDotWidth_acc_1900_nl;
  wire[9:0] AccumDotWidth_acc_2375_nl;
  wire[10:0] nl_AccumDotWidth_acc_2375_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1899_nl;
  wire[23:0] nl_AccumDotWidth_acc_1899_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1898_nl;
  wire[23:0] nl_AccumDotWidth_acc_1898_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1889_nl;
  wire[23:0] nl_AccumDotWidth_acc_1889_nl;
  wire[9:0] AccumDotWidth_acc_2374_nl;
  wire[10:0] nl_AccumDotWidth_acc_2374_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1888_nl;
  wire[23:0] nl_AccumDotWidth_acc_1888_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1887_nl;
  wire[23:0] nl_AccumDotWidth_acc_1887_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1878_nl;
  wire[23:0] nl_AccumDotWidth_acc_1878_nl;
  wire[9:0] AccumDotWidth_acc_2373_nl;
  wire[10:0] nl_AccumDotWidth_acc_2373_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1877_nl;
  wire[23:0] nl_AccumDotWidth_acc_1877_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1876_nl;
  wire[23:0] nl_AccumDotWidth_acc_1876_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1867_nl;
  wire[23:0] nl_AccumDotWidth_acc_1867_nl;
  wire[9:0] AccumDotWidth_acc_2372_nl;
  wire[10:0] nl_AccumDotWidth_acc_2372_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1866_nl;
  wire[23:0] nl_AccumDotWidth_acc_1866_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1865_nl;
  wire[23:0] nl_AccumDotWidth_acc_1865_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1856_nl;
  wire[23:0] nl_AccumDotWidth_acc_1856_nl;
  wire[9:0] AccumDotWidth_acc_2371_nl;
  wire[10:0] nl_AccumDotWidth_acc_2371_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1855_nl;
  wire[23:0] nl_AccumDotWidth_acc_1855_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1854_nl;
  wire[23:0] nl_AccumDotWidth_acc_1854_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1845_nl;
  wire[23:0] nl_AccumDotWidth_acc_1845_nl;
  wire[9:0] AccumDotWidth_acc_2370_nl;
  wire[10:0] nl_AccumDotWidth_acc_2370_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1844_nl;
  wire[23:0] nl_AccumDotWidth_acc_1844_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1843_nl;
  wire[23:0] nl_AccumDotWidth_acc_1843_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1834_nl;
  wire[23:0] nl_AccumDotWidth_acc_1834_nl;
  wire[9:0] AccumDotWidth_acc_2369_nl;
  wire[10:0] nl_AccumDotWidth_acc_2369_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1833_nl;
  wire[23:0] nl_AccumDotWidth_acc_1833_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1832_nl;
  wire[23:0] nl_AccumDotWidth_acc_1832_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1822_nl;
  wire[24:0] nl_AccumDotWidth_acc_1822_nl;
  wire[9:0] AccumDotWidth_acc_2368_nl;
  wire[10:0] nl_AccumDotWidth_acc_2368_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1821_nl;
  wire[23:0] nl_AccumDotWidth_acc_1821_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1819_nl;
  wire[23:0] nl_AccumDotWidth_acc_1819_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1805_nl;
  wire[24:0] nl_AccumDotWidth_acc_1805_nl;
  wire[9:0] AccumDotWidth_acc_2367_nl;
  wire[10:0] nl_AccumDotWidth_acc_2367_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1804_nl;
  wire[23:0] nl_AccumDotWidth_acc_1804_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1802_nl;
  wire[23:0] nl_AccumDotWidth_acc_1802_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1788_nl;
  wire[24:0] nl_AccumDotWidth_acc_1788_nl;
  wire[9:0] AccumDotWidth_acc_2366_nl;
  wire[10:0] nl_AccumDotWidth_acc_2366_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1787_nl;
  wire[23:0] nl_AccumDotWidth_acc_1787_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1785_nl;
  wire[23:0] nl_AccumDotWidth_acc_1785_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1771_nl;
  wire[24:0] nl_AccumDotWidth_acc_1771_nl;
  wire[9:0] AccumDotWidth_acc_2365_nl;
  wire[10:0] nl_AccumDotWidth_acc_2365_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1770_nl;
  wire[23:0] nl_AccumDotWidth_acc_1770_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1768_nl;
  wire[23:0] nl_AccumDotWidth_acc_1768_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1754_nl;
  wire[24:0] nl_AccumDotWidth_acc_1754_nl;
  wire[9:0] AccumDotWidth_acc_2364_nl;
  wire[10:0] nl_AccumDotWidth_acc_2364_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1753_nl;
  wire[23:0] nl_AccumDotWidth_acc_1753_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1751_nl;
  wire[23:0] nl_AccumDotWidth_acc_1751_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1737_nl;
  wire[24:0] nl_AccumDotWidth_acc_1737_nl;
  wire[9:0] AccumDotWidth_acc_2363_nl;
  wire[10:0] nl_AccumDotWidth_acc_2363_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1736_nl;
  wire[23:0] nl_AccumDotWidth_acc_1736_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1734_nl;
  wire[23:0] nl_AccumDotWidth_acc_1734_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1720_nl;
  wire[24:0] nl_AccumDotWidth_acc_1720_nl;
  wire[9:0] AccumDotWidth_acc_2362_nl;
  wire[10:0] nl_AccumDotWidth_acc_2362_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1719_nl;
  wire[23:0] nl_AccumDotWidth_acc_1719_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1717_nl;
  wire[23:0] nl_AccumDotWidth_acc_1717_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1703_nl;
  wire[24:0] nl_AccumDotWidth_acc_1703_nl;
  wire[9:0] AccumDotWidth_acc_2361_nl;
  wire[10:0] nl_AccumDotWidth_acc_2361_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1702_nl;
  wire[23:0] nl_AccumDotWidth_acc_1702_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1700_nl;
  wire[23:0] nl_AccumDotWidth_acc_1700_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1686_nl;
  wire[24:0] nl_AccumDotWidth_acc_1686_nl;
  wire[21:0] AccumDotWidth_acc_1681_nl;
  wire[23:0] nl_AccumDotWidth_acc_1681_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1685_nl;
  wire[24:0] nl_AccumDotWidth_acc_1685_nl;
  wire[21:0] AccumDotWidth_acc_1679_nl;
  wire[23:0] nl_AccumDotWidth_acc_1679_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1683_nl;
  wire[23:0] nl_AccumDotWidth_acc_1683_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1678_nl;
  wire[23:0] nl_AccumDotWidth_acc_1678_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1677_nl;
  wire[23:0] nl_AccumDotWidth_acc_1677_nl;
  wire[9:0] AccumDotWidth_acc_2360_nl;
  wire[10:0] nl_AccumDotWidth_acc_2360_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1660_nl;
  wire[24:0] nl_AccumDotWidth_acc_1660_nl;
  wire[21:0] AccumDotWidth_acc_1655_nl;
  wire[23:0] nl_AccumDotWidth_acc_1655_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1659_nl;
  wire[24:0] nl_AccumDotWidth_acc_1659_nl;
  wire[21:0] AccumDotWidth_acc_1653_nl;
  wire[23:0] nl_AccumDotWidth_acc_1653_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1657_nl;
  wire[23:0] nl_AccumDotWidth_acc_1657_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1652_nl;
  wire[23:0] nl_AccumDotWidth_acc_1652_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1651_nl;
  wire[23:0] nl_AccumDotWidth_acc_1651_nl;
  wire[9:0] AccumDotWidth_acc_2359_nl;
  wire[10:0] nl_AccumDotWidth_acc_2359_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1634_nl;
  wire[24:0] nl_AccumDotWidth_acc_1634_nl;
  wire[21:0] AccumDotWidth_acc_1629_nl;
  wire[23:0] nl_AccumDotWidth_acc_1629_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1633_nl;
  wire[24:0] nl_AccumDotWidth_acc_1633_nl;
  wire[21:0] AccumDotWidth_acc_1627_nl;
  wire[23:0] nl_AccumDotWidth_acc_1627_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1631_nl;
  wire[23:0] nl_AccumDotWidth_acc_1631_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1626_nl;
  wire[23:0] nl_AccumDotWidth_acc_1626_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1625_nl;
  wire[23:0] nl_AccumDotWidth_acc_1625_nl;
  wire[9:0] AccumDotWidth_acc_2358_nl;
  wire[10:0] nl_AccumDotWidth_acc_2358_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1608_nl;
  wire[24:0] nl_AccumDotWidth_acc_1608_nl;
  wire[21:0] AccumDotWidth_acc_1603_nl;
  wire[23:0] nl_AccumDotWidth_acc_1603_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1607_nl;
  wire[24:0] nl_AccumDotWidth_acc_1607_nl;
  wire[21:0] AccumDotWidth_acc_1601_nl;
  wire[23:0] nl_AccumDotWidth_acc_1601_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1605_nl;
  wire[23:0] nl_AccumDotWidth_acc_1605_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1600_nl;
  wire[23:0] nl_AccumDotWidth_acc_1600_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1599_nl;
  wire[23:0] nl_AccumDotWidth_acc_1599_nl;
  wire[9:0] AccumDotWidth_acc_2357_nl;
  wire[10:0] nl_AccumDotWidth_acc_2357_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1582_nl;
  wire[24:0] nl_AccumDotWidth_acc_1582_nl;
  wire[21:0] AccumDotWidth_acc_1577_nl;
  wire[23:0] nl_AccumDotWidth_acc_1577_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1581_nl;
  wire[24:0] nl_AccumDotWidth_acc_1581_nl;
  wire[21:0] AccumDotWidth_acc_1575_nl;
  wire[23:0] nl_AccumDotWidth_acc_1575_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1579_nl;
  wire[23:0] nl_AccumDotWidth_acc_1579_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1574_nl;
  wire[23:0] nl_AccumDotWidth_acc_1574_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1573_nl;
  wire[23:0] nl_AccumDotWidth_acc_1573_nl;
  wire[9:0] AccumDotWidth_acc_2356_nl;
  wire[10:0] nl_AccumDotWidth_acc_2356_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1556_nl;
  wire[24:0] nl_AccumDotWidth_acc_1556_nl;
  wire[21:0] AccumDotWidth_acc_1551_nl;
  wire[23:0] nl_AccumDotWidth_acc_1551_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1555_nl;
  wire[24:0] nl_AccumDotWidth_acc_1555_nl;
  wire[21:0] AccumDotWidth_acc_1549_nl;
  wire[23:0] nl_AccumDotWidth_acc_1549_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1553_nl;
  wire[23:0] nl_AccumDotWidth_acc_1553_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1548_nl;
  wire[23:0] nl_AccumDotWidth_acc_1548_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1547_nl;
  wire[23:0] nl_AccumDotWidth_acc_1547_nl;
  wire[9:0] AccumDotWidth_acc_2355_nl;
  wire[10:0] nl_AccumDotWidth_acc_2355_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1530_nl;
  wire[24:0] nl_AccumDotWidth_acc_1530_nl;
  wire[21:0] AccumDotWidth_acc_1525_nl;
  wire[23:0] nl_AccumDotWidth_acc_1525_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1529_nl;
  wire[24:0] nl_AccumDotWidth_acc_1529_nl;
  wire[21:0] AccumDotWidth_acc_1523_nl;
  wire[23:0] nl_AccumDotWidth_acc_1523_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1527_nl;
  wire[23:0] nl_AccumDotWidth_acc_1527_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1522_nl;
  wire[23:0] nl_AccumDotWidth_acc_1522_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1521_nl;
  wire[23:0] nl_AccumDotWidth_acc_1521_nl;
  wire[9:0] AccumDotWidth_acc_2354_nl;
  wire[10:0] nl_AccumDotWidth_acc_2354_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1504_nl;
  wire[24:0] nl_AccumDotWidth_acc_1504_nl;
  wire[21:0] AccumDotWidth_acc_1499_nl;
  wire[23:0] nl_AccumDotWidth_acc_1499_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1503_nl;
  wire[24:0] nl_AccumDotWidth_acc_1503_nl;
  wire[21:0] AccumDotWidth_acc_1497_nl;
  wire[23:0] nl_AccumDotWidth_acc_1497_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1501_nl;
  wire[23:0] nl_AccumDotWidth_acc_1501_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1496_nl;
  wire[23:0] nl_AccumDotWidth_acc_1496_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1495_nl;
  wire[23:0] nl_AccumDotWidth_acc_1495_nl;
  wire[9:0] AccumDotWidth_acc_2353_nl;
  wire[10:0] nl_AccumDotWidth_acc_2353_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1478_nl;
  wire[24:0] nl_AccumDotWidth_acc_1478_nl;
  wire[21:0] AccumDotWidth_acc_1473_nl;
  wire[23:0] nl_AccumDotWidth_acc_1473_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1477_nl;
  wire[24:0] nl_AccumDotWidth_acc_1477_nl;
  wire[21:0] AccumDotWidth_acc_1471_nl;
  wire[23:0] nl_AccumDotWidth_acc_1471_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1475_nl;
  wire[23:0] nl_AccumDotWidth_acc_1475_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1470_nl;
  wire[23:0] nl_AccumDotWidth_acc_1470_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1469_nl;
  wire[23:0] nl_AccumDotWidth_acc_1469_nl;
  wire[9:0] AccumDotWidth_acc_2352_nl;
  wire[10:0] nl_AccumDotWidth_acc_2352_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1452_nl;
  wire[24:0] nl_AccumDotWidth_acc_1452_nl;
  wire[21:0] AccumDotWidth_acc_1447_nl;
  wire[23:0] nl_AccumDotWidth_acc_1447_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1451_nl;
  wire[24:0] nl_AccumDotWidth_acc_1451_nl;
  wire[21:0] AccumDotWidth_acc_1445_nl;
  wire[23:0] nl_AccumDotWidth_acc_1445_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1449_nl;
  wire[23:0] nl_AccumDotWidth_acc_1449_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1444_nl;
  wire[23:0] nl_AccumDotWidth_acc_1444_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1443_nl;
  wire[23:0] nl_AccumDotWidth_acc_1443_nl;
  wire[9:0] AccumDotWidth_acc_2351_nl;
  wire[10:0] nl_AccumDotWidth_acc_2351_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1426_nl;
  wire[24:0] nl_AccumDotWidth_acc_1426_nl;
  wire[21:0] AccumDotWidth_acc_1421_nl;
  wire[23:0] nl_AccumDotWidth_acc_1421_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1425_nl;
  wire[24:0] nl_AccumDotWidth_acc_1425_nl;
  wire[21:0] AccumDotWidth_acc_1419_nl;
  wire[23:0] nl_AccumDotWidth_acc_1419_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1423_nl;
  wire[23:0] nl_AccumDotWidth_acc_1423_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1418_nl;
  wire[23:0] nl_AccumDotWidth_acc_1418_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1417_nl;
  wire[23:0] nl_AccumDotWidth_acc_1417_nl;
  wire[9:0] AccumDotWidth_acc_2350_nl;
  wire[10:0] nl_AccumDotWidth_acc_2350_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1400_nl;
  wire[24:0] nl_AccumDotWidth_acc_1400_nl;
  wire[21:0] AccumDotWidth_acc_1395_nl;
  wire[23:0] nl_AccumDotWidth_acc_1395_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1399_nl;
  wire[24:0] nl_AccumDotWidth_acc_1399_nl;
  wire[21:0] AccumDotWidth_acc_1393_nl;
  wire[23:0] nl_AccumDotWidth_acc_1393_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1397_nl;
  wire[23:0] nl_AccumDotWidth_acc_1397_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1392_nl;
  wire[23:0] nl_AccumDotWidth_acc_1392_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1391_nl;
  wire[23:0] nl_AccumDotWidth_acc_1391_nl;
  wire[9:0] AccumDotWidth_acc_2349_nl;
  wire[10:0] nl_AccumDotWidth_acc_2349_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1374_nl;
  wire[24:0] nl_AccumDotWidth_acc_1374_nl;
  wire[21:0] AccumDotWidth_acc_1369_nl;
  wire[23:0] nl_AccumDotWidth_acc_1369_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1373_nl;
  wire[24:0] nl_AccumDotWidth_acc_1373_nl;
  wire[21:0] AccumDotWidth_acc_1367_nl;
  wire[23:0] nl_AccumDotWidth_acc_1367_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1371_nl;
  wire[23:0] nl_AccumDotWidth_acc_1371_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1366_nl;
  wire[23:0] nl_AccumDotWidth_acc_1366_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1365_nl;
  wire[23:0] nl_AccumDotWidth_acc_1365_nl;
  wire[9:0] AccumDotWidth_acc_2348_nl;
  wire[10:0] nl_AccumDotWidth_acc_2348_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1348_nl;
  wire[24:0] nl_AccumDotWidth_acc_1348_nl;
  wire[21:0] AccumDotWidth_acc_1343_nl;
  wire[23:0] nl_AccumDotWidth_acc_1343_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1347_nl;
  wire[24:0] nl_AccumDotWidth_acc_1347_nl;
  wire[21:0] AccumDotWidth_acc_1341_nl;
  wire[23:0] nl_AccumDotWidth_acc_1341_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1345_nl;
  wire[23:0] nl_AccumDotWidth_acc_1345_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1340_nl;
  wire[23:0] nl_AccumDotWidth_acc_1340_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1339_nl;
  wire[23:0] nl_AccumDotWidth_acc_1339_nl;
  wire[9:0] AccumDotWidth_acc_2347_nl;
  wire[10:0] nl_AccumDotWidth_acc_2347_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1322_nl;
  wire[24:0] nl_AccumDotWidth_acc_1322_nl;
  wire[21:0] AccumDotWidth_acc_1317_nl;
  wire[23:0] nl_AccumDotWidth_acc_1317_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1321_nl;
  wire[24:0] nl_AccumDotWidth_acc_1321_nl;
  wire[21:0] AccumDotWidth_acc_1315_nl;
  wire[23:0] nl_AccumDotWidth_acc_1315_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1319_nl;
  wire[23:0] nl_AccumDotWidth_acc_1319_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1314_nl;
  wire[23:0] nl_AccumDotWidth_acc_1314_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1313_nl;
  wire[23:0] nl_AccumDotWidth_acc_1313_nl;
  wire[9:0] AccumDotWidth_acc_2346_nl;
  wire[10:0] nl_AccumDotWidth_acc_2346_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1296_nl;
  wire[24:0] nl_AccumDotWidth_acc_1296_nl;
  wire[21:0] AccumDotWidth_acc_1291_nl;
  wire[23:0] nl_AccumDotWidth_acc_1291_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1295_nl;
  wire[24:0] nl_AccumDotWidth_acc_1295_nl;
  wire[21:0] AccumDotWidth_acc_1289_nl;
  wire[23:0] nl_AccumDotWidth_acc_1289_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1293_nl;
  wire[23:0] nl_AccumDotWidth_acc_1293_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1288_nl;
  wire[23:0] nl_AccumDotWidth_acc_1288_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1287_nl;
  wire[23:0] nl_AccumDotWidth_acc_1287_nl;
  wire[9:0] AccumDotWidth_acc_2345_nl;
  wire[10:0] nl_AccumDotWidth_acc_2345_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1270_nl;
  wire[24:0] nl_AccumDotWidth_acc_1270_nl;
  wire[9:0] AccumDotWidth_acc_2344_nl;
  wire[10:0] nl_AccumDotWidth_acc_2344_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1269_nl;
  wire[23:0] nl_AccumDotWidth_acc_1269_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1267_nl;
  wire[23:0] nl_AccumDotWidth_acc_1267_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1253_nl;
  wire[24:0] nl_AccumDotWidth_acc_1253_nl;
  wire[9:0] AccumDotWidth_acc_2343_nl;
  wire[10:0] nl_AccumDotWidth_acc_2343_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1252_nl;
  wire[23:0] nl_AccumDotWidth_acc_1252_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1250_nl;
  wire[23:0] nl_AccumDotWidth_acc_1250_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1236_nl;
  wire[24:0] nl_AccumDotWidth_acc_1236_nl;
  wire[9:0] AccumDotWidth_acc_2342_nl;
  wire[10:0] nl_AccumDotWidth_acc_2342_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1235_nl;
  wire[23:0] nl_AccumDotWidth_acc_1235_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1233_nl;
  wire[23:0] nl_AccumDotWidth_acc_1233_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1219_nl;
  wire[24:0] nl_AccumDotWidth_acc_1219_nl;
  wire[9:0] AccumDotWidth_acc_2341_nl;
  wire[10:0] nl_AccumDotWidth_acc_2341_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1218_nl;
  wire[23:0] nl_AccumDotWidth_acc_1218_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1216_nl;
  wire[23:0] nl_AccumDotWidth_acc_1216_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1202_nl;
  wire[24:0] nl_AccumDotWidth_acc_1202_nl;
  wire[9:0] AccumDotWidth_acc_2340_nl;
  wire[10:0] nl_AccumDotWidth_acc_2340_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1201_nl;
  wire[23:0] nl_AccumDotWidth_acc_1201_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1199_nl;
  wire[23:0] nl_AccumDotWidth_acc_1199_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1185_nl;
  wire[24:0] nl_AccumDotWidth_acc_1185_nl;
  wire[9:0] AccumDotWidth_acc_2339_nl;
  wire[10:0] nl_AccumDotWidth_acc_2339_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1184_nl;
  wire[23:0] nl_AccumDotWidth_acc_1184_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1182_nl;
  wire[23:0] nl_AccumDotWidth_acc_1182_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1168_nl;
  wire[24:0] nl_AccumDotWidth_acc_1168_nl;
  wire[9:0] AccumDotWidth_acc_2338_nl;
  wire[10:0] nl_AccumDotWidth_acc_2338_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1167_nl;
  wire[23:0] nl_AccumDotWidth_acc_1167_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1165_nl;
  wire[23:0] nl_AccumDotWidth_acc_1165_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1151_nl;
  wire[24:0] nl_AccumDotWidth_acc_1151_nl;
  wire[9:0] AccumDotWidth_acc_2337_nl;
  wire[10:0] nl_AccumDotWidth_acc_2337_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1150_nl;
  wire[23:0] nl_AccumDotWidth_acc_1150_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1148_nl;
  wire[23:0] nl_AccumDotWidth_acc_1148_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1134_nl;
  wire[24:0] nl_AccumDotWidth_acc_1134_nl;
  wire[9:0] AccumDotWidth_acc_2336_nl;
  wire[10:0] nl_AccumDotWidth_acc_2336_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1133_nl;
  wire[23:0] nl_AccumDotWidth_acc_1133_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1131_nl;
  wire[23:0] nl_AccumDotWidth_acc_1131_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1117_nl;
  wire[24:0] nl_AccumDotWidth_acc_1117_nl;
  wire[9:0] AccumDotWidth_acc_2335_nl;
  wire[10:0] nl_AccumDotWidth_acc_2335_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1116_nl;
  wire[23:0] nl_AccumDotWidth_acc_1116_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1114_nl;
  wire[23:0] nl_AccumDotWidth_acc_1114_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1100_nl;
  wire[24:0] nl_AccumDotWidth_acc_1100_nl;
  wire[9:0] AccumDotWidth_acc_2334_nl;
  wire[10:0] nl_AccumDotWidth_acc_2334_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1099_nl;
  wire[23:0] nl_AccumDotWidth_acc_1099_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1097_nl;
  wire[23:0] nl_AccumDotWidth_acc_1097_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1083_nl;
  wire[24:0] nl_AccumDotWidth_acc_1083_nl;
  wire[9:0] AccumDotWidth_acc_2333_nl;
  wire[10:0] nl_AccumDotWidth_acc_2333_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1082_nl;
  wire[23:0] nl_AccumDotWidth_acc_1082_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1080_nl;
  wire[23:0] nl_AccumDotWidth_acc_1080_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1066_nl;
  wire[24:0] nl_AccumDotWidth_acc_1066_nl;
  wire[9:0] AccumDotWidth_acc_2332_nl;
  wire[10:0] nl_AccumDotWidth_acc_2332_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1065_nl;
  wire[23:0] nl_AccumDotWidth_acc_1065_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1063_nl;
  wire[23:0] nl_AccumDotWidth_acc_1063_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1049_nl;
  wire[24:0] nl_AccumDotWidth_acc_1049_nl;
  wire[9:0] AccumDotWidth_acc_2331_nl;
  wire[10:0] nl_AccumDotWidth_acc_2331_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1048_nl;
  wire[23:0] nl_AccumDotWidth_acc_1048_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1046_nl;
  wire[23:0] nl_AccumDotWidth_acc_1046_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1032_nl;
  wire[24:0] nl_AccumDotWidth_acc_1032_nl;
  wire[9:0] AccumDotWidth_acc_2330_nl;
  wire[10:0] nl_AccumDotWidth_acc_2330_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1031_nl;
  wire[23:0] nl_AccumDotWidth_acc_1031_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1029_nl;
  wire[23:0] nl_AccumDotWidth_acc_1029_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1015_nl;
  wire[24:0] nl_AccumDotWidth_acc_1015_nl;
  wire[9:0] AccumDotWidth_acc_2329_nl;
  wire[10:0] nl_AccumDotWidth_acc_2329_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1014_nl;
  wire[23:0] nl_AccumDotWidth_acc_1014_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_1012_nl;
  wire[23:0] nl_AccumDotWidth_acc_1012_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_998_nl;
  wire[24:0] nl_AccumDotWidth_acc_998_nl;
  wire[21:0] AccumDotWidth_acc_993_nl;
  wire[23:0] nl_AccumDotWidth_acc_993_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_997_nl;
  wire[24:0] nl_AccumDotWidth_acc_997_nl;
  wire[21:0] AccumDotWidth_acc_991_nl;
  wire[23:0] nl_AccumDotWidth_acc_991_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_995_nl;
  wire[23:0] nl_AccumDotWidth_acc_995_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_990_nl;
  wire[23:0] nl_AccumDotWidth_acc_990_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_989_nl;
  wire[23:0] nl_AccumDotWidth_acc_989_nl;
  wire[9:0] AccumDotWidth_acc_2328_nl;
  wire[10:0] nl_AccumDotWidth_acc_2328_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_972_nl;
  wire[24:0] nl_AccumDotWidth_acc_972_nl;
  wire[21:0] AccumDotWidth_acc_967_nl;
  wire[23:0] nl_AccumDotWidth_acc_967_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_971_nl;
  wire[24:0] nl_AccumDotWidth_acc_971_nl;
  wire[21:0] AccumDotWidth_acc_965_nl;
  wire[23:0] nl_AccumDotWidth_acc_965_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_969_nl;
  wire[23:0] nl_AccumDotWidth_acc_969_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_964_nl;
  wire[23:0] nl_AccumDotWidth_acc_964_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_963_nl;
  wire[23:0] nl_AccumDotWidth_acc_963_nl;
  wire[9:0] AccumDotWidth_acc_2327_nl;
  wire[10:0] nl_AccumDotWidth_acc_2327_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_946_nl;
  wire[24:0] nl_AccumDotWidth_acc_946_nl;
  wire[21:0] AccumDotWidth_acc_941_nl;
  wire[23:0] nl_AccumDotWidth_acc_941_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_945_nl;
  wire[24:0] nl_AccumDotWidth_acc_945_nl;
  wire[21:0] AccumDotWidth_acc_939_nl;
  wire[23:0] nl_AccumDotWidth_acc_939_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_943_nl;
  wire[23:0] nl_AccumDotWidth_acc_943_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_938_nl;
  wire[23:0] nl_AccumDotWidth_acc_938_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_937_nl;
  wire[23:0] nl_AccumDotWidth_acc_937_nl;
  wire[9:0] AccumDotWidth_acc_2326_nl;
  wire[10:0] nl_AccumDotWidth_acc_2326_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_920_nl;
  wire[24:0] nl_AccumDotWidth_acc_920_nl;
  wire[21:0] AccumDotWidth_acc_915_nl;
  wire[23:0] nl_AccumDotWidth_acc_915_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_919_nl;
  wire[24:0] nl_AccumDotWidth_acc_919_nl;
  wire[21:0] AccumDotWidth_acc_913_nl;
  wire[23:0] nl_AccumDotWidth_acc_913_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_917_nl;
  wire[23:0] nl_AccumDotWidth_acc_917_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_912_nl;
  wire[23:0] nl_AccumDotWidth_acc_912_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_911_nl;
  wire[23:0] nl_AccumDotWidth_acc_911_nl;
  wire[9:0] AccumDotWidth_acc_2325_nl;
  wire[10:0] nl_AccumDotWidth_acc_2325_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_894_nl;
  wire[24:0] nl_AccumDotWidth_acc_894_nl;
  wire[21:0] AccumDotWidth_acc_889_nl;
  wire[23:0] nl_AccumDotWidth_acc_889_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_893_nl;
  wire[24:0] nl_AccumDotWidth_acc_893_nl;
  wire[21:0] AccumDotWidth_acc_887_nl;
  wire[23:0] nl_AccumDotWidth_acc_887_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_891_nl;
  wire[23:0] nl_AccumDotWidth_acc_891_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_886_nl;
  wire[23:0] nl_AccumDotWidth_acc_886_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_885_nl;
  wire[23:0] nl_AccumDotWidth_acc_885_nl;
  wire[9:0] AccumDotWidth_acc_2324_nl;
  wire[10:0] nl_AccumDotWidth_acc_2324_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_868_nl;
  wire[24:0] nl_AccumDotWidth_acc_868_nl;
  wire[21:0] AccumDotWidth_acc_863_nl;
  wire[23:0] nl_AccumDotWidth_acc_863_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_867_nl;
  wire[24:0] nl_AccumDotWidth_acc_867_nl;
  wire[21:0] AccumDotWidth_acc_861_nl;
  wire[23:0] nl_AccumDotWidth_acc_861_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_865_nl;
  wire[23:0] nl_AccumDotWidth_acc_865_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_860_nl;
  wire[23:0] nl_AccumDotWidth_acc_860_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_859_nl;
  wire[23:0] nl_AccumDotWidth_acc_859_nl;
  wire[9:0] AccumDotWidth_acc_2323_nl;
  wire[10:0] nl_AccumDotWidth_acc_2323_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_842_nl;
  wire[24:0] nl_AccumDotWidth_acc_842_nl;
  wire[21:0] AccumDotWidth_acc_837_nl;
  wire[23:0] nl_AccumDotWidth_acc_837_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_841_nl;
  wire[24:0] nl_AccumDotWidth_acc_841_nl;
  wire[21:0] AccumDotWidth_acc_835_nl;
  wire[23:0] nl_AccumDotWidth_acc_835_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_839_nl;
  wire[23:0] nl_AccumDotWidth_acc_839_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_834_nl;
  wire[23:0] nl_AccumDotWidth_acc_834_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_833_nl;
  wire[23:0] nl_AccumDotWidth_acc_833_nl;
  wire[9:0] AccumDotWidth_acc_2322_nl;
  wire[10:0] nl_AccumDotWidth_acc_2322_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_816_nl;
  wire[24:0] nl_AccumDotWidth_acc_816_nl;
  wire[21:0] AccumDotWidth_acc_811_nl;
  wire[23:0] nl_AccumDotWidth_acc_811_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_815_nl;
  wire[24:0] nl_AccumDotWidth_acc_815_nl;
  wire[21:0] AccumDotWidth_acc_809_nl;
  wire[23:0] nl_AccumDotWidth_acc_809_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_813_nl;
  wire[23:0] nl_AccumDotWidth_acc_813_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_808_nl;
  wire[23:0] nl_AccumDotWidth_acc_808_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_807_nl;
  wire[23:0] nl_AccumDotWidth_acc_807_nl;
  wire[9:0] AccumDotWidth_acc_2321_nl;
  wire[10:0] nl_AccumDotWidth_acc_2321_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_790_nl;
  wire[24:0] nl_AccumDotWidth_acc_790_nl;
  wire[21:0] AccumDotWidth_acc_785_nl;
  wire[23:0] nl_AccumDotWidth_acc_785_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_789_nl;
  wire[24:0] nl_AccumDotWidth_acc_789_nl;
  wire[21:0] AccumDotWidth_acc_783_nl;
  wire[23:0] nl_AccumDotWidth_acc_783_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_787_nl;
  wire[23:0] nl_AccumDotWidth_acc_787_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_782_nl;
  wire[23:0] nl_AccumDotWidth_acc_782_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_781_nl;
  wire[23:0] nl_AccumDotWidth_acc_781_nl;
  wire[9:0] AccumDotWidth_acc_2320_nl;
  wire[10:0] nl_AccumDotWidth_acc_2320_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_764_nl;
  wire[24:0] nl_AccumDotWidth_acc_764_nl;
  wire[21:0] AccumDotWidth_acc_759_nl;
  wire[23:0] nl_AccumDotWidth_acc_759_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_763_nl;
  wire[24:0] nl_AccumDotWidth_acc_763_nl;
  wire[21:0] AccumDotWidth_acc_757_nl;
  wire[23:0] nl_AccumDotWidth_acc_757_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_761_nl;
  wire[23:0] nl_AccumDotWidth_acc_761_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_756_nl;
  wire[23:0] nl_AccumDotWidth_acc_756_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_755_nl;
  wire[23:0] nl_AccumDotWidth_acc_755_nl;
  wire[9:0] AccumDotWidth_acc_2319_nl;
  wire[10:0] nl_AccumDotWidth_acc_2319_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_738_nl;
  wire[24:0] nl_AccumDotWidth_acc_738_nl;
  wire[21:0] AccumDotWidth_acc_733_nl;
  wire[23:0] nl_AccumDotWidth_acc_733_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_737_nl;
  wire[24:0] nl_AccumDotWidth_acc_737_nl;
  wire[21:0] AccumDotWidth_acc_731_nl;
  wire[23:0] nl_AccumDotWidth_acc_731_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_735_nl;
  wire[23:0] nl_AccumDotWidth_acc_735_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_730_nl;
  wire[23:0] nl_AccumDotWidth_acc_730_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_729_nl;
  wire[23:0] nl_AccumDotWidth_acc_729_nl;
  wire[9:0] AccumDotWidth_acc_2318_nl;
  wire[10:0] nl_AccumDotWidth_acc_2318_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_712_nl;
  wire[24:0] nl_AccumDotWidth_acc_712_nl;
  wire[21:0] AccumDotWidth_acc_707_nl;
  wire[23:0] nl_AccumDotWidth_acc_707_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_711_nl;
  wire[24:0] nl_AccumDotWidth_acc_711_nl;
  wire[21:0] AccumDotWidth_acc_705_nl;
  wire[23:0] nl_AccumDotWidth_acc_705_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_709_nl;
  wire[23:0] nl_AccumDotWidth_acc_709_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_704_nl;
  wire[23:0] nl_AccumDotWidth_acc_704_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_703_nl;
  wire[23:0] nl_AccumDotWidth_acc_703_nl;
  wire[9:0] AccumDotWidth_acc_2317_nl;
  wire[10:0] nl_AccumDotWidth_acc_2317_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_686_nl;
  wire[24:0] nl_AccumDotWidth_acc_686_nl;
  wire[21:0] AccumDotWidth_acc_681_nl;
  wire[23:0] nl_AccumDotWidth_acc_681_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_685_nl;
  wire[24:0] nl_AccumDotWidth_acc_685_nl;
  wire[21:0] AccumDotWidth_acc_679_nl;
  wire[23:0] nl_AccumDotWidth_acc_679_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_683_nl;
  wire[23:0] nl_AccumDotWidth_acc_683_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_678_nl;
  wire[23:0] nl_AccumDotWidth_acc_678_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_677_nl;
  wire[23:0] nl_AccumDotWidth_acc_677_nl;
  wire[9:0] AccumDotWidth_acc_2316_nl;
  wire[10:0] nl_AccumDotWidth_acc_2316_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_660_nl;
  wire[24:0] nl_AccumDotWidth_acc_660_nl;
  wire[21:0] AccumDotWidth_acc_655_nl;
  wire[23:0] nl_AccumDotWidth_acc_655_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_659_nl;
  wire[24:0] nl_AccumDotWidth_acc_659_nl;
  wire[21:0] AccumDotWidth_acc_653_nl;
  wire[23:0] nl_AccumDotWidth_acc_653_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_657_nl;
  wire[23:0] nl_AccumDotWidth_acc_657_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_652_nl;
  wire[23:0] nl_AccumDotWidth_acc_652_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_651_nl;
  wire[23:0] nl_AccumDotWidth_acc_651_nl;
  wire[9:0] AccumDotWidth_acc_2315_nl;
  wire[10:0] nl_AccumDotWidth_acc_2315_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_634_nl;
  wire[24:0] nl_AccumDotWidth_acc_634_nl;
  wire[21:0] AccumDotWidth_acc_629_nl;
  wire[23:0] nl_AccumDotWidth_acc_629_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_633_nl;
  wire[24:0] nl_AccumDotWidth_acc_633_nl;
  wire[21:0] AccumDotWidth_acc_627_nl;
  wire[23:0] nl_AccumDotWidth_acc_627_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_631_nl;
  wire[23:0] nl_AccumDotWidth_acc_631_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_626_nl;
  wire[23:0] nl_AccumDotWidth_acc_626_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_625_nl;
  wire[23:0] nl_AccumDotWidth_acc_625_nl;
  wire[9:0] AccumDotWidth_acc_2314_nl;
  wire[10:0] nl_AccumDotWidth_acc_2314_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_608_nl;
  wire[24:0] nl_AccumDotWidth_acc_608_nl;
  wire[21:0] AccumDotWidth_acc_603_nl;
  wire[23:0] nl_AccumDotWidth_acc_603_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_607_nl;
  wire[24:0] nl_AccumDotWidth_acc_607_nl;
  wire[21:0] AccumDotWidth_acc_601_nl;
  wire[23:0] nl_AccumDotWidth_acc_601_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_605_nl;
  wire[23:0] nl_AccumDotWidth_acc_605_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_600_nl;
  wire[23:0] nl_AccumDotWidth_acc_600_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_599_nl;
  wire[23:0] nl_AccumDotWidth_acc_599_nl;
  wire[9:0] AccumDotWidth_acc_2313_nl;
  wire[10:0] nl_AccumDotWidth_acc_2313_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_582_nl;
  wire[24:0] nl_AccumDotWidth_acc_582_nl;
  wire[9:0] AccumDotWidth_acc_2312_nl;
  wire[10:0] nl_AccumDotWidth_acc_2312_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_581_nl;
  wire[23:0] nl_AccumDotWidth_acc_581_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_579_nl;
  wire[23:0] nl_AccumDotWidth_acc_579_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_565_nl;
  wire[24:0] nl_AccumDotWidth_acc_565_nl;
  wire[9:0] AccumDotWidth_acc_2311_nl;
  wire[10:0] nl_AccumDotWidth_acc_2311_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_564_nl;
  wire[23:0] nl_AccumDotWidth_acc_564_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_562_nl;
  wire[23:0] nl_AccumDotWidth_acc_562_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_548_nl;
  wire[24:0] nl_AccumDotWidth_acc_548_nl;
  wire[9:0] AccumDotWidth_acc_2310_nl;
  wire[10:0] nl_AccumDotWidth_acc_2310_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_547_nl;
  wire[23:0] nl_AccumDotWidth_acc_547_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_545_nl;
  wire[23:0] nl_AccumDotWidth_acc_545_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_531_nl;
  wire[24:0] nl_AccumDotWidth_acc_531_nl;
  wire[9:0] AccumDotWidth_acc_2309_nl;
  wire[10:0] nl_AccumDotWidth_acc_2309_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_530_nl;
  wire[23:0] nl_AccumDotWidth_acc_530_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_528_nl;
  wire[23:0] nl_AccumDotWidth_acc_528_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_514_nl;
  wire[24:0] nl_AccumDotWidth_acc_514_nl;
  wire[9:0] AccumDotWidth_acc_2308_nl;
  wire[10:0] nl_AccumDotWidth_acc_2308_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_513_nl;
  wire[23:0] nl_AccumDotWidth_acc_513_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_511_nl;
  wire[23:0] nl_AccumDotWidth_acc_511_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_497_nl;
  wire[24:0] nl_AccumDotWidth_acc_497_nl;
  wire[9:0] AccumDotWidth_acc_2307_nl;
  wire[10:0] nl_AccumDotWidth_acc_2307_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_496_nl;
  wire[23:0] nl_AccumDotWidth_acc_496_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_494_nl;
  wire[23:0] nl_AccumDotWidth_acc_494_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_480_nl;
  wire[24:0] nl_AccumDotWidth_acc_480_nl;
  wire[9:0] AccumDotWidth_acc_2306_nl;
  wire[10:0] nl_AccumDotWidth_acc_2306_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_479_nl;
  wire[23:0] nl_AccumDotWidth_acc_479_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_477_nl;
  wire[23:0] nl_AccumDotWidth_acc_477_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_463_nl;
  wire[24:0] nl_AccumDotWidth_acc_463_nl;
  wire[9:0] AccumDotWidth_acc_2305_nl;
  wire[10:0] nl_AccumDotWidth_acc_2305_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_462_nl;
  wire[23:0] nl_AccumDotWidth_acc_462_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_460_nl;
  wire[23:0] nl_AccumDotWidth_acc_460_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_447_nl;
  wire[23:0] nl_AccumDotWidth_acc_447_nl;
  wire[9:0] AccumDotWidth_acc_2304_nl;
  wire[10:0] nl_AccumDotWidth_acc_2304_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_446_nl;
  wire[23:0] nl_AccumDotWidth_acc_446_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_445_nl;
  wire[23:0] nl_AccumDotWidth_acc_445_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_436_nl;
  wire[23:0] nl_AccumDotWidth_acc_436_nl;
  wire[9:0] AccumDotWidth_acc_2303_nl;
  wire[10:0] nl_AccumDotWidth_acc_2303_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_435_nl;
  wire[23:0] nl_AccumDotWidth_acc_435_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_434_nl;
  wire[23:0] nl_AccumDotWidth_acc_434_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_425_nl;
  wire[23:0] nl_AccumDotWidth_acc_425_nl;
  wire[9:0] AccumDotWidth_acc_2302_nl;
  wire[10:0] nl_AccumDotWidth_acc_2302_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_424_nl;
  wire[23:0] nl_AccumDotWidth_acc_424_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_423_nl;
  wire[23:0] nl_AccumDotWidth_acc_423_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_414_nl;
  wire[23:0] nl_AccumDotWidth_acc_414_nl;
  wire[9:0] AccumDotWidth_acc_2301_nl;
  wire[10:0] nl_AccumDotWidth_acc_2301_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_413_nl;
  wire[23:0] nl_AccumDotWidth_acc_413_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_412_nl;
  wire[23:0] nl_AccumDotWidth_acc_412_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_403_nl;
  wire[23:0] nl_AccumDotWidth_acc_403_nl;
  wire[9:0] AccumDotWidth_acc_2300_nl;
  wire[10:0] nl_AccumDotWidth_acc_2300_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_402_nl;
  wire[23:0] nl_AccumDotWidth_acc_402_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_401_nl;
  wire[23:0] nl_AccumDotWidth_acc_401_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_392_nl;
  wire[23:0] nl_AccumDotWidth_acc_392_nl;
  wire[9:0] AccumDotWidth_acc_2299_nl;
  wire[10:0] nl_AccumDotWidth_acc_2299_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_391_nl;
  wire[23:0] nl_AccumDotWidth_acc_391_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_390_nl;
  wire[23:0] nl_AccumDotWidth_acc_390_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_381_nl;
  wire[23:0] nl_AccumDotWidth_acc_381_nl;
  wire[9:0] AccumDotWidth_acc_2298_nl;
  wire[10:0] nl_AccumDotWidth_acc_2298_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_380_nl;
  wire[23:0] nl_AccumDotWidth_acc_380_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_379_nl;
  wire[23:0] nl_AccumDotWidth_acc_379_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_370_nl;
  wire[23:0] nl_AccumDotWidth_acc_370_nl;
  wire[9:0] AccumDotWidth_acc_2297_nl;
  wire[10:0] nl_AccumDotWidth_acc_2297_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_369_nl;
  wire[23:0] nl_AccumDotWidth_acc_369_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_368_nl;
  wire[23:0] nl_AccumDotWidth_acc_368_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_358_nl;
  wire[24:0] nl_AccumDotWidth_acc_358_nl;
  wire[9:0] AccumDotWidth_acc_2296_nl;
  wire[10:0] nl_AccumDotWidth_acc_2296_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_357_nl;
  wire[23:0] nl_AccumDotWidth_acc_357_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_355_nl;
  wire[23:0] nl_AccumDotWidth_acc_355_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_341_nl;
  wire[24:0] nl_AccumDotWidth_acc_341_nl;
  wire[9:0] AccumDotWidth_acc_2295_nl;
  wire[10:0] nl_AccumDotWidth_acc_2295_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_340_nl;
  wire[23:0] nl_AccumDotWidth_acc_340_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_338_nl;
  wire[23:0] nl_AccumDotWidth_acc_338_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_324_nl;
  wire[24:0] nl_AccumDotWidth_acc_324_nl;
  wire[9:0] AccumDotWidth_acc_2294_nl;
  wire[10:0] nl_AccumDotWidth_acc_2294_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_323_nl;
  wire[23:0] nl_AccumDotWidth_acc_323_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_321_nl;
  wire[23:0] nl_AccumDotWidth_acc_321_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_307_nl;
  wire[24:0] nl_AccumDotWidth_acc_307_nl;
  wire[9:0] AccumDotWidth_acc_2293_nl;
  wire[10:0] nl_AccumDotWidth_acc_2293_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_306_nl;
  wire[23:0] nl_AccumDotWidth_acc_306_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_304_nl;
  wire[23:0] nl_AccumDotWidth_acc_304_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_290_nl;
  wire[24:0] nl_AccumDotWidth_acc_290_nl;
  wire[9:0] AccumDotWidth_acc_2292_nl;
  wire[10:0] nl_AccumDotWidth_acc_2292_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_289_nl;
  wire[23:0] nl_AccumDotWidth_acc_289_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_287_nl;
  wire[23:0] nl_AccumDotWidth_acc_287_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_273_nl;
  wire[24:0] nl_AccumDotWidth_acc_273_nl;
  wire[9:0] AccumDotWidth_acc_2291_nl;
  wire[10:0] nl_AccumDotWidth_acc_2291_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_272_nl;
  wire[23:0] nl_AccumDotWidth_acc_272_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_270_nl;
  wire[23:0] nl_AccumDotWidth_acc_270_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_256_nl;
  wire[24:0] nl_AccumDotWidth_acc_256_nl;
  wire[9:0] AccumDotWidth_acc_2290_nl;
  wire[10:0] nl_AccumDotWidth_acc_2290_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_255_nl;
  wire[23:0] nl_AccumDotWidth_acc_255_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_253_nl;
  wire[23:0] nl_AccumDotWidth_acc_253_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_239_nl;
  wire[24:0] nl_AccumDotWidth_acc_239_nl;
  wire[9:0] AccumDotWidth_acc_2289_nl;
  wire[10:0] nl_AccumDotWidth_acc_2289_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_238_nl;
  wire[23:0] nl_AccumDotWidth_acc_238_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_236_nl;
  wire[23:0] nl_AccumDotWidth_acc_236_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_222_nl;
  wire[24:0] nl_AccumDotWidth_acc_222_nl;
  wire[9:0] AccumDotWidth_acc_2288_nl;
  wire[10:0] nl_AccumDotWidth_acc_2288_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_221_nl;
  wire[23:0] nl_AccumDotWidth_acc_221_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_219_nl;
  wire[23:0] nl_AccumDotWidth_acc_219_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_205_nl;
  wire[24:0] nl_AccumDotWidth_acc_205_nl;
  wire[9:0] AccumDotWidth_acc_2287_nl;
  wire[10:0] nl_AccumDotWidth_acc_2287_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_204_nl;
  wire[23:0] nl_AccumDotWidth_acc_204_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_202_nl;
  wire[23:0] nl_AccumDotWidth_acc_202_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_188_nl;
  wire[24:0] nl_AccumDotWidth_acc_188_nl;
  wire[9:0] AccumDotWidth_acc_2286_nl;
  wire[10:0] nl_AccumDotWidth_acc_2286_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_187_nl;
  wire[23:0] nl_AccumDotWidth_acc_187_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_185_nl;
  wire[23:0] nl_AccumDotWidth_acc_185_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_171_nl;
  wire[24:0] nl_AccumDotWidth_acc_171_nl;
  wire[9:0] AccumDotWidth_acc_2285_nl;
  wire[10:0] nl_AccumDotWidth_acc_2285_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_170_nl;
  wire[23:0] nl_AccumDotWidth_acc_170_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_168_nl;
  wire[23:0] nl_AccumDotWidth_acc_168_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_154_nl;
  wire[24:0] nl_AccumDotWidth_acc_154_nl;
  wire[9:0] AccumDotWidth_acc_2284_nl;
  wire[10:0] nl_AccumDotWidth_acc_2284_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_153_nl;
  wire[23:0] nl_AccumDotWidth_acc_153_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_151_nl;
  wire[23:0] nl_AccumDotWidth_acc_151_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_137_nl;
  wire[24:0] nl_AccumDotWidth_acc_137_nl;
  wire[9:0] AccumDotWidth_acc_2283_nl;
  wire[10:0] nl_AccumDotWidth_acc_2283_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_136_nl;
  wire[23:0] nl_AccumDotWidth_acc_136_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_134_nl;
  wire[23:0] nl_AccumDotWidth_acc_134_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_120_nl;
  wire[24:0] nl_AccumDotWidth_acc_120_nl;
  wire[9:0] AccumDotWidth_acc_2282_nl;
  wire[10:0] nl_AccumDotWidth_acc_2282_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_119_nl;
  wire[23:0] nl_AccumDotWidth_acc_119_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_117_nl;
  wire[23:0] nl_AccumDotWidth_acc_117_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_103_nl;
  wire[24:0] nl_AccumDotWidth_acc_103_nl;
  wire[9:0] AccumDotWidth_acc_2281_nl;
  wire[10:0] nl_AccumDotWidth_acc_2281_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_102_nl;
  wire[23:0] nl_AccumDotWidth_acc_102_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_100_nl;
  wire[23:0] nl_AccumDotWidth_acc_100_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_87_nl;
  wire[23:0] nl_AccumDotWidth_acc_87_nl;
  wire[9:0] AccumDotWidth_acc_2280_nl;
  wire[10:0] nl_AccumDotWidth_acc_2280_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_86_nl;
  wire[23:0] nl_AccumDotWidth_acc_86_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_85_nl;
  wire[23:0] nl_AccumDotWidth_acc_85_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_76_nl;
  wire[23:0] nl_AccumDotWidth_acc_76_nl;
  wire[9:0] AccumDotWidth_acc_2279_nl;
  wire[10:0] nl_AccumDotWidth_acc_2279_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_75_nl;
  wire[23:0] nl_AccumDotWidth_acc_75_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_74_nl;
  wire[23:0] nl_AccumDotWidth_acc_74_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_65_nl;
  wire[23:0] nl_AccumDotWidth_acc_65_nl;
  wire[9:0] AccumDotWidth_acc_2278_nl;
  wire[10:0] nl_AccumDotWidth_acc_2278_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_64_nl;
  wire[23:0] nl_AccumDotWidth_acc_64_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_63_nl;
  wire[23:0] nl_AccumDotWidth_acc_63_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_54_nl;
  wire[23:0] nl_AccumDotWidth_acc_54_nl;
  wire[9:0] AccumDotWidth_acc_2277_nl;
  wire[10:0] nl_AccumDotWidth_acc_2277_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_53_nl;
  wire[23:0] nl_AccumDotWidth_acc_53_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_52_nl;
  wire[23:0] nl_AccumDotWidth_acc_52_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_43_nl;
  wire[23:0] nl_AccumDotWidth_acc_43_nl;
  wire[9:0] AccumDotWidth_acc_2276_nl;
  wire[10:0] nl_AccumDotWidth_acc_2276_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_42_nl;
  wire[23:0] nl_AccumDotWidth_acc_42_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_41_nl;
  wire[23:0] nl_AccumDotWidth_acc_41_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_32_nl;
  wire[23:0] nl_AccumDotWidth_acc_32_nl;
  wire[9:0] AccumDotWidth_acc_2275_nl;
  wire[10:0] nl_AccumDotWidth_acc_2275_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_31_nl;
  wire[23:0] nl_AccumDotWidth_acc_31_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_30_nl;
  wire[23:0] nl_AccumDotWidth_acc_30_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_21_nl;
  wire[23:0] nl_AccumDotWidth_acc_21_nl;
  wire[9:0] AccumDotWidth_acc_2274_nl;
  wire[10:0] nl_AccumDotWidth_acc_2274_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_20_nl;
  wire[23:0] nl_AccumDotWidth_acc_20_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_19_nl;
  wire[23:0] nl_AccumDotWidth_acc_19_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_nl;
  wire[23:0] nl_AccumDotWidth_acc_nl;
  wire[9:0] AccumDotWidth_acc_2273_nl;
  wire[10:0] nl_AccumDotWidth_acc_2273_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_9_nl;
  wire[23:0] nl_AccumDotWidth_acc_9_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[21:0] AccumDotWidth_acc_8_nl;
  wire[23:0] nl_AccumDotWidth_acc_8_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[29:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [219:0] nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat;
  assign nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat = {1'b0 ,
      layer5_out_rsci_idat_218_198 , 1'b0 , layer5_out_rsci_idat_196_176 , 1'b0 ,
      layer5_out_rsci_idat_174_154 , 1'b0 , layer5_out_rsci_idat_152_132 , 1'b0 ,
      layer5_out_rsci_idat_130_110 , 1'b0 , layer5_out_rsci_idat_108_88 , 1'b0 ,
      layer5_out_rsci_idat_86_66 , 1'b0 , layer5_out_rsci_idat_64_44 , 1'b0 , layer5_out_rsci_idat_42_22
      , 1'b0 , layer5_out_rsci_idat_20_0};
  econ_4x4_d10_core_input_1_rsci econ_4x4_d10_core_input_1_rsci_inst (
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_layer5_out_rsci econ_4x4_d10_core_layer5_out_rsci_inst (
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .core_wten(core_wten),
      .layer5_out_rsci_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse),
      .layer5_out_rsci_idat(nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat[219:0])
    );
  econ_4x4_d10_core_const_size_in_1_rsci econ_4x4_d10_core_const_size_in_1_rsci_inst
      (
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_out_1_rsci econ_4x4_d10_core_const_size_out_1_rsci_inst
      (
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w2_rsci econ_4x4_d10_core_w2_rsci_inst (
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b2_rsci econ_4x4_d10_core_b2_rsci_inst (
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_w4_rsci econ_4x4_d10_core_w4_rsci_inst (
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b4_rsci econ_4x4_d10_core_b4_rsci_inst (
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj econ_4x4_d10_core_input_1_rsc_triosy_obj_inst
      (
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj econ_4x4_d10_core_layer5_out_rsc_triosy_obj_inst
      (
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_inst
      (
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_inst
      (
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj econ_4x4_d10_core_w2_rsc_triosy_obj_inst (
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj econ_4x4_d10_core_b2_rsc_triosy_obj_inst (
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj econ_4x4_d10_core_w4_rsc_triosy_obj_inst (
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj econ_4x4_d10_core_b4_rsc_triosy_obj_inst (
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz),
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_staller econ_4x4_d10_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .b4_rsci_wen_comp(b4_rsci_wen_comp)
    );
  econ_4x4_d10_core_core_fsm econ_4x4_d10_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign layer5_out_and_cse = core_wen & main_stage_0_2;
  assign nl_MultLoop_acc_1146_nl = MultLoop_acc_1138_itm_1 + MultLoop_acc_1137_itm_1;
  assign MultLoop_acc_1146_nl = nl_MultLoop_acc_1146_nl[21:0];
  assign nl_MultLoop_acc_1145_nl = MultLoop_acc_1136_itm_1 + MultLoop_acc_1135_itm_1;
  assign MultLoop_acc_1145_nl = nl_MultLoop_acc_1145_nl[21:0];
  assign nl_MultLoop_acc_1150_nl = (MultLoop_acc_1146_nl) + (MultLoop_acc_1145_nl);
  assign MultLoop_acc_1150_nl = nl_MultLoop_acc_1150_nl[21:0];
  assign nl_MultLoop_acc_1149_nl = MultLoop_acc_1134_itm_1 + MultLoop_acc_1133_itm_1
      + MultLoop_acc_1132_itm_1 + MultLoop_acc_1131_itm_1;
  assign MultLoop_acc_1149_nl = nl_MultLoop_acc_1149_nl[21:0];
  assign nl_MultLoop_acc_1152_nl = (MultLoop_acc_1150_nl) + (MultLoop_acc_1149_nl);
  assign MultLoop_acc_1152_nl = nl_MultLoop_acc_1152_nl[21:0];
  assign nl_MultLoop_acc_1151_nl = MultLoop_acc_1126_itm_1 + MultLoop_acc_1125_itm_1
      + MultLoop_acc_1130_itm_1 + MultLoop_acc_1129_itm_1 + MultLoop_acc_1128_itm_1
      + MultLoop_acc_1127_itm_1 + MultLoop_acc_1124_itm_1 + MultLoop_acc_1123_itm_1;
  assign MultLoop_acc_1151_nl = nl_MultLoop_acc_1151_nl[21:0];
  assign nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1 = (MultLoop_acc_1152_nl) + (MultLoop_acc_1151_nl);
  assign MultLoop_1280_MultLoop_acc_3_ncse_sva_1 = nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1[21:0];
  assign nl_MultLoop_acc_1273_nl = MultLoop_acc_1265_itm_1 + MultLoop_acc_1264_itm_1;
  assign MultLoop_acc_1273_nl = nl_MultLoop_acc_1273_nl[21:0];
  assign nl_MultLoop_acc_1272_nl = MultLoop_acc_1263_itm_1 + MultLoop_acc_1262_itm_1;
  assign MultLoop_acc_1272_nl = nl_MultLoop_acc_1272_nl[21:0];
  assign nl_MultLoop_acc_1277_nl = (MultLoop_acc_1273_nl) + (MultLoop_acc_1272_nl);
  assign MultLoop_acc_1277_nl = nl_MultLoop_acc_1277_nl[21:0];
  assign nl_MultLoop_acc_1276_nl = MultLoop_acc_1261_itm_1 + MultLoop_acc_1260_itm_1
      + MultLoop_acc_1259_itm_1 + MultLoop_acc_1258_itm_1;
  assign MultLoop_acc_1276_nl = nl_MultLoop_acc_1276_nl[21:0];
  assign nl_MultLoop_acc_1279_nl = (MultLoop_acc_1277_nl) + (MultLoop_acc_1276_nl);
  assign MultLoop_acc_1279_nl = nl_MultLoop_acc_1279_nl[21:0];
  assign nl_MultLoop_acc_1278_nl = MultLoop_acc_1253_itm_1 + MultLoop_acc_1252_itm_1
      + MultLoop_acc_1257_itm_1 + MultLoop_acc_1256_itm_1 + MultLoop_acc_1255_itm_1
      + MultLoop_acc_1254_itm_1 + MultLoop_acc_1251_itm_1 + MultLoop_acc_1250_itm_1;
  assign MultLoop_acc_1278_nl = nl_MultLoop_acc_1278_nl[21:0];
  assign nl_layer4_out_0_sva_1 = (MultLoop_acc_1279_nl) + (MultLoop_acc_1278_nl);
  assign layer4_out_0_sva_1 = nl_layer4_out_0_sva_1[21:0];
  assign nl_MultLoop_acc_1019_nl = MultLoop_acc_1011_itm_1 + MultLoop_acc_1010_itm_1;
  assign MultLoop_acc_1019_nl = nl_MultLoop_acc_1019_nl[21:0];
  assign nl_MultLoop_acc_1018_nl = MultLoop_acc_1009_itm_1 + MultLoop_acc_1008_itm_1;
  assign MultLoop_acc_1018_nl = nl_MultLoop_acc_1018_nl[21:0];
  assign nl_MultLoop_acc_1023_nl = (MultLoop_acc_1019_nl) + (MultLoop_acc_1018_nl);
  assign MultLoop_acc_1023_nl = nl_MultLoop_acc_1023_nl[21:0];
  assign nl_MultLoop_acc_1022_nl = MultLoop_acc_1007_itm_1 + MultLoop_acc_1006_itm_1
      + MultLoop_acc_1005_itm_1 + MultLoop_acc_1004_itm_1;
  assign MultLoop_acc_1022_nl = nl_MultLoop_acc_1022_nl[21:0];
  assign nl_MultLoop_acc_1025_nl = (MultLoop_acc_1023_nl) + (MultLoop_acc_1022_nl);
  assign MultLoop_acc_1025_nl = nl_MultLoop_acc_1025_nl[21:0];
  assign nl_MultLoop_acc_1024_nl = MultLoop_acc_999_itm_1 + MultLoop_acc_998_itm_1
      + MultLoop_acc_1003_itm_1 + MultLoop_acc_1002_itm_1 + MultLoop_acc_1001_itm_1
      + MultLoop_acc_1000_itm_1 + MultLoop_acc_997_itm_1 + MultLoop_acc_996_itm_1;
  assign MultLoop_acc_1024_nl = nl_MultLoop_acc_1024_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1 = (MultLoop_acc_1025_nl)
      + (MultLoop_acc_1024_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1[21:0];
  assign nl_MultLoop_acc_134_nl = MultLoop_acc_130_itm_1 + MultLoop_acc_121_itm_1;
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[21:0];
  assign nl_MultLoop_acc_129_nl = MultLoop_acc_120_itm_1 + MultLoop_acc_119_itm_1;
  assign MultLoop_acc_129_nl = nl_MultLoop_acc_129_nl[21:0];
  assign nl_MultLoop_acc_136_nl = (MultLoop_acc_134_nl) + (MultLoop_acc_129_nl);
  assign MultLoop_acc_136_nl = nl_MultLoop_acc_136_nl[21:0];
  assign nl_MultLoop_acc_133_nl = MultLoop_acc_118_itm_1 + MultLoop_acc_117_itm_1
      + MultLoop_acc_116_itm_1 + MultLoop_acc_115_itm_1;
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[21:0];
  assign nl_MultLoop_acc_nl = (MultLoop_acc_136_nl) + (MultLoop_acc_133_nl);
  assign MultLoop_acc_nl = nl_MultLoop_acc_nl[21:0];
  assign nl_MultLoop_acc_135_nl = MultLoop_acc_110_itm_1 + MultLoop_acc_109_itm_1
      + MultLoop_acc_114_itm_1 + MultLoop_acc_113_itm_1 + MultLoop_acc_112_itm_1
      + MultLoop_acc_111_itm_1 + MultLoop_acc_108_itm_1 + MultLoop_acc_107_itm_1;
  assign MultLoop_acc_135_nl = nl_MultLoop_acc_135_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1 = (MultLoop_acc_nl)
      + (MultLoop_acc_135_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1[21:0];
  assign nl_MultLoop_acc_892_nl = MultLoop_acc_884_itm_1 + MultLoop_acc_883_itm_1;
  assign MultLoop_acc_892_nl = nl_MultLoop_acc_892_nl[21:0];
  assign nl_MultLoop_acc_891_nl = MultLoop_acc_882_itm_1 + MultLoop_acc_881_itm_1;
  assign MultLoop_acc_891_nl = nl_MultLoop_acc_891_nl[21:0];
  assign nl_MultLoop_acc_896_nl = (MultLoop_acc_892_nl) + (MultLoop_acc_891_nl);
  assign MultLoop_acc_896_nl = nl_MultLoop_acc_896_nl[21:0];
  assign nl_MultLoop_acc_895_nl = MultLoop_acc_880_itm_1 + MultLoop_acc_879_itm_1
      + MultLoop_acc_878_itm_1 + MultLoop_acc_877_itm_1;
  assign MultLoop_acc_895_nl = nl_MultLoop_acc_895_nl[21:0];
  assign nl_MultLoop_acc_898_nl = (MultLoop_acc_896_nl) + (MultLoop_acc_895_nl);
  assign MultLoop_acc_898_nl = nl_MultLoop_acc_898_nl[21:0];
  assign nl_MultLoop_acc_897_nl = MultLoop_acc_872_itm_1 + MultLoop_acc_871_itm_1
      + MultLoop_acc_876_itm_1 + MultLoop_acc_875_itm_1 + MultLoop_acc_874_itm_1
      + MultLoop_acc_873_itm_1 + MultLoop_acc_870_itm_1 + MultLoop_acc_869_itm_1;
  assign MultLoop_acc_897_nl = nl_MultLoop_acc_897_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1 = (MultLoop_acc_898_nl)
      + (MultLoop_acc_897_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1[21:0];
  assign nl_MultLoop_acc_257_nl = MultLoop_acc_249_itm_1 + MultLoop_acc_248_itm_1;
  assign MultLoop_acc_257_nl = nl_MultLoop_acc_257_nl[21:0];
  assign nl_MultLoop_acc_256_nl = MultLoop_acc_247_itm_1 + MultLoop_acc_246_itm_1;
  assign MultLoop_acc_256_nl = nl_MultLoop_acc_256_nl[21:0];
  assign nl_MultLoop_acc_261_nl = (MultLoop_acc_257_nl) + (MultLoop_acc_256_nl);
  assign MultLoop_acc_261_nl = nl_MultLoop_acc_261_nl[21:0];
  assign nl_MultLoop_acc_260_nl = MultLoop_acc_245_itm_1 + MultLoop_acc_244_itm_1
      + MultLoop_acc_243_itm_1 + MultLoop_acc_242_itm_1;
  assign MultLoop_acc_260_nl = nl_MultLoop_acc_260_nl[21:0];
  assign nl_MultLoop_acc_263_nl = (MultLoop_acc_261_nl) + (MultLoop_acc_260_nl);
  assign MultLoop_acc_263_nl = nl_MultLoop_acc_263_nl[21:0];
  assign nl_MultLoop_acc_262_nl = MultLoop_acc_237_itm_1 + MultLoop_acc_236_itm_1
      + MultLoop_acc_241_itm_1 + MultLoop_acc_240_itm_1 + MultLoop_acc_239_itm_1
      + MultLoop_acc_238_itm_1 + MultLoop_acc_235_itm_1 + MultLoop_acc_234_itm_1;
  assign MultLoop_acc_262_nl = nl_MultLoop_acc_262_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1 = (MultLoop_acc_263_nl)
      + (MultLoop_acc_262_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1[21:0];
  assign nl_MultLoop_acc_765_nl = MultLoop_acc_757_itm_1 + MultLoop_acc_756_itm_1;
  assign MultLoop_acc_765_nl = nl_MultLoop_acc_765_nl[21:0];
  assign nl_MultLoop_acc_764_nl = MultLoop_acc_755_itm_1 + MultLoop_acc_754_itm_1;
  assign MultLoop_acc_764_nl = nl_MultLoop_acc_764_nl[21:0];
  assign nl_MultLoop_acc_769_nl = (MultLoop_acc_765_nl) + (MultLoop_acc_764_nl);
  assign MultLoop_acc_769_nl = nl_MultLoop_acc_769_nl[21:0];
  assign nl_MultLoop_acc_768_nl = MultLoop_acc_753_itm_1 + MultLoop_acc_752_itm_1
      + MultLoop_acc_751_itm_1 + MultLoop_acc_750_itm_1;
  assign MultLoop_acc_768_nl = nl_MultLoop_acc_768_nl[21:0];
  assign nl_MultLoop_acc_771_nl = (MultLoop_acc_769_nl) + (MultLoop_acc_768_nl);
  assign MultLoop_acc_771_nl = nl_MultLoop_acc_771_nl[21:0];
  assign nl_MultLoop_acc_770_nl = MultLoop_acc_745_itm_1 + MultLoop_acc_744_itm_1
      + MultLoop_acc_749_itm_1 + MultLoop_acc_748_itm_1 + MultLoop_acc_747_itm_1
      + MultLoop_acc_746_itm_1 + MultLoop_acc_743_itm_1 + MultLoop_acc_742_itm_1;
  assign MultLoop_acc_770_nl = nl_MultLoop_acc_770_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1 = (MultLoop_acc_771_nl)
      + (MultLoop_acc_770_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1[21:0];
  assign nl_MultLoop_acc_384_nl = MultLoop_acc_376_itm_1 + MultLoop_acc_375_itm_1;
  assign MultLoop_acc_384_nl = nl_MultLoop_acc_384_nl[21:0];
  assign nl_MultLoop_acc_383_nl = MultLoop_acc_374_itm_1 + MultLoop_acc_373_itm_1;
  assign MultLoop_acc_383_nl = nl_MultLoop_acc_383_nl[21:0];
  assign nl_MultLoop_acc_388_nl = (MultLoop_acc_384_nl) + (MultLoop_acc_383_nl);
  assign MultLoop_acc_388_nl = nl_MultLoop_acc_388_nl[21:0];
  assign nl_MultLoop_acc_387_nl = MultLoop_acc_372_itm_1 + MultLoop_acc_371_itm_1
      + MultLoop_acc_370_itm_1 + MultLoop_acc_369_itm_1;
  assign MultLoop_acc_387_nl = nl_MultLoop_acc_387_nl[21:0];
  assign nl_MultLoop_acc_390_nl = (MultLoop_acc_388_nl) + (MultLoop_acc_387_nl);
  assign MultLoop_acc_390_nl = nl_MultLoop_acc_390_nl[21:0];
  assign nl_MultLoop_acc_389_nl = MultLoop_acc_364_itm_1 + MultLoop_acc_363_itm_1
      + MultLoop_acc_368_itm_1 + MultLoop_acc_367_itm_1 + MultLoop_acc_366_itm_1
      + MultLoop_acc_365_itm_1 + MultLoop_acc_362_itm_1 + MultLoop_acc_361_itm_1;
  assign MultLoop_acc_389_nl = nl_MultLoop_acc_389_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1 = (MultLoop_acc_390_nl)
      + (MultLoop_acc_389_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1[21:0];
  assign nl_MultLoop_acc_638_nl = MultLoop_acc_630_itm_1 + MultLoop_acc_629_itm_1;
  assign MultLoop_acc_638_nl = nl_MultLoop_acc_638_nl[21:0];
  assign nl_MultLoop_acc_637_nl = MultLoop_acc_628_itm_1 + MultLoop_acc_627_itm_1;
  assign MultLoop_acc_637_nl = nl_MultLoop_acc_637_nl[21:0];
  assign nl_MultLoop_acc_642_nl = (MultLoop_acc_638_nl) + (MultLoop_acc_637_nl);
  assign MultLoop_acc_642_nl = nl_MultLoop_acc_642_nl[21:0];
  assign nl_MultLoop_acc_641_nl = MultLoop_acc_626_itm_1 + MultLoop_acc_625_itm_1
      + MultLoop_acc_624_itm_1 + MultLoop_acc_623_itm_1;
  assign MultLoop_acc_641_nl = nl_MultLoop_acc_641_nl[21:0];
  assign nl_MultLoop_acc_644_nl = (MultLoop_acc_642_nl) + (MultLoop_acc_641_nl);
  assign MultLoop_acc_644_nl = nl_MultLoop_acc_644_nl[21:0];
  assign nl_MultLoop_acc_643_nl = MultLoop_acc_618_itm_1 + MultLoop_acc_617_itm_1
      + MultLoop_acc_622_itm_1 + MultLoop_acc_621_itm_1 + MultLoop_acc_620_itm_1
      + MultLoop_acc_619_itm_1 + MultLoop_acc_616_itm_1 + MultLoop_acc_615_itm_1;
  assign MultLoop_acc_643_nl = nl_MultLoop_acc_643_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1 = (MultLoop_acc_644_nl)
      + (MultLoop_acc_643_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1[21:0];
  assign nl_MultLoop_acc_511_nl = MultLoop_acc_503_itm_1 + MultLoop_acc_502_itm_1;
  assign MultLoop_acc_511_nl = nl_MultLoop_acc_511_nl[21:0];
  assign nl_MultLoop_acc_510_nl = MultLoop_acc_501_itm_1 + MultLoop_acc_500_itm_1;
  assign MultLoop_acc_510_nl = nl_MultLoop_acc_510_nl[21:0];
  assign nl_MultLoop_acc_515_nl = (MultLoop_acc_511_nl) + (MultLoop_acc_510_nl);
  assign MultLoop_acc_515_nl = nl_MultLoop_acc_515_nl[21:0];
  assign nl_MultLoop_acc_514_nl = MultLoop_acc_499_itm_1 + MultLoop_acc_498_itm_1
      + MultLoop_acc_497_itm_1 + MultLoop_acc_496_itm_1;
  assign MultLoop_acc_514_nl = nl_MultLoop_acc_514_nl[21:0];
  assign nl_MultLoop_acc_517_nl = (MultLoop_acc_515_nl) + (MultLoop_acc_514_nl);
  assign MultLoop_acc_517_nl = nl_MultLoop_acc_517_nl[21:0];
  assign nl_MultLoop_acc_516_nl = MultLoop_acc_491_itm_1 + MultLoop_acc_490_itm_1
      + MultLoop_acc_495_itm_1 + MultLoop_acc_494_itm_1 + MultLoop_acc_493_itm_1
      + MultLoop_acc_492_itm_1 + MultLoop_acc_489_itm_1 + MultLoop_acc_488_itm_1;
  assign MultLoop_acc_516_nl = nl_MultLoop_acc_516_nl[21:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1 = (MultLoop_acc_517_nl)
      + (MultLoop_acc_516_nl);
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1[21:0];
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1023:1016]));
  assign MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10239:10232]));
  assign MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9215:9208]));
  assign MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8191:8184]));
  assign MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7167:7160]));
  assign MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6143:6136]));
  assign MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5119:5112]));
  assign MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4095:4088]));
  assign MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3071:3064]));
  assign MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2047:2040]));
  assign MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[20:0]),
      (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nl_AccumDotWidth_acc_2400_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2400_nl = nl_AccumDotWidth_acc_2400_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign nl_AccumDotWidth_acc_2271_nl = conv_s2s_21_22({(AccumDotWidth_acc_2400_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2271_nl = nl_AccumDotWidth_acc_2271_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign nl_AccumDotWidth_acc_2270_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2270_nl = nl_AccumDotWidth_acc_2270_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign nl_AccumDotWidth_acc_2269_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2269_nl = nl_AccumDotWidth_acc_2269_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2271_nl) + (AccumDotWidth_acc_2270_nl) + (AccumDotWidth_acc_2269_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2399_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2399_nl = nl_AccumDotWidth_acc_2399_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign nl_AccumDotWidth_acc_2260_nl = conv_s2s_21_22({(AccumDotWidth_acc_2399_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2260_nl = nl_AccumDotWidth_acc_2260_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign nl_AccumDotWidth_acc_2259_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2259_nl = nl_AccumDotWidth_acc_2259_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign nl_AccumDotWidth_acc_2258_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2258_nl = nl_AccumDotWidth_acc_2258_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2260_nl) + (AccumDotWidth_acc_2259_nl) + (AccumDotWidth_acc_2258_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2398_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2398_nl = nl_AccumDotWidth_acc_2398_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign nl_AccumDotWidth_acc_2249_nl = conv_s2s_21_22({(AccumDotWidth_acc_2398_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2249_nl = nl_AccumDotWidth_acc_2249_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign nl_AccumDotWidth_acc_2248_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2248_nl = nl_AccumDotWidth_acc_2248_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign nl_AccumDotWidth_acc_2247_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2247_nl = nl_AccumDotWidth_acc_2247_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2249_nl) + (AccumDotWidth_acc_2248_nl) + (AccumDotWidth_acc_2247_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2397_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2397_nl = nl_AccumDotWidth_acc_2397_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign nl_AccumDotWidth_acc_2238_nl = conv_s2s_21_22({(AccumDotWidth_acc_2397_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2238_nl = nl_AccumDotWidth_acc_2238_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign nl_AccumDotWidth_acc_2237_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2237_nl = nl_AccumDotWidth_acc_2237_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign nl_AccumDotWidth_acc_2236_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2236_nl = nl_AccumDotWidth_acc_2236_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2238_nl) + (AccumDotWidth_acc_2237_nl) + (AccumDotWidth_acc_2236_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2396_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2396_nl = nl_AccumDotWidth_acc_2396_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign nl_AccumDotWidth_acc_2227_nl = conv_s2s_21_22({(AccumDotWidth_acc_2396_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2227_nl = nl_AccumDotWidth_acc_2227_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign nl_AccumDotWidth_acc_2226_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2226_nl = nl_AccumDotWidth_acc_2226_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign nl_AccumDotWidth_acc_2225_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2225_nl = nl_AccumDotWidth_acc_2225_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2227_nl) + (AccumDotWidth_acc_2226_nl) + (AccumDotWidth_acc_2225_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2395_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2395_nl = nl_AccumDotWidth_acc_2395_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign nl_AccumDotWidth_acc_2216_nl = conv_s2s_21_22({(AccumDotWidth_acc_2395_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2216_nl = nl_AccumDotWidth_acc_2216_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign nl_AccumDotWidth_acc_2215_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2215_nl = nl_AccumDotWidth_acc_2215_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign nl_AccumDotWidth_acc_2214_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2214_nl = nl_AccumDotWidth_acc_2214_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2216_nl) + (AccumDotWidth_acc_2215_nl) + (AccumDotWidth_acc_2214_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2394_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2394_nl = nl_AccumDotWidth_acc_2394_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign nl_AccumDotWidth_acc_2205_nl = conv_s2s_21_22({(AccumDotWidth_acc_2394_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2205_nl = nl_AccumDotWidth_acc_2205_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign nl_AccumDotWidth_acc_2204_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2204_nl = nl_AccumDotWidth_acc_2204_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign nl_AccumDotWidth_acc_2203_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2203_nl = nl_AccumDotWidth_acc_2203_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2205_nl) + (AccumDotWidth_acc_2204_nl) + (AccumDotWidth_acc_2203_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2393_nl = (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2393_nl = nl_AccumDotWidth_acc_2393_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign nl_AccumDotWidth_acc_2194_nl = conv_s2s_21_22({(AccumDotWidth_acc_2393_nl)
      , (ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2194_nl = nl_AccumDotWidth_acc_2194_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign nl_AccumDotWidth_acc_2193_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2193_nl = nl_AccumDotWidth_acc_2193_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign nl_AccumDotWidth_acc_2192_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2192_nl = nl_AccumDotWidth_acc_2192_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2194_nl) + (AccumDotWidth_acc_2193_nl) + (AccumDotWidth_acc_2192_nl);
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2392_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2392_nl = nl_AccumDotWidth_acc_2392_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign nl_AccumDotWidth_acc_2182_nl = conv_s2s_21_22({(AccumDotWidth_acc_2392_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2182_nl = nl_AccumDotWidth_acc_2182_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign nl_AccumDotWidth_acc_2181_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2181_nl = nl_AccumDotWidth_acc_2181_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign nl_AccumDotWidth_acc_2179_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2179_nl = nl_AccumDotWidth_acc_2179_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2182_nl) + (AccumDotWidth_acc_2181_nl) + (AccumDotWidth_acc_2179_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2391_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2391_nl = nl_AccumDotWidth_acc_2391_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign nl_AccumDotWidth_acc_2165_nl = conv_s2s_21_22({(AccumDotWidth_acc_2391_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2165_nl = nl_AccumDotWidth_acc_2165_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign nl_AccumDotWidth_acc_2164_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2164_nl = nl_AccumDotWidth_acc_2164_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign nl_AccumDotWidth_acc_2162_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2162_nl = nl_AccumDotWidth_acc_2162_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2165_nl) + (AccumDotWidth_acc_2164_nl) + (AccumDotWidth_acc_2162_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2390_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2390_nl = nl_AccumDotWidth_acc_2390_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign nl_AccumDotWidth_acc_2148_nl = conv_s2s_21_22({(AccumDotWidth_acc_2390_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2148_nl = nl_AccumDotWidth_acc_2148_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign nl_AccumDotWidth_acc_2147_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2147_nl = nl_AccumDotWidth_acc_2147_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign nl_AccumDotWidth_acc_2145_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2145_nl = nl_AccumDotWidth_acc_2145_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2148_nl) + (AccumDotWidth_acc_2147_nl) + (AccumDotWidth_acc_2145_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2389_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2389_nl = nl_AccumDotWidth_acc_2389_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign nl_AccumDotWidth_acc_2131_nl = conv_s2s_21_22({(AccumDotWidth_acc_2389_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2131_nl = nl_AccumDotWidth_acc_2131_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign nl_AccumDotWidth_acc_2130_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2130_nl = nl_AccumDotWidth_acc_2130_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign nl_AccumDotWidth_acc_2128_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2128_nl = nl_AccumDotWidth_acc_2128_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2131_nl) + (AccumDotWidth_acc_2130_nl) + (AccumDotWidth_acc_2128_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2388_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2388_nl = nl_AccumDotWidth_acc_2388_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign nl_AccumDotWidth_acc_2114_nl = conv_s2s_21_22({(AccumDotWidth_acc_2388_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2114_nl = nl_AccumDotWidth_acc_2114_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign nl_AccumDotWidth_acc_2113_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2113_nl = nl_AccumDotWidth_acc_2113_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign nl_AccumDotWidth_acc_2111_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2111_nl = nl_AccumDotWidth_acc_2111_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2114_nl) + (AccumDotWidth_acc_2113_nl) + (AccumDotWidth_acc_2111_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2387_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2387_nl = nl_AccumDotWidth_acc_2387_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign nl_AccumDotWidth_acc_2097_nl = conv_s2s_21_22({(AccumDotWidth_acc_2387_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2097_nl = nl_AccumDotWidth_acc_2097_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign nl_AccumDotWidth_acc_2096_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2096_nl = nl_AccumDotWidth_acc_2096_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign nl_AccumDotWidth_acc_2094_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2094_nl = nl_AccumDotWidth_acc_2094_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2097_nl) + (AccumDotWidth_acc_2096_nl) + (AccumDotWidth_acc_2094_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2386_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2386_nl = nl_AccumDotWidth_acc_2386_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign nl_AccumDotWidth_acc_2080_nl = conv_s2s_21_22({(AccumDotWidth_acc_2386_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2080_nl = nl_AccumDotWidth_acc_2080_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign nl_AccumDotWidth_acc_2079_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2079_nl = nl_AccumDotWidth_acc_2079_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign nl_AccumDotWidth_acc_2077_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2077_nl = nl_AccumDotWidth_acc_2077_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2080_nl) + (AccumDotWidth_acc_2079_nl) + (AccumDotWidth_acc_2077_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2385_nl = (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2385_nl = nl_AccumDotWidth_acc_2385_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign nl_AccumDotWidth_acc_2063_nl = conv_s2s_21_22({(AccumDotWidth_acc_2385_nl)
      , (ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2063_nl = nl_AccumDotWidth_acc_2063_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign nl_AccumDotWidth_acc_2062_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2062_nl = nl_AccumDotWidth_acc_2062_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign nl_AccumDotWidth_acc_2060_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2060_nl = nl_AccumDotWidth_acc_2060_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2063_nl) + (AccumDotWidth_acc_2062_nl) + (AccumDotWidth_acc_2060_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2384_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2384_nl = nl_AccumDotWidth_acc_2384_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign nl_AccumDotWidth_acc_2046_nl = conv_s2s_21_22({(AccumDotWidth_acc_2384_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2046_nl = nl_AccumDotWidth_acc_2046_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign nl_AccumDotWidth_acc_2045_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2045_nl = nl_AccumDotWidth_acc_2045_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign nl_AccumDotWidth_acc_2043_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2043_nl = nl_AccumDotWidth_acc_2043_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2046_nl) + (AccumDotWidth_acc_2045_nl) + (AccumDotWidth_acc_2043_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2383_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2383_nl = nl_AccumDotWidth_acc_2383_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign nl_AccumDotWidth_acc_2029_nl = conv_s2s_21_22({(AccumDotWidth_acc_2383_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2029_nl = nl_AccumDotWidth_acc_2029_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign nl_AccumDotWidth_acc_2028_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2028_nl = nl_AccumDotWidth_acc_2028_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign nl_AccumDotWidth_acc_2026_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2026_nl = nl_AccumDotWidth_acc_2026_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2029_nl) + (AccumDotWidth_acc_2028_nl) + (AccumDotWidth_acc_2026_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2382_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2382_nl = nl_AccumDotWidth_acc_2382_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign nl_AccumDotWidth_acc_2012_nl = conv_s2s_21_22({(AccumDotWidth_acc_2382_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2012_nl = nl_AccumDotWidth_acc_2012_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign nl_AccumDotWidth_acc_2011_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_2011_nl = nl_AccumDotWidth_acc_2011_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign nl_AccumDotWidth_acc_2009_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_2009_nl = nl_AccumDotWidth_acc_2009_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_2012_nl) + (AccumDotWidth_acc_2011_nl) + (AccumDotWidth_acc_2009_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2381_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2381_nl = nl_AccumDotWidth_acc_2381_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign nl_AccumDotWidth_acc_1995_nl = conv_s2s_21_22({(AccumDotWidth_acc_2381_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1995_nl = nl_AccumDotWidth_acc_1995_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign nl_AccumDotWidth_acc_1994_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1994_nl = nl_AccumDotWidth_acc_1994_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign nl_AccumDotWidth_acc_1992_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1992_nl = nl_AccumDotWidth_acc_1992_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1995_nl) + (AccumDotWidth_acc_1994_nl) + (AccumDotWidth_acc_1992_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2380_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2380_nl = nl_AccumDotWidth_acc_2380_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign nl_AccumDotWidth_acc_1978_nl = conv_s2s_21_22({(AccumDotWidth_acc_2380_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1978_nl = nl_AccumDotWidth_acc_1978_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign nl_AccumDotWidth_acc_1977_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1977_nl = nl_AccumDotWidth_acc_1977_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign nl_AccumDotWidth_acc_1975_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1975_nl = nl_AccumDotWidth_acc_1975_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1978_nl) + (AccumDotWidth_acc_1977_nl) + (AccumDotWidth_acc_1975_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2379_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2379_nl = nl_AccumDotWidth_acc_2379_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign nl_AccumDotWidth_acc_1961_nl = conv_s2s_21_22({(AccumDotWidth_acc_2379_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1961_nl = nl_AccumDotWidth_acc_1961_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign nl_AccumDotWidth_acc_1960_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1960_nl = nl_AccumDotWidth_acc_1960_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign nl_AccumDotWidth_acc_1958_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1958_nl = nl_AccumDotWidth_acc_1958_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1961_nl) + (AccumDotWidth_acc_1960_nl) + (AccumDotWidth_acc_1958_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2378_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2378_nl = nl_AccumDotWidth_acc_2378_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign nl_AccumDotWidth_acc_1944_nl = conv_s2s_21_22({(AccumDotWidth_acc_2378_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1944_nl = nl_AccumDotWidth_acc_1944_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign nl_AccumDotWidth_acc_1943_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1943_nl = nl_AccumDotWidth_acc_1943_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign nl_AccumDotWidth_acc_1941_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1941_nl = nl_AccumDotWidth_acc_1941_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1944_nl) + (AccumDotWidth_acc_1943_nl) + (AccumDotWidth_acc_1941_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2377_nl = (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2377_nl = nl_AccumDotWidth_acc_2377_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign nl_AccumDotWidth_acc_1927_nl = conv_s2s_21_22({(AccumDotWidth_acc_2377_nl)
      , (ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1927_nl = nl_AccumDotWidth_acc_1927_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign nl_AccumDotWidth_acc_1926_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1926_nl = nl_AccumDotWidth_acc_1926_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign nl_AccumDotWidth_acc_1924_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1924_nl = nl_AccumDotWidth_acc_1924_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1927_nl) + (AccumDotWidth_acc_1926_nl) + (AccumDotWidth_acc_1924_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2376_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2376_nl = nl_AccumDotWidth_acc_2376_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign nl_AccumDotWidth_acc_1911_nl = conv_s2s_21_22({(AccumDotWidth_acc_2376_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1911_nl = nl_AccumDotWidth_acc_1911_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign nl_AccumDotWidth_acc_1910_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1910_nl = nl_AccumDotWidth_acc_1910_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign nl_AccumDotWidth_acc_1909_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1909_nl = nl_AccumDotWidth_acc_1909_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1911_nl) + (AccumDotWidth_acc_1910_nl) + (AccumDotWidth_acc_1909_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2375_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2375_nl = nl_AccumDotWidth_acc_2375_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign nl_AccumDotWidth_acc_1900_nl = conv_s2s_21_22({(AccumDotWidth_acc_2375_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1900_nl = nl_AccumDotWidth_acc_1900_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign nl_AccumDotWidth_acc_1899_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1899_nl = nl_AccumDotWidth_acc_1899_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign nl_AccumDotWidth_acc_1898_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1898_nl = nl_AccumDotWidth_acc_1898_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1900_nl) + (AccumDotWidth_acc_1899_nl) + (AccumDotWidth_acc_1898_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2374_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2374_nl = nl_AccumDotWidth_acc_2374_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign nl_AccumDotWidth_acc_1889_nl = conv_s2s_21_22({(AccumDotWidth_acc_2374_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1889_nl = nl_AccumDotWidth_acc_1889_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign nl_AccumDotWidth_acc_1888_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1888_nl = nl_AccumDotWidth_acc_1888_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign nl_AccumDotWidth_acc_1887_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1887_nl = nl_AccumDotWidth_acc_1887_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1889_nl) + (AccumDotWidth_acc_1888_nl) + (AccumDotWidth_acc_1887_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2373_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2373_nl = nl_AccumDotWidth_acc_2373_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign nl_AccumDotWidth_acc_1878_nl = conv_s2s_21_22({(AccumDotWidth_acc_2373_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1878_nl = nl_AccumDotWidth_acc_1878_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign nl_AccumDotWidth_acc_1877_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1877_nl = nl_AccumDotWidth_acc_1877_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign nl_AccumDotWidth_acc_1876_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1876_nl = nl_AccumDotWidth_acc_1876_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1878_nl) + (AccumDotWidth_acc_1877_nl) + (AccumDotWidth_acc_1876_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2372_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2372_nl = nl_AccumDotWidth_acc_2372_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign nl_AccumDotWidth_acc_1867_nl = conv_s2s_21_22({(AccumDotWidth_acc_2372_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1867_nl = nl_AccumDotWidth_acc_1867_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign nl_AccumDotWidth_acc_1866_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1866_nl = nl_AccumDotWidth_acc_1866_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign nl_AccumDotWidth_acc_1865_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1865_nl = nl_AccumDotWidth_acc_1865_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1867_nl) + (AccumDotWidth_acc_1866_nl) + (AccumDotWidth_acc_1865_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2371_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2371_nl = nl_AccumDotWidth_acc_2371_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign nl_AccumDotWidth_acc_1856_nl = conv_s2s_21_22({(AccumDotWidth_acc_2371_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1856_nl = nl_AccumDotWidth_acc_1856_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign nl_AccumDotWidth_acc_1855_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1855_nl = nl_AccumDotWidth_acc_1855_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign nl_AccumDotWidth_acc_1854_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1854_nl = nl_AccumDotWidth_acc_1854_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1856_nl) + (AccumDotWidth_acc_1855_nl) + (AccumDotWidth_acc_1854_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2370_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2370_nl = nl_AccumDotWidth_acc_2370_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign nl_AccumDotWidth_acc_1845_nl = conv_s2s_21_22({(AccumDotWidth_acc_2370_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1845_nl = nl_AccumDotWidth_acc_1845_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign nl_AccumDotWidth_acc_1844_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1844_nl = nl_AccumDotWidth_acc_1844_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign nl_AccumDotWidth_acc_1843_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1843_nl = nl_AccumDotWidth_acc_1843_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1845_nl) + (AccumDotWidth_acc_1844_nl) + (AccumDotWidth_acc_1843_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2369_nl = (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2369_nl = nl_AccumDotWidth_acc_2369_nl[9:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign nl_AccumDotWidth_acc_1834_nl = conv_s2s_21_22({(AccumDotWidth_acc_2369_nl)
      , (ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1834_nl = nl_AccumDotWidth_acc_1834_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign nl_AccumDotWidth_acc_1833_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1833_nl = nl_AccumDotWidth_acc_1833_nl[21:0];
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign nl_AccumDotWidth_acc_1832_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1832_nl = nl_AccumDotWidth_acc_1832_nl[21:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1834_nl) + (AccumDotWidth_acc_1833_nl) + (AccumDotWidth_acc_1832_nl);
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2368_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2368_nl = nl_AccumDotWidth_acc_2368_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign nl_AccumDotWidth_acc_1822_nl = conv_s2s_21_22({(AccumDotWidth_acc_2368_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1822_nl = nl_AccumDotWidth_acc_1822_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign nl_AccumDotWidth_acc_1821_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1821_nl = nl_AccumDotWidth_acc_1821_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign nl_AccumDotWidth_acc_1819_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1819_nl = nl_AccumDotWidth_acc_1819_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1822_nl) + (AccumDotWidth_acc_1821_nl) + (AccumDotWidth_acc_1819_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2367_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2367_nl = nl_AccumDotWidth_acc_2367_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign nl_AccumDotWidth_acc_1805_nl = conv_s2s_21_22({(AccumDotWidth_acc_2367_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1805_nl = nl_AccumDotWidth_acc_1805_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign nl_AccumDotWidth_acc_1804_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1804_nl = nl_AccumDotWidth_acc_1804_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign nl_AccumDotWidth_acc_1802_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1802_nl = nl_AccumDotWidth_acc_1802_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1805_nl) + (AccumDotWidth_acc_1804_nl) + (AccumDotWidth_acc_1802_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2366_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2366_nl = nl_AccumDotWidth_acc_2366_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign nl_AccumDotWidth_acc_1788_nl = conv_s2s_21_22({(AccumDotWidth_acc_2366_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1788_nl = nl_AccumDotWidth_acc_1788_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign nl_AccumDotWidth_acc_1787_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1787_nl = nl_AccumDotWidth_acc_1787_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign nl_AccumDotWidth_acc_1785_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1785_nl = nl_AccumDotWidth_acc_1785_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1788_nl) + (AccumDotWidth_acc_1787_nl) + (AccumDotWidth_acc_1785_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2365_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2365_nl = nl_AccumDotWidth_acc_2365_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign nl_AccumDotWidth_acc_1771_nl = conv_s2s_21_22({(AccumDotWidth_acc_2365_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1771_nl = nl_AccumDotWidth_acc_1771_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign nl_AccumDotWidth_acc_1770_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1770_nl = nl_AccumDotWidth_acc_1770_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign nl_AccumDotWidth_acc_1768_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1768_nl = nl_AccumDotWidth_acc_1768_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1771_nl) + (AccumDotWidth_acc_1770_nl) + (AccumDotWidth_acc_1768_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2364_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2364_nl = nl_AccumDotWidth_acc_2364_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign nl_AccumDotWidth_acc_1754_nl = conv_s2s_21_22({(AccumDotWidth_acc_2364_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1754_nl = nl_AccumDotWidth_acc_1754_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign nl_AccumDotWidth_acc_1753_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1753_nl = nl_AccumDotWidth_acc_1753_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign nl_AccumDotWidth_acc_1751_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1751_nl = nl_AccumDotWidth_acc_1751_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1754_nl) + (AccumDotWidth_acc_1753_nl) + (AccumDotWidth_acc_1751_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2363_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2363_nl = nl_AccumDotWidth_acc_2363_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign nl_AccumDotWidth_acc_1737_nl = conv_s2s_21_22({(AccumDotWidth_acc_2363_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1737_nl = nl_AccumDotWidth_acc_1737_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign nl_AccumDotWidth_acc_1736_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1736_nl = nl_AccumDotWidth_acc_1736_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign nl_AccumDotWidth_acc_1734_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1734_nl = nl_AccumDotWidth_acc_1734_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1737_nl) + (AccumDotWidth_acc_1736_nl) + (AccumDotWidth_acc_1734_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2362_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2362_nl = nl_AccumDotWidth_acc_2362_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign nl_AccumDotWidth_acc_1720_nl = conv_s2s_21_22({(AccumDotWidth_acc_2362_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1720_nl = nl_AccumDotWidth_acc_1720_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign nl_AccumDotWidth_acc_1719_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1719_nl = nl_AccumDotWidth_acc_1719_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign nl_AccumDotWidth_acc_1717_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1717_nl = nl_AccumDotWidth_acc_1717_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1720_nl) + (AccumDotWidth_acc_1719_nl) + (AccumDotWidth_acc_1717_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2361_nl = (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2361_nl = nl_AccumDotWidth_acc_2361_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign nl_AccumDotWidth_acc_1703_nl = conv_s2s_21_22({(AccumDotWidth_acc_2361_nl)
      , (ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1703_nl = nl_AccumDotWidth_acc_1703_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign nl_AccumDotWidth_acc_1702_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1702_nl = nl_AccumDotWidth_acc_1702_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign nl_AccumDotWidth_acc_1700_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1700_nl = nl_AccumDotWidth_acc_1700_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1703_nl) + (AccumDotWidth_acc_1702_nl) + (AccumDotWidth_acc_1700_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumDotWidth_acc_1681_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1681_nl = nl_AccumDotWidth_acc_1681_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_1686_nl = (AccumDotWidth_acc_1681_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1686_nl = nl_AccumDotWidth_acc_1686_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_1679_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1679_nl = nl_AccumDotWidth_acc_1679_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign nl_AccumDotWidth_acc_1685_nl = (AccumDotWidth_acc_1679_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1685_nl = nl_AccumDotWidth_acc_1685_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign nl_AccumDotWidth_acc_1683_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1683_nl = nl_AccumDotWidth_acc_1683_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign nl_AccumDotWidth_acc_1678_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1678_nl = nl_AccumDotWidth_acc_1678_nl[21:0];
  assign nl_AccumDotWidth_acc_2360_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2360_nl = nl_AccumDotWidth_acc_2360_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_1677_nl = conv_s2s_21_22({(AccumDotWidth_acc_2360_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1677_nl = nl_AccumDotWidth_acc_1677_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1686_nl) + (AccumDotWidth_acc_1685_nl) + (AccumDotWidth_acc_1683_nl)
      + (AccumDotWidth_acc_1678_nl) + (AccumDotWidth_acc_1677_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumDotWidth_acc_1655_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1655_nl = nl_AccumDotWidth_acc_1655_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_1660_nl = (AccumDotWidth_acc_1655_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1660_nl = nl_AccumDotWidth_acc_1660_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_1653_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1653_nl = nl_AccumDotWidth_acc_1653_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign nl_AccumDotWidth_acc_1659_nl = (AccumDotWidth_acc_1653_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1659_nl = nl_AccumDotWidth_acc_1659_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign nl_AccumDotWidth_acc_1657_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1657_nl = nl_AccumDotWidth_acc_1657_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign nl_AccumDotWidth_acc_1652_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1652_nl = nl_AccumDotWidth_acc_1652_nl[21:0];
  assign nl_AccumDotWidth_acc_2359_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2359_nl = nl_AccumDotWidth_acc_2359_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_1651_nl = conv_s2s_21_22({(AccumDotWidth_acc_2359_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1651_nl = nl_AccumDotWidth_acc_1651_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1660_nl) + (AccumDotWidth_acc_1659_nl) + (AccumDotWidth_acc_1657_nl)
      + (AccumDotWidth_acc_1652_nl) + (AccumDotWidth_acc_1651_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumDotWidth_acc_1629_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1629_nl = nl_AccumDotWidth_acc_1629_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_1634_nl = (AccumDotWidth_acc_1629_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1634_nl = nl_AccumDotWidth_acc_1634_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_1627_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1627_nl = nl_AccumDotWidth_acc_1627_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign nl_AccumDotWidth_acc_1633_nl = (AccumDotWidth_acc_1627_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1633_nl = nl_AccumDotWidth_acc_1633_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign nl_AccumDotWidth_acc_1631_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1631_nl = nl_AccumDotWidth_acc_1631_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign nl_AccumDotWidth_acc_1626_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1626_nl = nl_AccumDotWidth_acc_1626_nl[21:0];
  assign nl_AccumDotWidth_acc_2358_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2358_nl = nl_AccumDotWidth_acc_2358_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_1625_nl = conv_s2s_21_22({(AccumDotWidth_acc_2358_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1625_nl = nl_AccumDotWidth_acc_1625_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1634_nl) + (AccumDotWidth_acc_1633_nl) + (AccumDotWidth_acc_1631_nl)
      + (AccumDotWidth_acc_1626_nl) + (AccumDotWidth_acc_1625_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumDotWidth_acc_1603_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1603_nl = nl_AccumDotWidth_acc_1603_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_1608_nl = (AccumDotWidth_acc_1603_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1608_nl = nl_AccumDotWidth_acc_1608_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_1601_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1601_nl = nl_AccumDotWidth_acc_1601_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign nl_AccumDotWidth_acc_1607_nl = (AccumDotWidth_acc_1601_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1607_nl = nl_AccumDotWidth_acc_1607_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign nl_AccumDotWidth_acc_1605_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1605_nl = nl_AccumDotWidth_acc_1605_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign nl_AccumDotWidth_acc_1600_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1600_nl = nl_AccumDotWidth_acc_1600_nl[21:0];
  assign nl_AccumDotWidth_acc_2357_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2357_nl = nl_AccumDotWidth_acc_2357_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_1599_nl = conv_s2s_21_22({(AccumDotWidth_acc_2357_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1599_nl = nl_AccumDotWidth_acc_1599_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1608_nl) + (AccumDotWidth_acc_1607_nl) + (AccumDotWidth_acc_1605_nl)
      + (AccumDotWidth_acc_1600_nl) + (AccumDotWidth_acc_1599_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumDotWidth_acc_1577_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1577_nl = nl_AccumDotWidth_acc_1577_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_1582_nl = (AccumDotWidth_acc_1577_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1582_nl = nl_AccumDotWidth_acc_1582_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_1575_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1575_nl = nl_AccumDotWidth_acc_1575_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign nl_AccumDotWidth_acc_1581_nl = (AccumDotWidth_acc_1575_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1581_nl = nl_AccumDotWidth_acc_1581_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign nl_AccumDotWidth_acc_1579_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1579_nl = nl_AccumDotWidth_acc_1579_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign nl_AccumDotWidth_acc_1574_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1574_nl = nl_AccumDotWidth_acc_1574_nl[21:0];
  assign nl_AccumDotWidth_acc_2356_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2356_nl = nl_AccumDotWidth_acc_2356_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_1573_nl = conv_s2s_21_22({(AccumDotWidth_acc_2356_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1573_nl = nl_AccumDotWidth_acc_1573_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1582_nl) + (AccumDotWidth_acc_1581_nl) + (AccumDotWidth_acc_1579_nl)
      + (AccumDotWidth_acc_1574_nl) + (AccumDotWidth_acc_1573_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumDotWidth_acc_1551_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1551_nl = nl_AccumDotWidth_acc_1551_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_1556_nl = (AccumDotWidth_acc_1551_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1556_nl = nl_AccumDotWidth_acc_1556_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_1549_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1549_nl = nl_AccumDotWidth_acc_1549_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign nl_AccumDotWidth_acc_1555_nl = (AccumDotWidth_acc_1549_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1555_nl = nl_AccumDotWidth_acc_1555_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign nl_AccumDotWidth_acc_1553_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1553_nl = nl_AccumDotWidth_acc_1553_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign nl_AccumDotWidth_acc_1548_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1548_nl = nl_AccumDotWidth_acc_1548_nl[21:0];
  assign nl_AccumDotWidth_acc_2355_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2355_nl = nl_AccumDotWidth_acc_2355_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_1547_nl = conv_s2s_21_22({(AccumDotWidth_acc_2355_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1547_nl = nl_AccumDotWidth_acc_1547_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1556_nl) + (AccumDotWidth_acc_1555_nl) + (AccumDotWidth_acc_1553_nl)
      + (AccumDotWidth_acc_1548_nl) + (AccumDotWidth_acc_1547_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumDotWidth_acc_1525_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1525_nl = nl_AccumDotWidth_acc_1525_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_1530_nl = (AccumDotWidth_acc_1525_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1530_nl = nl_AccumDotWidth_acc_1530_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_1523_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1523_nl = nl_AccumDotWidth_acc_1523_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign nl_AccumDotWidth_acc_1529_nl = (AccumDotWidth_acc_1523_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1529_nl = nl_AccumDotWidth_acc_1529_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign nl_AccumDotWidth_acc_1527_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1527_nl = nl_AccumDotWidth_acc_1527_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign nl_AccumDotWidth_acc_1522_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1522_nl = nl_AccumDotWidth_acc_1522_nl[21:0];
  assign nl_AccumDotWidth_acc_2354_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2354_nl = nl_AccumDotWidth_acc_2354_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_1521_nl = conv_s2s_21_22({(AccumDotWidth_acc_2354_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1521_nl = nl_AccumDotWidth_acc_1521_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1530_nl) + (AccumDotWidth_acc_1529_nl) + (AccumDotWidth_acc_1527_nl)
      + (AccumDotWidth_acc_1522_nl) + (AccumDotWidth_acc_1521_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1011:990])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumDotWidth_acc_1499_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1499_nl = nl_AccumDotWidth_acc_1499_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_1504_nl = (AccumDotWidth_acc_1499_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1504_nl = nl_AccumDotWidth_acc_1504_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1033:1012])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_1497_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1497_nl = nl_AccumDotWidth_acc_1497_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign nl_AccumDotWidth_acc_1503_nl = (AccumDotWidth_acc_1497_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1503_nl = nl_AccumDotWidth_acc_1503_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign nl_AccumDotWidth_acc_1501_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1501_nl = nl_AccumDotWidth_acc_1501_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign nl_AccumDotWidth_acc_1496_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1496_nl = nl_AccumDotWidth_acc_1496_nl[21:0];
  assign nl_AccumDotWidth_acc_2353_nl = (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2353_nl = nl_AccumDotWidth_acc_2353_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_1495_nl = conv_s2s_21_22({(AccumDotWidth_acc_2353_nl)
      , (ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1495_nl = nl_AccumDotWidth_acc_1495_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1504_nl) + (AccumDotWidth_acc_1503_nl) + (AccumDotWidth_acc_1501_nl)
      + (AccumDotWidth_acc_1496_nl) + (AccumDotWidth_acc_1495_nl);
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumDotWidth_acc_1473_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1473_nl = nl_AccumDotWidth_acc_1473_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_1478_nl = (AccumDotWidth_acc_1473_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1478_nl = nl_AccumDotWidth_acc_1478_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_1471_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1471_nl = nl_AccumDotWidth_acc_1471_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign nl_AccumDotWidth_acc_1477_nl = (AccumDotWidth_acc_1471_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1477_nl = nl_AccumDotWidth_acc_1477_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign nl_AccumDotWidth_acc_1475_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1475_nl = nl_AccumDotWidth_acc_1475_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign nl_AccumDotWidth_acc_1470_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1470_nl = nl_AccumDotWidth_acc_1470_nl[21:0];
  assign nl_AccumDotWidth_acc_2352_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2352_nl = nl_AccumDotWidth_acc_2352_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_1469_nl = conv_s2s_21_22({(AccumDotWidth_acc_2352_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1469_nl = nl_AccumDotWidth_acc_1469_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1478_nl) + (AccumDotWidth_acc_1477_nl) + (AccumDotWidth_acc_1475_nl)
      + (AccumDotWidth_acc_1470_nl) + (AccumDotWidth_acc_1469_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumDotWidth_acc_1447_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1447_nl = nl_AccumDotWidth_acc_1447_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_1452_nl = (AccumDotWidth_acc_1447_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1452_nl = nl_AccumDotWidth_acc_1452_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_1445_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1445_nl = nl_AccumDotWidth_acc_1445_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign nl_AccumDotWidth_acc_1451_nl = (AccumDotWidth_acc_1445_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1451_nl = nl_AccumDotWidth_acc_1451_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign nl_AccumDotWidth_acc_1449_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1449_nl = nl_AccumDotWidth_acc_1449_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign nl_AccumDotWidth_acc_1444_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1444_nl = nl_AccumDotWidth_acc_1444_nl[21:0];
  assign nl_AccumDotWidth_acc_2351_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2351_nl = nl_AccumDotWidth_acc_2351_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_1443_nl = conv_s2s_21_22({(AccumDotWidth_acc_2351_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1443_nl = nl_AccumDotWidth_acc_1443_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1452_nl) + (AccumDotWidth_acc_1451_nl) + (AccumDotWidth_acc_1449_nl)
      + (AccumDotWidth_acc_1444_nl) + (AccumDotWidth_acc_1443_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumDotWidth_acc_1421_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1421_nl = nl_AccumDotWidth_acc_1421_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_1426_nl = (AccumDotWidth_acc_1421_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1426_nl = nl_AccumDotWidth_acc_1426_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_1419_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1419_nl = nl_AccumDotWidth_acc_1419_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign nl_AccumDotWidth_acc_1425_nl = (AccumDotWidth_acc_1419_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1425_nl = nl_AccumDotWidth_acc_1425_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign nl_AccumDotWidth_acc_1423_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1423_nl = nl_AccumDotWidth_acc_1423_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign nl_AccumDotWidth_acc_1418_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1418_nl = nl_AccumDotWidth_acc_1418_nl[21:0];
  assign nl_AccumDotWidth_acc_2350_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2350_nl = nl_AccumDotWidth_acc_2350_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_1417_nl = conv_s2s_21_22({(AccumDotWidth_acc_2350_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1417_nl = nl_AccumDotWidth_acc_1417_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1426_nl) + (AccumDotWidth_acc_1425_nl) + (AccumDotWidth_acc_1423_nl)
      + (AccumDotWidth_acc_1418_nl) + (AccumDotWidth_acc_1417_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumDotWidth_acc_1395_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1395_nl = nl_AccumDotWidth_acc_1395_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_1400_nl = (AccumDotWidth_acc_1395_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1400_nl = nl_AccumDotWidth_acc_1400_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_1393_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1393_nl = nl_AccumDotWidth_acc_1393_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign nl_AccumDotWidth_acc_1399_nl = (AccumDotWidth_acc_1393_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1399_nl = nl_AccumDotWidth_acc_1399_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign nl_AccumDotWidth_acc_1397_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1397_nl = nl_AccumDotWidth_acc_1397_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign nl_AccumDotWidth_acc_1392_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1392_nl = nl_AccumDotWidth_acc_1392_nl[21:0];
  assign nl_AccumDotWidth_acc_2349_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2349_nl = nl_AccumDotWidth_acc_2349_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_1391_nl = conv_s2s_21_22({(AccumDotWidth_acc_2349_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1391_nl = nl_AccumDotWidth_acc_1391_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1400_nl) + (AccumDotWidth_acc_1399_nl) + (AccumDotWidth_acc_1397_nl)
      + (AccumDotWidth_acc_1392_nl) + (AccumDotWidth_acc_1391_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumDotWidth_acc_1369_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1369_nl = nl_AccumDotWidth_acc_1369_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_1374_nl = (AccumDotWidth_acc_1369_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1374_nl = nl_AccumDotWidth_acc_1374_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_1367_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1367_nl = nl_AccumDotWidth_acc_1367_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign nl_AccumDotWidth_acc_1373_nl = (AccumDotWidth_acc_1367_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1373_nl = nl_AccumDotWidth_acc_1373_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign nl_AccumDotWidth_acc_1371_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1371_nl = nl_AccumDotWidth_acc_1371_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign nl_AccumDotWidth_acc_1366_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1366_nl = nl_AccumDotWidth_acc_1366_nl[21:0];
  assign nl_AccumDotWidth_acc_2348_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2348_nl = nl_AccumDotWidth_acc_2348_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_1365_nl = conv_s2s_21_22({(AccumDotWidth_acc_2348_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1365_nl = nl_AccumDotWidth_acc_1365_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1374_nl) + (AccumDotWidth_acc_1373_nl) + (AccumDotWidth_acc_1371_nl)
      + (AccumDotWidth_acc_1366_nl) + (AccumDotWidth_acc_1365_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumDotWidth_acc_1343_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1343_nl = nl_AccumDotWidth_acc_1343_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_1348_nl = (AccumDotWidth_acc_1343_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1348_nl = nl_AccumDotWidth_acc_1348_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_1341_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1341_nl = nl_AccumDotWidth_acc_1341_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign nl_AccumDotWidth_acc_1347_nl = (AccumDotWidth_acc_1341_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1347_nl = nl_AccumDotWidth_acc_1347_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign nl_AccumDotWidth_acc_1345_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1345_nl = nl_AccumDotWidth_acc_1345_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign nl_AccumDotWidth_acc_1340_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1340_nl = nl_AccumDotWidth_acc_1340_nl[21:0];
  assign nl_AccumDotWidth_acc_2347_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2347_nl = nl_AccumDotWidth_acc_2347_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_1339_nl = conv_s2s_21_22({(AccumDotWidth_acc_2347_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1339_nl = nl_AccumDotWidth_acc_1339_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1348_nl) + (AccumDotWidth_acc_1347_nl) + (AccumDotWidth_acc_1345_nl)
      + (AccumDotWidth_acc_1340_nl) + (AccumDotWidth_acc_1339_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumDotWidth_acc_1317_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1317_nl = nl_AccumDotWidth_acc_1317_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_1322_nl = (AccumDotWidth_acc_1317_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1322_nl = nl_AccumDotWidth_acc_1322_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_1315_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1315_nl = nl_AccumDotWidth_acc_1315_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign nl_AccumDotWidth_acc_1321_nl = (AccumDotWidth_acc_1315_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1321_nl = nl_AccumDotWidth_acc_1321_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign nl_AccumDotWidth_acc_1319_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1319_nl = nl_AccumDotWidth_acc_1319_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign nl_AccumDotWidth_acc_1314_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1314_nl = nl_AccumDotWidth_acc_1314_nl[21:0];
  assign nl_AccumDotWidth_acc_2346_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2346_nl = nl_AccumDotWidth_acc_2346_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_1313_nl = conv_s2s_21_22({(AccumDotWidth_acc_2346_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1313_nl = nl_AccumDotWidth_acc_1313_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1322_nl) + (AccumDotWidth_acc_1321_nl) + (AccumDotWidth_acc_1319_nl)
      + (AccumDotWidth_acc_1314_nl) + (AccumDotWidth_acc_1313_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[945:924])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumDotWidth_acc_1291_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1291_nl = nl_AccumDotWidth_acc_1291_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_1296_nl = (AccumDotWidth_acc_1291_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1296_nl = nl_AccumDotWidth_acc_1296_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[967:946])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_1289_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1289_nl = nl_AccumDotWidth_acc_1289_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign nl_AccumDotWidth_acc_1295_nl = (AccumDotWidth_acc_1289_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1295_nl = nl_AccumDotWidth_acc_1295_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign nl_AccumDotWidth_acc_1293_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1293_nl = nl_AccumDotWidth_acc_1293_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign nl_AccumDotWidth_acc_1288_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_1288_nl = nl_AccumDotWidth_acc_1288_nl[21:0];
  assign nl_AccumDotWidth_acc_2345_nl = (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2345_nl = nl_AccumDotWidth_acc_2345_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_1287_nl = conv_s2s_21_22({(AccumDotWidth_acc_2345_nl)
      , (ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1287_nl = nl_AccumDotWidth_acc_1287_nl[21:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1296_nl) + (AccumDotWidth_acc_1295_nl) + (AccumDotWidth_acc_1293_nl)
      + (AccumDotWidth_acc_1288_nl) + (AccumDotWidth_acc_1287_nl);
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2344_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2344_nl = nl_AccumDotWidth_acc_2344_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_1270_nl = conv_s2s_21_22({(AccumDotWidth_acc_2344_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1270_nl = nl_AccumDotWidth_acc_1270_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_1269_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1269_nl = nl_AccumDotWidth_acc_1269_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_1267_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1267_nl = nl_AccumDotWidth_acc_1267_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1270_nl) + (AccumDotWidth_acc_1269_nl) + (AccumDotWidth_acc_1267_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2343_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2343_nl = nl_AccumDotWidth_acc_2343_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_1253_nl = conv_s2s_21_22({(AccumDotWidth_acc_2343_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1253_nl = nl_AccumDotWidth_acc_1253_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_1252_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1252_nl = nl_AccumDotWidth_acc_1252_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_1250_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1250_nl = nl_AccumDotWidth_acc_1250_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1253_nl) + (AccumDotWidth_acc_1252_nl) + (AccumDotWidth_acc_1250_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2342_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2342_nl = nl_AccumDotWidth_acc_2342_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_1236_nl = conv_s2s_21_22({(AccumDotWidth_acc_2342_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1236_nl = nl_AccumDotWidth_acc_1236_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_1235_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1235_nl = nl_AccumDotWidth_acc_1235_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_1233_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1233_nl = nl_AccumDotWidth_acc_1233_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1236_nl) + (AccumDotWidth_acc_1235_nl) + (AccumDotWidth_acc_1233_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2341_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2341_nl = nl_AccumDotWidth_acc_2341_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_1219_nl = conv_s2s_21_22({(AccumDotWidth_acc_2341_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1219_nl = nl_AccumDotWidth_acc_1219_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_1218_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1218_nl = nl_AccumDotWidth_acc_1218_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_1216_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1216_nl = nl_AccumDotWidth_acc_1216_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1219_nl) + (AccumDotWidth_acc_1218_nl) + (AccumDotWidth_acc_1216_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2340_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2340_nl = nl_AccumDotWidth_acc_2340_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_1202_nl = conv_s2s_21_22({(AccumDotWidth_acc_2340_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1202_nl = nl_AccumDotWidth_acc_1202_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_1201_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1201_nl = nl_AccumDotWidth_acc_1201_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_1199_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1199_nl = nl_AccumDotWidth_acc_1199_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1202_nl) + (AccumDotWidth_acc_1201_nl) + (AccumDotWidth_acc_1199_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2339_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2339_nl = nl_AccumDotWidth_acc_2339_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_1185_nl = conv_s2s_21_22({(AccumDotWidth_acc_2339_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1185_nl = nl_AccumDotWidth_acc_1185_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_1184_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1184_nl = nl_AccumDotWidth_acc_1184_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_1182_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1182_nl = nl_AccumDotWidth_acc_1182_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1185_nl) + (AccumDotWidth_acc_1184_nl) + (AccumDotWidth_acc_1182_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2338_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2338_nl = nl_AccumDotWidth_acc_2338_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_1168_nl = conv_s2s_21_22({(AccumDotWidth_acc_2338_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1168_nl = nl_AccumDotWidth_acc_1168_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_1167_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1167_nl = nl_AccumDotWidth_acc_1167_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_1165_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1165_nl = nl_AccumDotWidth_acc_1165_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1168_nl) + (AccumDotWidth_acc_1167_nl) + (AccumDotWidth_acc_1165_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2337_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2337_nl = nl_AccumDotWidth_acc_2337_nl[9:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[857:836])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_1151_nl = conv_s2s_21_22({(AccumDotWidth_acc_2337_nl)
      , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1151_nl = nl_AccumDotWidth_acc_1151_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[813:792])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_1150_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1150_nl = nl_AccumDotWidth_acc_1150_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[835:814])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[901:880])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_1148_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_1148_nl = nl_AccumDotWidth_acc_1148_nl[21:0];
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[879:858])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (AccumDotWidth_acc_1151_nl) + (AccumDotWidth_acc_1150_nl) + (AccumDotWidth_acc_1148_nl)
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2336_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2336_nl = nl_AccumDotWidth_acc_2336_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign nl_AccumDotWidth_acc_1134_nl = conv_s2s_21_22({(AccumDotWidth_acc_2336_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1134_nl = nl_AccumDotWidth_acc_1134_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign nl_AccumDotWidth_acc_1133_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1133_nl = nl_AccumDotWidth_acc_1133_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign nl_AccumDotWidth_acc_1131_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1131_nl = nl_AccumDotWidth_acc_1131_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1 = (AccumDotWidth_acc_1134_nl)
      + (AccumDotWidth_acc_1133_nl) + (AccumDotWidth_acc_1131_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2335_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2335_nl = nl_AccumDotWidth_acc_2335_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign nl_AccumDotWidth_acc_1117_nl = conv_s2s_21_22({(AccumDotWidth_acc_2335_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1117_nl = nl_AccumDotWidth_acc_1117_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign nl_AccumDotWidth_acc_1116_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1116_nl = nl_AccumDotWidth_acc_1116_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign nl_AccumDotWidth_acc_1114_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1114_nl = nl_AccumDotWidth_acc_1114_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1 = (AccumDotWidth_acc_1117_nl)
      + (AccumDotWidth_acc_1116_nl) + (AccumDotWidth_acc_1114_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2334_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2334_nl = nl_AccumDotWidth_acc_2334_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign nl_AccumDotWidth_acc_1100_nl = conv_s2s_21_22({(AccumDotWidth_acc_2334_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1100_nl = nl_AccumDotWidth_acc_1100_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign nl_AccumDotWidth_acc_1099_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1099_nl = nl_AccumDotWidth_acc_1099_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign nl_AccumDotWidth_acc_1097_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1097_nl = nl_AccumDotWidth_acc_1097_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1 = (AccumDotWidth_acc_1100_nl)
      + (AccumDotWidth_acc_1099_nl) + (AccumDotWidth_acc_1097_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2333_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2333_nl = nl_AccumDotWidth_acc_2333_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign nl_AccumDotWidth_acc_1083_nl = conv_s2s_21_22({(AccumDotWidth_acc_2333_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1083_nl = nl_AccumDotWidth_acc_1083_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign nl_AccumDotWidth_acc_1082_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1082_nl = nl_AccumDotWidth_acc_1082_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign nl_AccumDotWidth_acc_1080_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1080_nl = nl_AccumDotWidth_acc_1080_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = (AccumDotWidth_acc_1083_nl)
      + (AccumDotWidth_acc_1082_nl) + (AccumDotWidth_acc_1080_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2332_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2332_nl = nl_AccumDotWidth_acc_2332_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign nl_AccumDotWidth_acc_1066_nl = conv_s2s_21_22({(AccumDotWidth_acc_2332_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1066_nl = nl_AccumDotWidth_acc_1066_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign nl_AccumDotWidth_acc_1065_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1065_nl = nl_AccumDotWidth_acc_1065_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign nl_AccumDotWidth_acc_1063_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1063_nl = nl_AccumDotWidth_acc_1063_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = (AccumDotWidth_acc_1066_nl)
      + (AccumDotWidth_acc_1065_nl) + (AccumDotWidth_acc_1063_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2331_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2331_nl = nl_AccumDotWidth_acc_2331_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign nl_AccumDotWidth_acc_1049_nl = conv_s2s_21_22({(AccumDotWidth_acc_2331_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1049_nl = nl_AccumDotWidth_acc_1049_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign nl_AccumDotWidth_acc_1048_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1048_nl = nl_AccumDotWidth_acc_1048_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign nl_AccumDotWidth_acc_1046_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1046_nl = nl_AccumDotWidth_acc_1046_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1 = (AccumDotWidth_acc_1049_nl)
      + (AccumDotWidth_acc_1048_nl) + (AccumDotWidth_acc_1046_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2330_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2330_nl = nl_AccumDotWidth_acc_2330_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign nl_AccumDotWidth_acc_1032_nl = conv_s2s_21_22({(AccumDotWidth_acc_2330_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1032_nl = nl_AccumDotWidth_acc_1032_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign nl_AccumDotWidth_acc_1031_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1031_nl = nl_AccumDotWidth_acc_1031_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign nl_AccumDotWidth_acc_1029_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1029_nl = nl_AccumDotWidth_acc_1029_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1 = (AccumDotWidth_acc_1032_nl)
      + (AccumDotWidth_acc_1031_nl) + (AccumDotWidth_acc_1029_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2329_nl = (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2329_nl = nl_AccumDotWidth_acc_2329_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign nl_AccumDotWidth_acc_1015_nl = conv_s2s_21_22({(AccumDotWidth_acc_2329_nl)
      , (ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1015_nl = nl_AccumDotWidth_acc_1015_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign nl_AccumDotWidth_acc_1014_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1014_nl = nl_AccumDotWidth_acc_1014_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign nl_AccumDotWidth_acc_1012_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_1012_nl = nl_AccumDotWidth_acc_1012_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1 = (AccumDotWidth_acc_1015_nl)
      + (AccumDotWidth_acc_1014_nl) + (AccumDotWidth_acc_1012_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumDotWidth_acc_993_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_993_nl = nl_AccumDotWidth_acc_993_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_998_nl = (AccumDotWidth_acc_993_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_998_nl = nl_AccumDotWidth_acc_998_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_991_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_991_nl = nl_AccumDotWidth_acc_991_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign nl_AccumDotWidth_acc_997_nl = (AccumDotWidth_acc_991_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_997_nl = nl_AccumDotWidth_acc_997_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign nl_AccumDotWidth_acc_995_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_995_nl = nl_AccumDotWidth_acc_995_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign nl_AccumDotWidth_acc_990_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_990_nl = nl_AccumDotWidth_acc_990_nl[21:0];
  assign nl_AccumDotWidth_acc_2328_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2328_nl = nl_AccumDotWidth_acc_2328_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_989_nl = conv_s2s_21_22({(AccumDotWidth_acc_2328_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_989_nl = nl_AccumDotWidth_acc_989_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1 = (AccumDotWidth_acc_998_nl)
      + (AccumDotWidth_acc_997_nl) + (AccumDotWidth_acc_995_nl) + (AccumDotWidth_acc_990_nl)
      + (AccumDotWidth_acc_989_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumDotWidth_acc_967_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_967_nl = nl_AccumDotWidth_acc_967_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_972_nl = (AccumDotWidth_acc_967_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_972_nl = nl_AccumDotWidth_acc_972_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_965_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_965_nl = nl_AccumDotWidth_acc_965_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign nl_AccumDotWidth_acc_971_nl = (AccumDotWidth_acc_965_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_971_nl = nl_AccumDotWidth_acc_971_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign nl_AccumDotWidth_acc_969_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_969_nl = nl_AccumDotWidth_acc_969_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign nl_AccumDotWidth_acc_964_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_964_nl = nl_AccumDotWidth_acc_964_nl[21:0];
  assign nl_AccumDotWidth_acc_2327_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2327_nl = nl_AccumDotWidth_acc_2327_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_963_nl = conv_s2s_21_22({(AccumDotWidth_acc_2327_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_963_nl = nl_AccumDotWidth_acc_963_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1 = (AccumDotWidth_acc_972_nl)
      + (AccumDotWidth_acc_971_nl) + (AccumDotWidth_acc_969_nl) + (AccumDotWidth_acc_964_nl)
      + (AccumDotWidth_acc_963_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumDotWidth_acc_941_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_941_nl = nl_AccumDotWidth_acc_941_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_946_nl = (AccumDotWidth_acc_941_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_946_nl = nl_AccumDotWidth_acc_946_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_939_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_939_nl = nl_AccumDotWidth_acc_939_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign nl_AccumDotWidth_acc_945_nl = (AccumDotWidth_acc_939_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_945_nl = nl_AccumDotWidth_acc_945_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign nl_AccumDotWidth_acc_943_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_943_nl = nl_AccumDotWidth_acc_943_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign nl_AccumDotWidth_acc_938_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_938_nl = nl_AccumDotWidth_acc_938_nl[21:0];
  assign nl_AccumDotWidth_acc_2326_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2326_nl = nl_AccumDotWidth_acc_2326_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_937_nl = conv_s2s_21_22({(AccumDotWidth_acc_2326_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_937_nl = nl_AccumDotWidth_acc_937_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1 = (AccumDotWidth_acc_946_nl)
      + (AccumDotWidth_acc_945_nl) + (AccumDotWidth_acc_943_nl) + (AccumDotWidth_acc_938_nl)
      + (AccumDotWidth_acc_937_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumDotWidth_acc_915_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_915_nl = nl_AccumDotWidth_acc_915_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_920_nl = (AccumDotWidth_acc_915_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_920_nl = nl_AccumDotWidth_acc_920_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_913_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_913_nl = nl_AccumDotWidth_acc_913_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign nl_AccumDotWidth_acc_919_nl = (AccumDotWidth_acc_913_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_919_nl = nl_AccumDotWidth_acc_919_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign nl_AccumDotWidth_acc_917_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_917_nl = nl_AccumDotWidth_acc_917_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign nl_AccumDotWidth_acc_912_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_912_nl = nl_AccumDotWidth_acc_912_nl[21:0];
  assign nl_AccumDotWidth_acc_2325_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2325_nl = nl_AccumDotWidth_acc_2325_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_911_nl = conv_s2s_21_22({(AccumDotWidth_acc_2325_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_911_nl = nl_AccumDotWidth_acc_911_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1 = (AccumDotWidth_acc_920_nl)
      + (AccumDotWidth_acc_919_nl) + (AccumDotWidth_acc_917_nl) + (AccumDotWidth_acc_912_nl)
      + (AccumDotWidth_acc_911_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumDotWidth_acc_889_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_889_nl = nl_AccumDotWidth_acc_889_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_894_nl = (AccumDotWidth_acc_889_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_894_nl = nl_AccumDotWidth_acc_894_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_887_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_887_nl = nl_AccumDotWidth_acc_887_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign nl_AccumDotWidth_acc_893_nl = (AccumDotWidth_acc_887_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_893_nl = nl_AccumDotWidth_acc_893_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign nl_AccumDotWidth_acc_891_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_891_nl = nl_AccumDotWidth_acc_891_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign nl_AccumDotWidth_acc_886_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_886_nl = nl_AccumDotWidth_acc_886_nl[21:0];
  assign nl_AccumDotWidth_acc_2324_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2324_nl = nl_AccumDotWidth_acc_2324_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_885_nl = conv_s2s_21_22({(AccumDotWidth_acc_2324_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_885_nl = nl_AccumDotWidth_acc_885_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1 = (AccumDotWidth_acc_894_nl)
      + (AccumDotWidth_acc_893_nl) + (AccumDotWidth_acc_891_nl) + (AccumDotWidth_acc_886_nl)
      + (AccumDotWidth_acc_885_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumDotWidth_acc_863_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_863_nl = nl_AccumDotWidth_acc_863_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_868_nl = (AccumDotWidth_acc_863_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_868_nl = nl_AccumDotWidth_acc_868_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_861_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_861_nl = nl_AccumDotWidth_acc_861_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign nl_AccumDotWidth_acc_867_nl = (AccumDotWidth_acc_861_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_867_nl = nl_AccumDotWidth_acc_867_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign nl_AccumDotWidth_acc_865_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_865_nl = nl_AccumDotWidth_acc_865_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign nl_AccumDotWidth_acc_860_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_860_nl = nl_AccumDotWidth_acc_860_nl[21:0];
  assign nl_AccumDotWidth_acc_2323_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2323_nl = nl_AccumDotWidth_acc_2323_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_859_nl = conv_s2s_21_22({(AccumDotWidth_acc_2323_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_859_nl = nl_AccumDotWidth_acc_859_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1 = (AccumDotWidth_acc_868_nl)
      + (AccumDotWidth_acc_867_nl) + (AccumDotWidth_acc_865_nl) + (AccumDotWidth_acc_860_nl)
      + (AccumDotWidth_acc_859_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumDotWidth_acc_837_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_837_nl = nl_AccumDotWidth_acc_837_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_842_nl = (AccumDotWidth_acc_837_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_842_nl = nl_AccumDotWidth_acc_842_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_835_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_835_nl = nl_AccumDotWidth_acc_835_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign nl_AccumDotWidth_acc_841_nl = (AccumDotWidth_acc_835_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_841_nl = nl_AccumDotWidth_acc_841_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign nl_AccumDotWidth_acc_839_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_839_nl = nl_AccumDotWidth_acc_839_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign nl_AccumDotWidth_acc_834_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_834_nl = nl_AccumDotWidth_acc_834_nl[21:0];
  assign nl_AccumDotWidth_acc_2322_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2322_nl = nl_AccumDotWidth_acc_2322_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_833_nl = conv_s2s_21_22({(AccumDotWidth_acc_2322_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_833_nl = nl_AccumDotWidth_acc_833_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1 = (AccumDotWidth_acc_842_nl)
      + (AccumDotWidth_acc_841_nl) + (AccumDotWidth_acc_839_nl) + (AccumDotWidth_acc_834_nl)
      + (AccumDotWidth_acc_833_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[747:726])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumDotWidth_acc_811_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_811_nl = nl_AccumDotWidth_acc_811_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_816_nl = (AccumDotWidth_acc_811_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_816_nl = nl_AccumDotWidth_acc_816_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[769:748])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_809_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_809_nl = nl_AccumDotWidth_acc_809_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign nl_AccumDotWidth_acc_815_nl = (AccumDotWidth_acc_809_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_815_nl = nl_AccumDotWidth_acc_815_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign nl_AccumDotWidth_acc_813_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_813_nl = nl_AccumDotWidth_acc_813_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign nl_AccumDotWidth_acc_808_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_808_nl = nl_AccumDotWidth_acc_808_nl[21:0];
  assign nl_AccumDotWidth_acc_2321_nl = (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2321_nl = nl_AccumDotWidth_acc_2321_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_807_nl = conv_s2s_21_22({(AccumDotWidth_acc_2321_nl)
      , (ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_807_nl = nl_AccumDotWidth_acc_807_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1 = (AccumDotWidth_acc_816_nl)
      + (AccumDotWidth_acc_815_nl) + (AccumDotWidth_acc_813_nl) + (AccumDotWidth_acc_808_nl)
      + (AccumDotWidth_acc_807_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[127:120])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign nl_AccumDotWidth_acc_785_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_785_nl = nl_AccumDotWidth_acc_785_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_790_nl = (AccumDotWidth_acc_785_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_790_nl = nl_AccumDotWidth_acc_790_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[191:184])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_783_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_783_nl = nl_AccumDotWidth_acc_783_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign nl_AccumDotWidth_acc_789_nl = (AccumDotWidth_acc_783_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_789_nl = nl_AccumDotWidth_acc_789_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[63:56])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign nl_AccumDotWidth_acc_787_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_787_nl = nl_AccumDotWidth_acc_787_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign nl_AccumDotWidth_acc_782_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_782_nl = nl_AccumDotWidth_acc_782_nl[21:0];
  assign nl_AccumDotWidth_acc_2320_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2320_nl = nl_AccumDotWidth_acc_2320_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_781_nl = conv_s2s_21_22({(AccumDotWidth_acc_2320_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_781_nl = nl_AccumDotWidth_acc_781_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1 = (AccumDotWidth_acc_790_nl)
      + (AccumDotWidth_acc_789_nl) + (AccumDotWidth_acc_787_nl) + (AccumDotWidth_acc_782_nl)
      + (AccumDotWidth_acc_781_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[119:112])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign nl_AccumDotWidth_acc_759_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_759_nl = nl_AccumDotWidth_acc_759_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_764_nl = (AccumDotWidth_acc_759_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_764_nl = nl_AccumDotWidth_acc_764_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[183:176])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_757_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_757_nl = nl_AccumDotWidth_acc_757_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign nl_AccumDotWidth_acc_763_nl = (AccumDotWidth_acc_757_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_763_nl = nl_AccumDotWidth_acc_763_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[55:48])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign nl_AccumDotWidth_acc_761_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_761_nl = nl_AccumDotWidth_acc_761_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign nl_AccumDotWidth_acc_756_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_756_nl = nl_AccumDotWidth_acc_756_nl[21:0];
  assign nl_AccumDotWidth_acc_2319_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2319_nl = nl_AccumDotWidth_acc_2319_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_755_nl = conv_s2s_21_22({(AccumDotWidth_acc_2319_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_755_nl = nl_AccumDotWidth_acc_755_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1 = (AccumDotWidth_acc_764_nl)
      + (AccumDotWidth_acc_763_nl) + (AccumDotWidth_acc_761_nl) + (AccumDotWidth_acc_756_nl)
      + (AccumDotWidth_acc_755_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[111:104])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign nl_AccumDotWidth_acc_733_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_733_nl = nl_AccumDotWidth_acc_733_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_738_nl = (AccumDotWidth_acc_733_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_738_nl = nl_AccumDotWidth_acc_738_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[175:168])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_731_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_731_nl = nl_AccumDotWidth_acc_731_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign nl_AccumDotWidth_acc_737_nl = (AccumDotWidth_acc_731_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_737_nl = nl_AccumDotWidth_acc_737_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[47:40])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign nl_AccumDotWidth_acc_735_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_735_nl = nl_AccumDotWidth_acc_735_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign nl_AccumDotWidth_acc_730_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_730_nl = nl_AccumDotWidth_acc_730_nl[21:0];
  assign nl_AccumDotWidth_acc_2318_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2318_nl = nl_AccumDotWidth_acc_2318_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_729_nl = conv_s2s_21_22({(AccumDotWidth_acc_2318_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_729_nl = nl_AccumDotWidth_acc_729_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1 = (AccumDotWidth_acc_738_nl)
      + (AccumDotWidth_acc_737_nl) + (AccumDotWidth_acc_735_nl) + (AccumDotWidth_acc_730_nl)
      + (AccumDotWidth_acc_729_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[103:96])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign nl_AccumDotWidth_acc_707_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_707_nl = nl_AccumDotWidth_acc_707_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_712_nl = (AccumDotWidth_acc_707_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_712_nl = nl_AccumDotWidth_acc_712_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[167:160])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_705_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_705_nl = nl_AccumDotWidth_acc_705_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign nl_AccumDotWidth_acc_711_nl = (AccumDotWidth_acc_705_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_711_nl = nl_AccumDotWidth_acc_711_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[39:32])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign nl_AccumDotWidth_acc_709_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_709_nl = nl_AccumDotWidth_acc_709_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign nl_AccumDotWidth_acc_704_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_704_nl = nl_AccumDotWidth_acc_704_nl[21:0];
  assign nl_AccumDotWidth_acc_2317_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2317_nl = nl_AccumDotWidth_acc_2317_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_703_nl = conv_s2s_21_22({(AccumDotWidth_acc_2317_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_703_nl = nl_AccumDotWidth_acc_703_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1 = (AccumDotWidth_acc_712_nl)
      + (AccumDotWidth_acc_711_nl) + (AccumDotWidth_acc_709_nl) + (AccumDotWidth_acc_704_nl)
      + (AccumDotWidth_acc_703_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[95:88])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign nl_AccumDotWidth_acc_681_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_681_nl = nl_AccumDotWidth_acc_681_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_686_nl = (AccumDotWidth_acc_681_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_686_nl = nl_AccumDotWidth_acc_686_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[159:152])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_679_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_679_nl = nl_AccumDotWidth_acc_679_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign nl_AccumDotWidth_acc_685_nl = (AccumDotWidth_acc_679_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_685_nl = nl_AccumDotWidth_acc_685_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[31:24])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign nl_AccumDotWidth_acc_683_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_683_nl = nl_AccumDotWidth_acc_683_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign nl_AccumDotWidth_acc_678_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_678_nl = nl_AccumDotWidth_acc_678_nl[21:0];
  assign nl_AccumDotWidth_acc_2316_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2316_nl = nl_AccumDotWidth_acc_2316_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_677_nl = conv_s2s_21_22({(AccumDotWidth_acc_2316_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_677_nl = nl_AccumDotWidth_acc_677_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1 = (AccumDotWidth_acc_686_nl)
      + (AccumDotWidth_acc_685_nl) + (AccumDotWidth_acc_683_nl) + (AccumDotWidth_acc_678_nl)
      + (AccumDotWidth_acc_677_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[87:80])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign nl_AccumDotWidth_acc_655_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_655_nl = nl_AccumDotWidth_acc_655_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_660_nl = (AccumDotWidth_acc_655_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_660_nl = nl_AccumDotWidth_acc_660_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[151:144])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_653_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_653_nl = nl_AccumDotWidth_acc_653_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign nl_AccumDotWidth_acc_659_nl = (AccumDotWidth_acc_653_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_659_nl = nl_AccumDotWidth_acc_659_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[23:16])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign nl_AccumDotWidth_acc_657_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_657_nl = nl_AccumDotWidth_acc_657_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign nl_AccumDotWidth_acc_652_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_652_nl = nl_AccumDotWidth_acc_652_nl[21:0];
  assign nl_AccumDotWidth_acc_2315_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2315_nl = nl_AccumDotWidth_acc_2315_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_651_nl = conv_s2s_21_22({(AccumDotWidth_acc_2315_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_651_nl = nl_AccumDotWidth_acc_651_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1 = (AccumDotWidth_acc_660_nl)
      + (AccumDotWidth_acc_659_nl) + (AccumDotWidth_acc_657_nl) + (AccumDotWidth_acc_652_nl)
      + (AccumDotWidth_acc_651_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[79:72])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign nl_AccumDotWidth_acc_629_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_629_nl = nl_AccumDotWidth_acc_629_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_634_nl = (AccumDotWidth_acc_629_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_634_nl = nl_AccumDotWidth_acc_634_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[143:136])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_627_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_627_nl = nl_AccumDotWidth_acc_627_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign nl_AccumDotWidth_acc_633_nl = (AccumDotWidth_acc_627_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_633_nl = nl_AccumDotWidth_acc_633_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[15:8])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign nl_AccumDotWidth_acc_631_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_631_nl = nl_AccumDotWidth_acc_631_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign nl_AccumDotWidth_acc_626_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_626_nl = nl_AccumDotWidth_acc_626_nl[21:0];
  assign nl_AccumDotWidth_acc_2314_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2314_nl = nl_AccumDotWidth_acc_2314_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_625_nl = conv_s2s_21_22({(AccumDotWidth_acc_2314_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_625_nl = nl_AccumDotWidth_acc_625_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1 = (AccumDotWidth_acc_634_nl)
      + (AccumDotWidth_acc_633_nl) + (AccumDotWidth_acc_631_nl) + (AccumDotWidth_acc_626_nl)
      + (AccumDotWidth_acc_625_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[681:660])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[71:64])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign nl_AccumDotWidth_acc_603_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_603_nl = nl_AccumDotWidth_acc_603_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_608_nl = (AccumDotWidth_acc_603_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_608_nl = nl_AccumDotWidth_acc_608_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[703:682])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[135:128])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_601_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_601_nl = nl_AccumDotWidth_acc_601_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign nl_AccumDotWidth_acc_607_nl = (AccumDotWidth_acc_601_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_607_nl = nl_AccumDotWidth_acc_607_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[7:0])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign nl_AccumDotWidth_acc_605_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_605_nl = nl_AccumDotWidth_acc_605_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign nl_AccumDotWidth_acc_600_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign AccumDotWidth_acc_600_nl = nl_AccumDotWidth_acc_600_nl[21:0];
  assign nl_AccumDotWidth_acc_2313_nl = (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2313_nl = nl_AccumDotWidth_acc_2313_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_599_nl = conv_s2s_21_22({(AccumDotWidth_acc_2313_nl)
      , (ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_599_nl = nl_AccumDotWidth_acc_599_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1 = (AccumDotWidth_acc_608_nl)
      + (AccumDotWidth_acc_607_nl) + (AccumDotWidth_acc_605_nl) + (AccumDotWidth_acc_600_nl)
      + (AccumDotWidth_acc_599_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2312_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2312_nl = nl_AccumDotWidth_acc_2312_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[255:248])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[575:568])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_582_nl = conv_s2s_21_22({(AccumDotWidth_acc_2312_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_582_nl = nl_AccumDotWidth_acc_582_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[447:440])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_581_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_581_nl = nl_AccumDotWidth_acc_581_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[383:376])));
  assign nl_AccumDotWidth_acc_579_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_579_nl = nl_AccumDotWidth_acc_579_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[319:312])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[511:504])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1 = (AccumDotWidth_acc_582_nl)
      + (AccumDotWidth_acc_581_nl) + (AccumDotWidth_acc_579_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2311_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2311_nl = nl_AccumDotWidth_acc_2311_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[247:240])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[567:560])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_565_nl = conv_s2s_21_22({(AccumDotWidth_acc_2311_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_565_nl = nl_AccumDotWidth_acc_565_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[439:432])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_564_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_564_nl = nl_AccumDotWidth_acc_564_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[375:368])));
  assign nl_AccumDotWidth_acc_562_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_562_nl = nl_AccumDotWidth_acc_562_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[311:304])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[503:496])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1 = (AccumDotWidth_acc_565_nl)
      + (AccumDotWidth_acc_564_nl) + (AccumDotWidth_acc_562_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2310_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2310_nl = nl_AccumDotWidth_acc_2310_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[239:232])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[559:552])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_548_nl = conv_s2s_21_22({(AccumDotWidth_acc_2310_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_548_nl = nl_AccumDotWidth_acc_548_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[431:424])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_547_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_547_nl = nl_AccumDotWidth_acc_547_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[367:360])));
  assign nl_AccumDotWidth_acc_545_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_545_nl = nl_AccumDotWidth_acc_545_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[303:296])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[495:488])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1 = (AccumDotWidth_acc_548_nl)
      + (AccumDotWidth_acc_547_nl) + (AccumDotWidth_acc_545_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2309_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2309_nl = nl_AccumDotWidth_acc_2309_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[231:224])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[551:544])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_531_nl = conv_s2s_21_22({(AccumDotWidth_acc_2309_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_531_nl = nl_AccumDotWidth_acc_531_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[423:416])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_530_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_530_nl = nl_AccumDotWidth_acc_530_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[359:352])));
  assign nl_AccumDotWidth_acc_528_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_528_nl = nl_AccumDotWidth_acc_528_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[295:288])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[487:480])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1 = (AccumDotWidth_acc_531_nl)
      + (AccumDotWidth_acc_530_nl) + (AccumDotWidth_acc_528_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2308_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2308_nl = nl_AccumDotWidth_acc_2308_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[223:216])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[543:536])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_514_nl = conv_s2s_21_22({(AccumDotWidth_acc_2308_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_514_nl = nl_AccumDotWidth_acc_514_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[415:408])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_513_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_513_nl = nl_AccumDotWidth_acc_513_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[351:344])));
  assign nl_AccumDotWidth_acc_511_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_511_nl = nl_AccumDotWidth_acc_511_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[287:280])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[479:472])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1 = (AccumDotWidth_acc_514_nl)
      + (AccumDotWidth_acc_513_nl) + (AccumDotWidth_acc_511_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2307_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2307_nl = nl_AccumDotWidth_acc_2307_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[215:208])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[535:528])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_497_nl = conv_s2s_21_22({(AccumDotWidth_acc_2307_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_497_nl = nl_AccumDotWidth_acc_497_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[407:400])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_496_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_496_nl = nl_AccumDotWidth_acc_496_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[343:336])));
  assign nl_AccumDotWidth_acc_494_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_494_nl = nl_AccumDotWidth_acc_494_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[279:272])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[471:464])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1 = (AccumDotWidth_acc_497_nl)
      + (AccumDotWidth_acc_496_nl) + (AccumDotWidth_acc_494_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2306_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2306_nl = nl_AccumDotWidth_acc_2306_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[207:200])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[527:520])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_480_nl = conv_s2s_21_22({(AccumDotWidth_acc_2306_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_480_nl = nl_AccumDotWidth_acc_480_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[399:392])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_479_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_479_nl = nl_AccumDotWidth_acc_479_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[335:328])));
  assign nl_AccumDotWidth_acc_477_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_477_nl = nl_AccumDotWidth_acc_477_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[271:264])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[463:456])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1 = (AccumDotWidth_acc_480_nl)
      + (AccumDotWidth_acc_479_nl) + (AccumDotWidth_acc_477_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2305_nl = (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2305_nl = nl_AccumDotWidth_acc_2305_nl[9:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[199:192])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[519:512])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[593:572])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_463_nl = conv_s2s_21_22({(AccumDotWidth_acc_2305_nl)
      , (ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_463_nl = nl_AccumDotWidth_acc_463_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[391:384])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[549:528])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_462_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_462_nl = nl_AccumDotWidth_acc_462_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[571:550])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[637:616])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[327:320])));
  assign nl_AccumDotWidth_acc_460_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_460_nl = nl_AccumDotWidth_acc_460_nl[21:0];
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[615:594])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[263:256])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[455:448])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1 = (AccumDotWidth_acc_463_nl)
      + (AccumDotWidth_acc_462_nl) + (AccumDotWidth_acc_460_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2304_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2304_nl = nl_AccumDotWidth_acc_2304_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign nl_AccumDotWidth_acc_447_nl = conv_s2s_21_22({(AccumDotWidth_acc_2304_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_447_nl = nl_AccumDotWidth_acc_447_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign nl_AccumDotWidth_acc_446_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_446_nl = nl_AccumDotWidth_acc_446_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign nl_AccumDotWidth_acc_445_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_445_nl = nl_AccumDotWidth_acc_445_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1 = (AccumDotWidth_acc_447_nl)
      + (AccumDotWidth_acc_446_nl) + (AccumDotWidth_acc_445_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2303_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2303_nl = nl_AccumDotWidth_acc_2303_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign nl_AccumDotWidth_acc_436_nl = conv_s2s_21_22({(AccumDotWidth_acc_2303_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_436_nl = nl_AccumDotWidth_acc_436_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign nl_AccumDotWidth_acc_435_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_435_nl = nl_AccumDotWidth_acc_435_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign nl_AccumDotWidth_acc_434_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_434_nl = nl_AccumDotWidth_acc_434_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1 = (AccumDotWidth_acc_436_nl)
      + (AccumDotWidth_acc_435_nl) + (AccumDotWidth_acc_434_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2302_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2302_nl = nl_AccumDotWidth_acc_2302_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign nl_AccumDotWidth_acc_425_nl = conv_s2s_21_22({(AccumDotWidth_acc_2302_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_425_nl = nl_AccumDotWidth_acc_425_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign nl_AccumDotWidth_acc_424_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_424_nl = nl_AccumDotWidth_acc_424_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign nl_AccumDotWidth_acc_423_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_423_nl = nl_AccumDotWidth_acc_423_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1 = (AccumDotWidth_acc_425_nl)
      + (AccumDotWidth_acc_424_nl) + (AccumDotWidth_acc_423_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2301_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2301_nl = nl_AccumDotWidth_acc_2301_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign nl_AccumDotWidth_acc_414_nl = conv_s2s_21_22({(AccumDotWidth_acc_2301_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_414_nl = nl_AccumDotWidth_acc_414_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign nl_AccumDotWidth_acc_413_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_413_nl = nl_AccumDotWidth_acc_413_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign nl_AccumDotWidth_acc_412_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_412_nl = nl_AccumDotWidth_acc_412_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1 = (AccumDotWidth_acc_414_nl)
      + (AccumDotWidth_acc_413_nl) + (AccumDotWidth_acc_412_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2300_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2300_nl = nl_AccumDotWidth_acc_2300_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign nl_AccumDotWidth_acc_403_nl = conv_s2s_21_22({(AccumDotWidth_acc_2300_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_403_nl = nl_AccumDotWidth_acc_403_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign nl_AccumDotWidth_acc_402_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_402_nl = nl_AccumDotWidth_acc_402_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign nl_AccumDotWidth_acc_401_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_401_nl = nl_AccumDotWidth_acc_401_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1 = (AccumDotWidth_acc_403_nl)
      + (AccumDotWidth_acc_402_nl) + (AccumDotWidth_acc_401_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2299_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2299_nl = nl_AccumDotWidth_acc_2299_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign nl_AccumDotWidth_acc_392_nl = conv_s2s_21_22({(AccumDotWidth_acc_2299_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_392_nl = nl_AccumDotWidth_acc_392_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign nl_AccumDotWidth_acc_391_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_391_nl = nl_AccumDotWidth_acc_391_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign nl_AccumDotWidth_acc_390_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_390_nl = nl_AccumDotWidth_acc_390_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1 = (AccumDotWidth_acc_392_nl)
      + (AccumDotWidth_acc_391_nl) + (AccumDotWidth_acc_390_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2298_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2298_nl = nl_AccumDotWidth_acc_2298_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign nl_AccumDotWidth_acc_381_nl = conv_s2s_21_22({(AccumDotWidth_acc_2298_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_381_nl = nl_AccumDotWidth_acc_381_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign nl_AccumDotWidth_acc_380_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_380_nl = nl_AccumDotWidth_acc_380_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign nl_AccumDotWidth_acc_379_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_379_nl = nl_AccumDotWidth_acc_379_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1 = (AccumDotWidth_acc_381_nl)
      + (AccumDotWidth_acc_380_nl) + (AccumDotWidth_acc_379_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2297_nl = (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2297_nl = nl_AccumDotWidth_acc_2297_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign nl_AccumDotWidth_acc_370_nl = conv_s2s_21_22({(AccumDotWidth_acc_2297_nl)
      , (ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_370_nl = nl_AccumDotWidth_acc_370_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign nl_AccumDotWidth_acc_369_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_369_nl = nl_AccumDotWidth_acc_369_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign nl_AccumDotWidth_acc_368_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_368_nl = nl_AccumDotWidth_acc_368_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1 = (AccumDotWidth_acc_370_nl)
      + (AccumDotWidth_acc_369_nl) + (AccumDotWidth_acc_368_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2296_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2296_nl = nl_AccumDotWidth_acc_2296_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_358_nl = conv_s2s_21_22({(AccumDotWidth_acc_2296_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_358_nl = nl_AccumDotWidth_acc_358_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_357_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_357_nl = nl_AccumDotWidth_acc_357_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign nl_AccumDotWidth_acc_355_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_355_nl = nl_AccumDotWidth_acc_355_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1 = (AccumDotWidth_acc_358_nl)
      + (AccumDotWidth_acc_357_nl) + (AccumDotWidth_acc_355_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2295_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2295_nl = nl_AccumDotWidth_acc_2295_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_341_nl = conv_s2s_21_22({(AccumDotWidth_acc_2295_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_341_nl = nl_AccumDotWidth_acc_341_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_340_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_340_nl = nl_AccumDotWidth_acc_340_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign nl_AccumDotWidth_acc_338_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_338_nl = nl_AccumDotWidth_acc_338_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1 = (AccumDotWidth_acc_341_nl)
      + (AccumDotWidth_acc_340_nl) + (AccumDotWidth_acc_338_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2294_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2294_nl = nl_AccumDotWidth_acc_2294_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_324_nl = conv_s2s_21_22({(AccumDotWidth_acc_2294_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_324_nl = nl_AccumDotWidth_acc_324_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_323_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_323_nl = nl_AccumDotWidth_acc_323_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign nl_AccumDotWidth_acc_321_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_321_nl = nl_AccumDotWidth_acc_321_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1 = (AccumDotWidth_acc_324_nl)
      + (AccumDotWidth_acc_323_nl) + (AccumDotWidth_acc_321_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2293_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2293_nl = nl_AccumDotWidth_acc_2293_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_307_nl = conv_s2s_21_22({(AccumDotWidth_acc_2293_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_307_nl = nl_AccumDotWidth_acc_307_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_306_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_306_nl = nl_AccumDotWidth_acc_306_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign nl_AccumDotWidth_acc_304_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_304_nl = nl_AccumDotWidth_acc_304_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1 = (AccumDotWidth_acc_307_nl)
      + (AccumDotWidth_acc_306_nl) + (AccumDotWidth_acc_304_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2292_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2292_nl = nl_AccumDotWidth_acc_2292_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_290_nl = conv_s2s_21_22({(AccumDotWidth_acc_2292_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_290_nl = nl_AccumDotWidth_acc_290_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_289_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_289_nl = nl_AccumDotWidth_acc_289_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign nl_AccumDotWidth_acc_287_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_287_nl = nl_AccumDotWidth_acc_287_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1 = (AccumDotWidth_acc_290_nl)
      + (AccumDotWidth_acc_289_nl) + (AccumDotWidth_acc_287_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2291_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2291_nl = nl_AccumDotWidth_acc_2291_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_273_nl = conv_s2s_21_22({(AccumDotWidth_acc_2291_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_273_nl = nl_AccumDotWidth_acc_273_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_272_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_272_nl = nl_AccumDotWidth_acc_272_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign nl_AccumDotWidth_acc_270_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_270_nl = nl_AccumDotWidth_acc_270_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1 = (AccumDotWidth_acc_273_nl)
      + (AccumDotWidth_acc_272_nl) + (AccumDotWidth_acc_270_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2290_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2290_nl = nl_AccumDotWidth_acc_2290_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_256_nl = conv_s2s_21_22({(AccumDotWidth_acc_2290_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_256_nl = nl_AccumDotWidth_acc_256_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_255_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_255_nl = nl_AccumDotWidth_acc_255_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign nl_AccumDotWidth_acc_253_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_253_nl = nl_AccumDotWidth_acc_253_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1 = (AccumDotWidth_acc_256_nl)
      + (AccumDotWidth_acc_255_nl) + (AccumDotWidth_acc_253_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2289_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2289_nl = nl_AccumDotWidth_acc_2289_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[263:242])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_239_nl = conv_s2s_21_22({(AccumDotWidth_acc_2289_nl)
      , (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_239_nl = nl_AccumDotWidth_acc_239_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[219:198])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_238_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_238_nl = nl_AccumDotWidth_acc_238_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[505:484])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign nl_AccumDotWidth_acc_236_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_236_nl = nl_AccumDotWidth_acc_236_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[483:462])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[241:220])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1 = (AccumDotWidth_acc_239_nl)
      + (AccumDotWidth_acc_238_nl) + (AccumDotWidth_acc_236_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2288_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2288_nl = nl_AccumDotWidth_acc_2288_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[639:632])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1343:1336])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_222_nl = conv_s2s_21_22({(AccumDotWidth_acc_2288_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_222_nl = nl_AccumDotWidth_acc_222_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1215:1208])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_221_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_221_nl = nl_AccumDotWidth_acc_221_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1279:1272])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[767:760])));
  assign nl_AccumDotWidth_acc_219_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_219_nl = nl_AccumDotWidth_acc_219_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[703:696])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1 = (AccumDotWidth_acc_222_nl)
      + (AccumDotWidth_acc_221_nl) + (AccumDotWidth_acc_219_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2287_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2287_nl = nl_AccumDotWidth_acc_2287_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[631:624])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1335:1328])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_205_nl = conv_s2s_21_22({(AccumDotWidth_acc_2287_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_205_nl = nl_AccumDotWidth_acc_205_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1207:1200])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_204_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_204_nl = nl_AccumDotWidth_acc_204_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1271:1264])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[759:752])));
  assign nl_AccumDotWidth_acc_202_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_202_nl = nl_AccumDotWidth_acc_202_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[695:688])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1 = (AccumDotWidth_acc_205_nl)
      + (AccumDotWidth_acc_204_nl) + (AccumDotWidth_acc_202_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2286_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2286_nl = nl_AccumDotWidth_acc_2286_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[623:616])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1327:1320])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_188_nl = conv_s2s_21_22({(AccumDotWidth_acc_2286_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_188_nl = nl_AccumDotWidth_acc_188_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1199:1192])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_187_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_187_nl = nl_AccumDotWidth_acc_187_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1263:1256])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[751:744])));
  assign nl_AccumDotWidth_acc_185_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_185_nl = nl_AccumDotWidth_acc_185_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[687:680])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1 = (AccumDotWidth_acc_188_nl)
      + (AccumDotWidth_acc_187_nl) + (AccumDotWidth_acc_185_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2285_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2285_nl = nl_AccumDotWidth_acc_2285_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[615:608])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1319:1312])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_171_nl = conv_s2s_21_22({(AccumDotWidth_acc_2285_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_171_nl = nl_AccumDotWidth_acc_171_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1191:1184])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_170_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_170_nl = nl_AccumDotWidth_acc_170_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1255:1248])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[743:736])));
  assign nl_AccumDotWidth_acc_168_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_168_nl = nl_AccumDotWidth_acc_168_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[679:672])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1 = (AccumDotWidth_acc_171_nl)
      + (AccumDotWidth_acc_170_nl) + (AccumDotWidth_acc_168_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2284_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2284_nl = nl_AccumDotWidth_acc_2284_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[607:600])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1311:1304])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_154_nl = conv_s2s_21_22({(AccumDotWidth_acc_2284_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_154_nl = nl_AccumDotWidth_acc_154_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1183:1176])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_153_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_153_nl = nl_AccumDotWidth_acc_153_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1247:1240])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[735:728])));
  assign nl_AccumDotWidth_acc_151_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_151_nl = nl_AccumDotWidth_acc_151_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[671:664])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1 = (AccumDotWidth_acc_154_nl)
      + (AccumDotWidth_acc_153_nl) + (AccumDotWidth_acc_151_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2283_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2283_nl = nl_AccumDotWidth_acc_2283_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[599:592])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1303:1296])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_137_nl = conv_s2s_21_22({(AccumDotWidth_acc_2283_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_137_nl = nl_AccumDotWidth_acc_137_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1175:1168])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_136_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_136_nl = nl_AccumDotWidth_acc_136_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1239:1232])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[727:720])));
  assign nl_AccumDotWidth_acc_134_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_134_nl = nl_AccumDotWidth_acc_134_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[663:656])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1 = (AccumDotWidth_acc_137_nl)
      + (AccumDotWidth_acc_136_nl) + (AccumDotWidth_acc_134_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2282_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2282_nl = nl_AccumDotWidth_acc_2282_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[591:584])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1295:1288])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_120_nl = conv_s2s_21_22({(AccumDotWidth_acc_2282_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_120_nl = nl_AccumDotWidth_acc_120_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1167:1160])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_119_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_119_nl = nl_AccumDotWidth_acc_119_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1231:1224])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[719:712])));
  assign nl_AccumDotWidth_acc_117_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_117_nl = nl_AccumDotWidth_acc_117_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[655:648])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1 = (AccumDotWidth_acc_120_nl)
      + (AccumDotWidth_acc_119_nl) + (AccumDotWidth_acc_117_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2281_nl = (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2281_nl = nl_AccumDotWidth_acc_2281_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[583:576])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[197:176])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1287:1280])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_103_nl = conv_s2s_21_22({(AccumDotWidth_acc_2281_nl)
      , (ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_103_nl = nl_AccumDotWidth_acc_103_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[153:132])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1159:1152])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_102_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_102_nl = nl_AccumDotWidth_acc_102_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1223:1216])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[439:418])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[711:704])));
  assign nl_AccumDotWidth_acc_100_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)));
  assign AccumDotWidth_acc_100_nl = nl_AccumDotWidth_acc_100_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[417:396])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[647:640])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[175:154])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1 = (AccumDotWidth_acc_103_nl)
      + (AccumDotWidth_acc_102_nl) + (AccumDotWidth_acc_100_nl) + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2280_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2280_nl = nl_AccumDotWidth_acc_2280_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[831:824])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[1023:1016])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1407:1400])));
  assign nl_AccumDotWidth_acc_87_nl = conv_s2s_21_22({(AccumDotWidth_acc_2280_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_87_nl = nl_AccumDotWidth_acc_87_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1599:1592])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[895:888])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1087:1080])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1471:1464])));
  assign nl_AccumDotWidth_acc_86_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_86_nl = nl_AccumDotWidth_acc_86_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1663:1656])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign nl_AccumDotWidth_acc_85_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_85_nl = nl_AccumDotWidth_acc_85_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1 = (AccumDotWidth_acc_87_nl)
      + (AccumDotWidth_acc_86_nl) + (AccumDotWidth_acc_85_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2279_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2279_nl = nl_AccumDotWidth_acc_2279_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[823:816])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[1015:1008])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1399:1392])));
  assign nl_AccumDotWidth_acc_76_nl = conv_s2s_21_22({(AccumDotWidth_acc_2279_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_76_nl = nl_AccumDotWidth_acc_76_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1591:1584])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[887:880])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1079:1072])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1463:1456])));
  assign nl_AccumDotWidth_acc_75_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_75_nl = nl_AccumDotWidth_acc_75_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1655:1648])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign nl_AccumDotWidth_acc_74_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_74_nl = nl_AccumDotWidth_acc_74_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1 = (AccumDotWidth_acc_76_nl)
      + (AccumDotWidth_acc_75_nl) + (AccumDotWidth_acc_74_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2278_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2278_nl = nl_AccumDotWidth_acc_2278_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[815:808])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[1007:1000])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1391:1384])));
  assign nl_AccumDotWidth_acc_65_nl = conv_s2s_21_22({(AccumDotWidth_acc_2278_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_65_nl = nl_AccumDotWidth_acc_65_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1583:1576])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[879:872])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1071:1064])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1455:1448])));
  assign nl_AccumDotWidth_acc_64_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_64_nl = nl_AccumDotWidth_acc_64_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1647:1640])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign nl_AccumDotWidth_acc_63_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_63_nl = nl_AccumDotWidth_acc_63_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1 = (AccumDotWidth_acc_65_nl)
      + (AccumDotWidth_acc_64_nl) + (AccumDotWidth_acc_63_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2277_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2277_nl = nl_AccumDotWidth_acc_2277_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[807:800])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[999:992])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1383:1376])));
  assign nl_AccumDotWidth_acc_54_nl = conv_s2s_21_22({(AccumDotWidth_acc_2277_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_54_nl = nl_AccumDotWidth_acc_54_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1575:1568])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[871:864])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1063:1056])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1447:1440])));
  assign nl_AccumDotWidth_acc_53_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_53_nl = nl_AccumDotWidth_acc_53_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1639:1632])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign nl_AccumDotWidth_acc_52_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_52_nl = nl_AccumDotWidth_acc_52_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1 = (AccumDotWidth_acc_54_nl)
      + (AccumDotWidth_acc_53_nl) + (AccumDotWidth_acc_52_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2276_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[31:24]);
  assign AccumDotWidth_acc_2276_nl = nl_AccumDotWidth_acc_2276_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[799:792])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[991:984])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1375:1368])));
  assign nl_AccumDotWidth_acc_43_nl = conv_s2s_21_22({(AccumDotWidth_acc_2276_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_43_nl = nl_AccumDotWidth_acc_43_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1567:1560])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[863:856])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1055:1048])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1439:1432])));
  assign nl_AccumDotWidth_acc_42_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_42_nl = nl_AccumDotWidth_acc_42_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1631:1624])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign nl_AccumDotWidth_acc_41_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_41_nl = nl_AccumDotWidth_acc_41_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1 = (AccumDotWidth_acc_43_nl)
      + (AccumDotWidth_acc_42_nl) + (AccumDotWidth_acc_41_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2275_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2275_nl = nl_AccumDotWidth_acc_2275_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[791:784])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[983:976])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1367:1360])));
  assign nl_AccumDotWidth_acc_32_nl = conv_s2s_21_22({(AccumDotWidth_acc_2275_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_32_nl = nl_AccumDotWidth_acc_32_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1559:1552])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[855:848])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1047:1040])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1431:1424])));
  assign nl_AccumDotWidth_acc_31_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_31_nl = nl_AccumDotWidth_acc_31_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1623:1616])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign nl_AccumDotWidth_acc_30_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_30_nl = nl_AccumDotWidth_acc_30_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1 = (AccumDotWidth_acc_32_nl)
      + (AccumDotWidth_acc_31_nl) + (AccumDotWidth_acc_30_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2274_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2274_nl = nl_AccumDotWidth_acc_2274_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[783:776])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[975:968])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1359:1352])));
  assign nl_AccumDotWidth_acc_21_nl = conv_s2s_21_22({(AccumDotWidth_acc_2274_nl)
      , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_21_nl = nl_AccumDotWidth_acc_21_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1551:1544])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[847:840])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1039:1032])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1423:1416])));
  assign nl_AccumDotWidth_acc_20_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_20_nl = nl_AccumDotWidth_acc_20_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1615:1608])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign nl_AccumDotWidth_acc_19_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_19_nl = nl_AccumDotWidth_acc_19_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1 = (AccumDotWidth_acc_21_nl)
      + (AccumDotWidth_acc_20_nl) + (AccumDotWidth_acc_19_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1[21:0];
  assign nl_AccumDotWidth_acc_2273_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[20:11])
      + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2273_nl = nl_AccumDotWidth_acc_2273_nl[9:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[21:0])) * $signed((w2_rsci_idat_mxwt[775:768])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[87:66])) * $signed((w2_rsci_idat_mxwt[967:960])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[285:264])) * $signed((w2_rsci_idat_mxwt[1351:1344])));
  assign nl_AccumDotWidth_acc_nl = conv_s2s_21_22({(AccumDotWidth_acc_2273_nl) ,
      (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9[10:0])})
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_nl = nl_AccumDotWidth_acc_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[351:330])) * $signed((w2_rsci_idat_mxwt[1543:1536])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[43:22])) * $signed((w2_rsci_idat_mxwt[839:832])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[109:88])) * $signed((w2_rsci_idat_mxwt[1031:1024])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[307:286])) * $signed((w2_rsci_idat_mxwt[1415:1408])));
  assign nl_AccumDotWidth_acc_9_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_9_nl = nl_AccumDotWidth_acc_9_nl[21:0];
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[373:352])) * $signed((w2_rsci_idat_mxwt[1607:1600])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[65:44])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[131:110])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[329:308])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign nl_AccumDotWidth_acc_8_nl = conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl)))
      + conv_s2s_21_22(readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl)));
  assign AccumDotWidth_acc_8_nl = nl_AccumDotWidth_acc_8_nl[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1 = (AccumDotWidth_acc_nl)
      + (AccumDotWidth_acc_9_nl) + (AccumDotWidth_acc_8_nl);
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1[21:0];
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[959:952])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[951:944])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[943:936])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[935:928])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[927:920])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[919:912])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[911:904])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[903:896])));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1151:1144])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1143:1136])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1135:1128])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1127:1120])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1119:1112])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1111:1104])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1103:1096])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1095:1088])));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[1055:1034])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[989:968])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[923:902])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[791:770])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[725:704])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[659:638])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1535:1528])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1527:1520])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1519:1512])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1511:1504])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1503:1496])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1495:1488])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1487:1480])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1479:1472])));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[527:506])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[461:440])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1727:1720])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1719:1712])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1711:1704])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1703:1696])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1695:1688])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1687:1680])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1679:1672])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = conv_s2u_30_30($signed((input_1_rsci_idat_mxwt[395:374])) * $signed((w2_rsci_idat_mxwt[1671:1664])));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_itm_29_9
      = readslicef_30_21_9((ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289 = MUX_v_21_2_2(21'b000000000000000000000,
      (nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_idat_218_198 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_42_22 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_64_44 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_86_66 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_108_88 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_130_110 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_152_132 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_174_154 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_196_176 <= 21'b000000000000000000000;
    end
    else if ( layer5_out_and_cse ) begin
      layer5_out_rsci_idat_218_198 <= MUX_v_21_2_2(21'b000000000000000000000, (MultLoop_1280_MultLoop_acc_3_ncse_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_20_0 <= MUX_v_21_2_2(21'b000000000000000000000, (layer4_out_0_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_42_22 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_64_44 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_86_66 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_108_88 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_130_110 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_152_132 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_174_154 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_196_176 <= MUX_v_21_2_2(21'b000000000000000000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      MultLoop_acc_1265_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1264_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1263_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1262_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1261_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1260_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1259_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1258_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1257_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1256_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1255_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1254_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1253_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1252_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1251_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1250_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1138_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1137_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1136_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1135_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1134_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1133_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1132_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1131_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1130_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1129_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1128_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1127_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1126_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1125_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1124_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1123_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1011_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1010_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1009_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1008_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1007_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1006_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1005_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1004_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1003_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1002_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1001_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_1000_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_999_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_998_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_997_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_996_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_884_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_883_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_882_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_881_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_880_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_879_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_878_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_877_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_876_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_875_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_874_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_873_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_872_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_871_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_870_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_869_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_757_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_756_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_755_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_754_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_753_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_752_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_751_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_750_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_749_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_748_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_747_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_746_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_745_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_744_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_743_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_742_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_630_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_629_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_628_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_627_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_626_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_625_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_624_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_623_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_622_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_621_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_620_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_619_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_618_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_617_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_616_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_615_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_503_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_502_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_501_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_500_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_499_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_498_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_497_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_496_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_495_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_494_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_493_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_492_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_491_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_490_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_489_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_488_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_376_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_375_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_374_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_373_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_372_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_371_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_370_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_369_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_368_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_367_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_366_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_365_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_364_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_363_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_362_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_361_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_249_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_248_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_247_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_246_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_245_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_244_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_243_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_242_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_241_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_240_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_239_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_238_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_237_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_236_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_235_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_234_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_130_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_121_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_120_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_119_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_118_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_117_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_116_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_115_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_114_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_113_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_112_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_111_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_110_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_109_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_108_itm_1 <= 22'b0000000000000000000000;
      MultLoop_acc_107_itm_1 <= 22'b0000000000000000000000;
      main_stage_0_2 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= 1'b1;
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= main_stage_0_2;
      MultLoop_acc_1265_itm_1 <= nl_MultLoop_acc_1265_itm_1[21:0];
      MultLoop_acc_1264_itm_1 <= nl_MultLoop_acc_1264_itm_1[21:0];
      MultLoop_acc_1263_itm_1 <= nl_MultLoop_acc_1263_itm_1[21:0];
      MultLoop_acc_1262_itm_1 <= nl_MultLoop_acc_1262_itm_1[21:0];
      MultLoop_acc_1261_itm_1 <= nl_MultLoop_acc_1261_itm_1[21:0];
      MultLoop_acc_1260_itm_1 <= nl_MultLoop_acc_1260_itm_1[21:0];
      MultLoop_acc_1259_itm_1 <= nl_MultLoop_acc_1259_itm_1[21:0];
      MultLoop_acc_1258_itm_1 <= nl_MultLoop_acc_1258_itm_1[21:0];
      MultLoop_acc_1257_itm_1 <= nl_MultLoop_acc_1257_itm_1[21:0];
      MultLoop_acc_1256_itm_1 <= nl_MultLoop_acc_1256_itm_1[21:0];
      MultLoop_acc_1255_itm_1 <= nl_MultLoop_acc_1255_itm_1[21:0];
      MultLoop_acc_1254_itm_1 <= nl_MultLoop_acc_1254_itm_1[21:0];
      MultLoop_acc_1253_itm_1 <= nl_MultLoop_acc_1253_itm_1[21:0];
      MultLoop_acc_1252_itm_1 <= nl_MultLoop_acc_1252_itm_1[21:0];
      MultLoop_acc_1251_itm_1 <= nl_MultLoop_acc_1251_itm_1[21:0];
      MultLoop_acc_1250_itm_1 <= nl_MultLoop_acc_1250_itm_1[21:0];
      MultLoop_acc_1138_itm_1 <= nl_MultLoop_acc_1138_itm_1[21:0];
      MultLoop_acc_1137_itm_1 <= nl_MultLoop_acc_1137_itm_1[21:0];
      MultLoop_acc_1136_itm_1 <= nl_MultLoop_acc_1136_itm_1[21:0];
      MultLoop_acc_1135_itm_1 <= nl_MultLoop_acc_1135_itm_1[21:0];
      MultLoop_acc_1134_itm_1 <= nl_MultLoop_acc_1134_itm_1[21:0];
      MultLoop_acc_1133_itm_1 <= nl_MultLoop_acc_1133_itm_1[21:0];
      MultLoop_acc_1132_itm_1 <= nl_MultLoop_acc_1132_itm_1[21:0];
      MultLoop_acc_1131_itm_1 <= nl_MultLoop_acc_1131_itm_1[21:0];
      MultLoop_acc_1130_itm_1 <= nl_MultLoop_acc_1130_itm_1[21:0];
      MultLoop_acc_1129_itm_1 <= nl_MultLoop_acc_1129_itm_1[21:0];
      MultLoop_acc_1128_itm_1 <= nl_MultLoop_acc_1128_itm_1[21:0];
      MultLoop_acc_1127_itm_1 <= nl_MultLoop_acc_1127_itm_1[21:0];
      MultLoop_acc_1126_itm_1 <= nl_MultLoop_acc_1126_itm_1[21:0];
      MultLoop_acc_1125_itm_1 <= nl_MultLoop_acc_1125_itm_1[21:0];
      MultLoop_acc_1124_itm_1 <= nl_MultLoop_acc_1124_itm_1[21:0];
      MultLoop_acc_1123_itm_1 <= nl_MultLoop_acc_1123_itm_1[21:0];
      MultLoop_acc_1011_itm_1 <= nl_MultLoop_acc_1011_itm_1[21:0];
      MultLoop_acc_1010_itm_1 <= nl_MultLoop_acc_1010_itm_1[21:0];
      MultLoop_acc_1009_itm_1 <= nl_MultLoop_acc_1009_itm_1[21:0];
      MultLoop_acc_1008_itm_1 <= nl_MultLoop_acc_1008_itm_1[21:0];
      MultLoop_acc_1007_itm_1 <= nl_MultLoop_acc_1007_itm_1[21:0];
      MultLoop_acc_1006_itm_1 <= nl_MultLoop_acc_1006_itm_1[21:0];
      MultLoop_acc_1005_itm_1 <= nl_MultLoop_acc_1005_itm_1[21:0];
      MultLoop_acc_1004_itm_1 <= nl_MultLoop_acc_1004_itm_1[21:0];
      MultLoop_acc_1003_itm_1 <= nl_MultLoop_acc_1003_itm_1[21:0];
      MultLoop_acc_1002_itm_1 <= nl_MultLoop_acc_1002_itm_1[21:0];
      MultLoop_acc_1001_itm_1 <= nl_MultLoop_acc_1001_itm_1[21:0];
      MultLoop_acc_1000_itm_1 <= nl_MultLoop_acc_1000_itm_1[21:0];
      MultLoop_acc_999_itm_1 <= nl_MultLoop_acc_999_itm_1[21:0];
      MultLoop_acc_998_itm_1 <= nl_MultLoop_acc_998_itm_1[21:0];
      MultLoop_acc_997_itm_1 <= nl_MultLoop_acc_997_itm_1[21:0];
      MultLoop_acc_996_itm_1 <= nl_MultLoop_acc_996_itm_1[21:0];
      MultLoop_acc_884_itm_1 <= nl_MultLoop_acc_884_itm_1[21:0];
      MultLoop_acc_883_itm_1 <= nl_MultLoop_acc_883_itm_1[21:0];
      MultLoop_acc_882_itm_1 <= nl_MultLoop_acc_882_itm_1[21:0];
      MultLoop_acc_881_itm_1 <= nl_MultLoop_acc_881_itm_1[21:0];
      MultLoop_acc_880_itm_1 <= nl_MultLoop_acc_880_itm_1[21:0];
      MultLoop_acc_879_itm_1 <= nl_MultLoop_acc_879_itm_1[21:0];
      MultLoop_acc_878_itm_1 <= nl_MultLoop_acc_878_itm_1[21:0];
      MultLoop_acc_877_itm_1 <= nl_MultLoop_acc_877_itm_1[21:0];
      MultLoop_acc_876_itm_1 <= nl_MultLoop_acc_876_itm_1[21:0];
      MultLoop_acc_875_itm_1 <= nl_MultLoop_acc_875_itm_1[21:0];
      MultLoop_acc_874_itm_1 <= nl_MultLoop_acc_874_itm_1[21:0];
      MultLoop_acc_873_itm_1 <= nl_MultLoop_acc_873_itm_1[21:0];
      MultLoop_acc_872_itm_1 <= nl_MultLoop_acc_872_itm_1[21:0];
      MultLoop_acc_871_itm_1 <= nl_MultLoop_acc_871_itm_1[21:0];
      MultLoop_acc_870_itm_1 <= nl_MultLoop_acc_870_itm_1[21:0];
      MultLoop_acc_869_itm_1 <= nl_MultLoop_acc_869_itm_1[21:0];
      MultLoop_acc_757_itm_1 <= nl_MultLoop_acc_757_itm_1[21:0];
      MultLoop_acc_756_itm_1 <= nl_MultLoop_acc_756_itm_1[21:0];
      MultLoop_acc_755_itm_1 <= nl_MultLoop_acc_755_itm_1[21:0];
      MultLoop_acc_754_itm_1 <= nl_MultLoop_acc_754_itm_1[21:0];
      MultLoop_acc_753_itm_1 <= nl_MultLoop_acc_753_itm_1[21:0];
      MultLoop_acc_752_itm_1 <= nl_MultLoop_acc_752_itm_1[21:0];
      MultLoop_acc_751_itm_1 <= nl_MultLoop_acc_751_itm_1[21:0];
      MultLoop_acc_750_itm_1 <= nl_MultLoop_acc_750_itm_1[21:0];
      MultLoop_acc_749_itm_1 <= nl_MultLoop_acc_749_itm_1[21:0];
      MultLoop_acc_748_itm_1 <= nl_MultLoop_acc_748_itm_1[21:0];
      MultLoop_acc_747_itm_1 <= nl_MultLoop_acc_747_itm_1[21:0];
      MultLoop_acc_746_itm_1 <= nl_MultLoop_acc_746_itm_1[21:0];
      MultLoop_acc_745_itm_1 <= nl_MultLoop_acc_745_itm_1[21:0];
      MultLoop_acc_744_itm_1 <= nl_MultLoop_acc_744_itm_1[21:0];
      MultLoop_acc_743_itm_1 <= nl_MultLoop_acc_743_itm_1[21:0];
      MultLoop_acc_742_itm_1 <= nl_MultLoop_acc_742_itm_1[21:0];
      MultLoop_acc_630_itm_1 <= nl_MultLoop_acc_630_itm_1[21:0];
      MultLoop_acc_629_itm_1 <= nl_MultLoop_acc_629_itm_1[21:0];
      MultLoop_acc_628_itm_1 <= nl_MultLoop_acc_628_itm_1[21:0];
      MultLoop_acc_627_itm_1 <= nl_MultLoop_acc_627_itm_1[21:0];
      MultLoop_acc_626_itm_1 <= nl_MultLoop_acc_626_itm_1[21:0];
      MultLoop_acc_625_itm_1 <= nl_MultLoop_acc_625_itm_1[21:0];
      MultLoop_acc_624_itm_1 <= nl_MultLoop_acc_624_itm_1[21:0];
      MultLoop_acc_623_itm_1 <= nl_MultLoop_acc_623_itm_1[21:0];
      MultLoop_acc_622_itm_1 <= nl_MultLoop_acc_622_itm_1[21:0];
      MultLoop_acc_621_itm_1 <= nl_MultLoop_acc_621_itm_1[21:0];
      MultLoop_acc_620_itm_1 <= nl_MultLoop_acc_620_itm_1[21:0];
      MultLoop_acc_619_itm_1 <= nl_MultLoop_acc_619_itm_1[21:0];
      MultLoop_acc_618_itm_1 <= nl_MultLoop_acc_618_itm_1[21:0];
      MultLoop_acc_617_itm_1 <= nl_MultLoop_acc_617_itm_1[21:0];
      MultLoop_acc_616_itm_1 <= nl_MultLoop_acc_616_itm_1[21:0];
      MultLoop_acc_615_itm_1 <= nl_MultLoop_acc_615_itm_1[21:0];
      MultLoop_acc_503_itm_1 <= nl_MultLoop_acc_503_itm_1[21:0];
      MultLoop_acc_502_itm_1 <= nl_MultLoop_acc_502_itm_1[21:0];
      MultLoop_acc_501_itm_1 <= nl_MultLoop_acc_501_itm_1[21:0];
      MultLoop_acc_500_itm_1 <= nl_MultLoop_acc_500_itm_1[21:0];
      MultLoop_acc_499_itm_1 <= nl_MultLoop_acc_499_itm_1[21:0];
      MultLoop_acc_498_itm_1 <= nl_MultLoop_acc_498_itm_1[21:0];
      MultLoop_acc_497_itm_1 <= nl_MultLoop_acc_497_itm_1[21:0];
      MultLoop_acc_496_itm_1 <= nl_MultLoop_acc_496_itm_1[21:0];
      MultLoop_acc_495_itm_1 <= nl_MultLoop_acc_495_itm_1[21:0];
      MultLoop_acc_494_itm_1 <= nl_MultLoop_acc_494_itm_1[21:0];
      MultLoop_acc_493_itm_1 <= nl_MultLoop_acc_493_itm_1[21:0];
      MultLoop_acc_492_itm_1 <= nl_MultLoop_acc_492_itm_1[21:0];
      MultLoop_acc_491_itm_1 <= nl_MultLoop_acc_491_itm_1[21:0];
      MultLoop_acc_490_itm_1 <= nl_MultLoop_acc_490_itm_1[21:0];
      MultLoop_acc_489_itm_1 <= nl_MultLoop_acc_489_itm_1[21:0];
      MultLoop_acc_488_itm_1 <= nl_MultLoop_acc_488_itm_1[21:0];
      MultLoop_acc_376_itm_1 <= nl_MultLoop_acc_376_itm_1[21:0];
      MultLoop_acc_375_itm_1 <= nl_MultLoop_acc_375_itm_1[21:0];
      MultLoop_acc_374_itm_1 <= nl_MultLoop_acc_374_itm_1[21:0];
      MultLoop_acc_373_itm_1 <= nl_MultLoop_acc_373_itm_1[21:0];
      MultLoop_acc_372_itm_1 <= nl_MultLoop_acc_372_itm_1[21:0];
      MultLoop_acc_371_itm_1 <= nl_MultLoop_acc_371_itm_1[21:0];
      MultLoop_acc_370_itm_1 <= nl_MultLoop_acc_370_itm_1[21:0];
      MultLoop_acc_369_itm_1 <= nl_MultLoop_acc_369_itm_1[21:0];
      MultLoop_acc_368_itm_1 <= nl_MultLoop_acc_368_itm_1[21:0];
      MultLoop_acc_367_itm_1 <= nl_MultLoop_acc_367_itm_1[21:0];
      MultLoop_acc_366_itm_1 <= nl_MultLoop_acc_366_itm_1[21:0];
      MultLoop_acc_365_itm_1 <= nl_MultLoop_acc_365_itm_1[21:0];
      MultLoop_acc_364_itm_1 <= nl_MultLoop_acc_364_itm_1[21:0];
      MultLoop_acc_363_itm_1 <= nl_MultLoop_acc_363_itm_1[21:0];
      MultLoop_acc_362_itm_1 <= nl_MultLoop_acc_362_itm_1[21:0];
      MultLoop_acc_361_itm_1 <= nl_MultLoop_acc_361_itm_1[21:0];
      MultLoop_acc_249_itm_1 <= nl_MultLoop_acc_249_itm_1[21:0];
      MultLoop_acc_248_itm_1 <= nl_MultLoop_acc_248_itm_1[21:0];
      MultLoop_acc_247_itm_1 <= nl_MultLoop_acc_247_itm_1[21:0];
      MultLoop_acc_246_itm_1 <= nl_MultLoop_acc_246_itm_1[21:0];
      MultLoop_acc_245_itm_1 <= nl_MultLoop_acc_245_itm_1[21:0];
      MultLoop_acc_244_itm_1 <= nl_MultLoop_acc_244_itm_1[21:0];
      MultLoop_acc_243_itm_1 <= nl_MultLoop_acc_243_itm_1[21:0];
      MultLoop_acc_242_itm_1 <= nl_MultLoop_acc_242_itm_1[21:0];
      MultLoop_acc_241_itm_1 <= nl_MultLoop_acc_241_itm_1[21:0];
      MultLoop_acc_240_itm_1 <= nl_MultLoop_acc_240_itm_1[21:0];
      MultLoop_acc_239_itm_1 <= nl_MultLoop_acc_239_itm_1[21:0];
      MultLoop_acc_238_itm_1 <= nl_MultLoop_acc_238_itm_1[21:0];
      MultLoop_acc_237_itm_1 <= nl_MultLoop_acc_237_itm_1[21:0];
      MultLoop_acc_236_itm_1 <= nl_MultLoop_acc_236_itm_1[21:0];
      MultLoop_acc_235_itm_1 <= nl_MultLoop_acc_235_itm_1[21:0];
      MultLoop_acc_234_itm_1 <= nl_MultLoop_acc_234_itm_1[21:0];
      MultLoop_acc_130_itm_1 <= nl_MultLoop_acc_130_itm_1[21:0];
      MultLoop_acc_121_itm_1 <= nl_MultLoop_acc_121_itm_1[21:0];
      MultLoop_acc_120_itm_1 <= nl_MultLoop_acc_120_itm_1[21:0];
      MultLoop_acc_119_itm_1 <= nl_MultLoop_acc_119_itm_1[21:0];
      MultLoop_acc_118_itm_1 <= nl_MultLoop_acc_118_itm_1[21:0];
      MultLoop_acc_117_itm_1 <= nl_MultLoop_acc_117_itm_1[21:0];
      MultLoop_acc_116_itm_1 <= nl_MultLoop_acc_116_itm_1[21:0];
      MultLoop_acc_115_itm_1 <= nl_MultLoop_acc_115_itm_1[21:0];
      MultLoop_acc_114_itm_1 <= nl_MultLoop_acc_114_itm_1[21:0];
      MultLoop_acc_113_itm_1 <= nl_MultLoop_acc_113_itm_1[21:0];
      MultLoop_acc_112_itm_1 <= nl_MultLoop_acc_112_itm_1[21:0];
      MultLoop_acc_111_itm_1 <= nl_MultLoop_acc_111_itm_1[21:0];
      MultLoop_acc_110_itm_1 <= nl_MultLoop_acc_110_itm_1[21:0];
      MultLoop_acc_109_itm_1 <= nl_MultLoop_acc_109_itm_1[21:0];
      MultLoop_acc_108_itm_1 <= nl_MultLoop_acc_108_itm_1[21:0];
      MultLoop_acc_107_itm_1 <= nl_MultLoop_acc_107_itm_1[21:0];
      main_stage_0_2 <= fsm_output[1];
    end
  end
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(MultLoop_1280_MultLoop_acc_3_ncse_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(layer4_out_0_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_MultLoop_acc_1289_nl = (MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[7:0]);
  assign MultLoop_acc_1289_nl = nl_MultLoop_acc_1289_nl[10:0];
  assign nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[7:0]));
  assign MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1217_nl = ({(MultLoop_acc_1289_nl) , (MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1217_nl = nl_MultLoop_acc_1217_nl[21:0];
  assign nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[15:8]));
  assign MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[23:16]));
  assign MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1216_nl = (readslicef_29_22_7((MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1216_nl = nl_MultLoop_acc_1216_nl[21:0];
  assign nl_MultLoop_acc_1249_nl = (MultLoop_acc_1217_nl) + (MultLoop_acc_1216_nl);
  assign MultLoop_acc_1249_nl = nl_MultLoop_acc_1249_nl[21:0];
  assign nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[31:24]));
  assign MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[39:32]));
  assign MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1215_nl = (readslicef_29_22_7((MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1215_nl = nl_MultLoop_acc_1215_nl[21:0];
  assign nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[47:40]));
  assign MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[55:48]));
  assign MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1214_nl = (readslicef_29_22_7((MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1214_nl = nl_MultLoop_acc_1214_nl[21:0];
  assign nl_MultLoop_acc_1248_nl = (MultLoop_acc_1215_nl) + (MultLoop_acc_1214_nl);
  assign MultLoop_acc_1248_nl = nl_MultLoop_acc_1248_nl[21:0];
  assign nl_MultLoop_acc_1265_itm_1  = (MultLoop_acc_1249_nl) + (MultLoop_acc_1248_nl);
  assign nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[63:56]));
  assign MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[71:64]));
  assign MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1213_nl = (readslicef_29_22_7((MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1213_nl = nl_MultLoop_acc_1213_nl[21:0];
  assign nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[79:72]));
  assign MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[87:80]));
  assign MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1212_nl = (readslicef_29_22_7((MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1212_nl = nl_MultLoop_acc_1212_nl[21:0];
  assign nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[95:88]));
  assign MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[103:96]));
  assign MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1211_nl = (readslicef_29_22_7((MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1211_nl = nl_MultLoop_acc_1211_nl[21:0];
  assign nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[111:104]));
  assign MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[119:112]));
  assign MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1210_nl = (readslicef_29_22_7((MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1210_nl = nl_MultLoop_acc_1210_nl[21:0];
  assign nl_MultLoop_acc_1264_itm_1  = (MultLoop_acc_1213_nl) + (MultLoop_acc_1212_nl)
      + (MultLoop_acc_1211_nl) + (MultLoop_acc_1210_nl);
  assign nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[127:120]));
  assign MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[135:128]));
  assign MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1209_nl = (readslicef_29_22_7((MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1209_nl = nl_MultLoop_acc_1209_nl[21:0];
  assign nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[143:136]));
  assign MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[151:144]));
  assign MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1208_nl = (readslicef_29_22_7((MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1208_nl = nl_MultLoop_acc_1208_nl[21:0];
  assign nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[159:152]));
  assign MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[167:160]));
  assign MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1207_nl = (readslicef_29_22_7((MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1207_nl = nl_MultLoop_acc_1207_nl[21:0];
  assign nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[175:168]));
  assign MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[183:176]));
  assign MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1206_nl = (readslicef_29_22_7((MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1206_nl = nl_MultLoop_acc_1206_nl[21:0];
  assign nl_MultLoop_acc_1263_itm_1  = (MultLoop_acc_1209_nl) + (MultLoop_acc_1208_nl)
      + (MultLoop_acc_1207_nl) + (MultLoop_acc_1206_nl);
  assign nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[191:184]));
  assign MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[199:192]));
  assign MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1205_nl = (readslicef_29_22_7((MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1205_nl = nl_MultLoop_acc_1205_nl[21:0];
  assign nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[207:200]));
  assign MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[215:208]));
  assign MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1204_nl = (readslicef_29_22_7((MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1204_nl = nl_MultLoop_acc_1204_nl[21:0];
  assign nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[223:216]));
  assign MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[231:224]));
  assign MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1203_nl = (readslicef_29_22_7((MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1203_nl = nl_MultLoop_acc_1203_nl[21:0];
  assign nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[239:232]));
  assign MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[247:240]));
  assign MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1202_nl = (readslicef_29_22_7((MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1202_nl = nl_MultLoop_acc_1202_nl[21:0];
  assign nl_MultLoop_acc_1262_itm_1  = (MultLoop_acc_1205_nl) + (MultLoop_acc_1204_nl)
      + (MultLoop_acc_1203_nl) + (MultLoop_acc_1202_nl);
  assign nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[255:248]));
  assign MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[263:256]));
  assign MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1201_nl = (readslicef_29_22_7((MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1201_nl = nl_MultLoop_acc_1201_nl[21:0];
  assign nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[271:264]));
  assign MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[279:272]));
  assign MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1200_nl = (readslicef_29_22_7((MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1200_nl = nl_MultLoop_acc_1200_nl[21:0];
  assign nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[287:280]));
  assign MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[295:288]));
  assign MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1199_nl = (readslicef_29_22_7((MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1199_nl = nl_MultLoop_acc_1199_nl[21:0];
  assign nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[303:296]));
  assign MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[311:304]));
  assign MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1198_nl = (readslicef_29_22_7((MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1198_nl = nl_MultLoop_acc_1198_nl[21:0];
  assign nl_MultLoop_acc_1261_itm_1  = (MultLoop_acc_1201_nl) + (MultLoop_acc_1200_nl)
      + (MultLoop_acc_1199_nl) + (MultLoop_acc_1198_nl);
  assign nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[319:312]));
  assign MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[327:320]));
  assign MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1197_nl = (readslicef_29_22_7((MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1197_nl = nl_MultLoop_acc_1197_nl[21:0];
  assign nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[335:328]));
  assign MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[343:336]));
  assign MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1196_nl = (readslicef_29_22_7((MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1196_nl = nl_MultLoop_acc_1196_nl[21:0];
  assign nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[351:344]));
  assign MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[359:352]));
  assign MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1195_nl = (readslicef_29_22_7((MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1195_nl = nl_MultLoop_acc_1195_nl[21:0];
  assign nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[367:360]));
  assign MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[375:368]));
  assign MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1194_nl = (readslicef_29_22_7((MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1194_nl = nl_MultLoop_acc_1194_nl[21:0];
  assign nl_MultLoop_acc_1260_itm_1  = (MultLoop_acc_1197_nl) + (MultLoop_acc_1196_nl)
      + (MultLoop_acc_1195_nl) + (MultLoop_acc_1194_nl);
  assign nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[383:376]));
  assign MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[391:384]));
  assign MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1193_nl = (readslicef_29_22_7((MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1193_nl = nl_MultLoop_acc_1193_nl[21:0];
  assign nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[399:392]));
  assign MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[407:400]));
  assign MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1192_nl = (readslicef_29_22_7((MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1192_nl = nl_MultLoop_acc_1192_nl[21:0];
  assign nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[415:408]));
  assign MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[423:416]));
  assign MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1191_nl = (readslicef_29_22_7((MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1191_nl = nl_MultLoop_acc_1191_nl[21:0];
  assign nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[431:424]));
  assign MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[439:432]));
  assign MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1190_nl = (readslicef_29_22_7((MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1190_nl = nl_MultLoop_acc_1190_nl[21:0];
  assign nl_MultLoop_acc_1259_itm_1  = (MultLoop_acc_1193_nl) + (MultLoop_acc_1192_nl)
      + (MultLoop_acc_1191_nl) + (MultLoop_acc_1190_nl);
  assign nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[447:440]));
  assign MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[455:448]));
  assign MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1189_nl = (readslicef_29_22_7((MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1189_nl = nl_MultLoop_acc_1189_nl[21:0];
  assign nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[463:456]));
  assign MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[471:464]));
  assign MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1188_nl = (readslicef_29_22_7((MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1188_nl = nl_MultLoop_acc_1188_nl[21:0];
  assign nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[479:472]));
  assign MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[487:480]));
  assign MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1187_nl = (readslicef_29_22_7((MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1187_nl = nl_MultLoop_acc_1187_nl[21:0];
  assign nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[495:488]));
  assign MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[503:496]));
  assign MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1186_nl = (readslicef_29_22_7((MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1186_nl = nl_MultLoop_acc_1186_nl[21:0];
  assign nl_MultLoop_acc_1258_itm_1  = (MultLoop_acc_1189_nl) + (MultLoop_acc_1188_nl)
      + (MultLoop_acc_1187_nl) + (MultLoop_acc_1186_nl);
  assign nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[511:504]));
  assign MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[519:512]));
  assign MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1185_nl = (readslicef_29_22_7((MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1185_nl = nl_MultLoop_acc_1185_nl[21:0];
  assign nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[527:520]));
  assign MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[535:528]));
  assign MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1184_nl = (readslicef_29_22_7((MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1184_nl = nl_MultLoop_acc_1184_nl[21:0];
  assign nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[543:536]));
  assign MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[551:544]));
  assign MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1183_nl = (readslicef_29_22_7((MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1183_nl = nl_MultLoop_acc_1183_nl[21:0];
  assign nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[559:552]));
  assign MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[567:560]));
  assign MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1182_nl = (readslicef_29_22_7((MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1182_nl = nl_MultLoop_acc_1182_nl[21:0];
  assign nl_MultLoop_acc_1257_itm_1  = (MultLoop_acc_1185_nl) + (MultLoop_acc_1184_nl)
      + (MultLoop_acc_1183_nl) + (MultLoop_acc_1182_nl);
  assign nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[575:568]));
  assign MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[583:576]));
  assign MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1181_nl = (readslicef_29_22_7((MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1181_nl = nl_MultLoop_acc_1181_nl[21:0];
  assign nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[591:584]));
  assign MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[599:592]));
  assign MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1180_nl = (readslicef_29_22_7((MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1180_nl = nl_MultLoop_acc_1180_nl[21:0];
  assign nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[607:600]));
  assign MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[615:608]));
  assign MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1179_nl = (readslicef_29_22_7((MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1179_nl = nl_MultLoop_acc_1179_nl[21:0];
  assign nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[623:616]));
  assign MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[631:624]));
  assign MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1178_nl = (readslicef_29_22_7((MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1178_nl = nl_MultLoop_acc_1178_nl[21:0];
  assign nl_MultLoop_acc_1256_itm_1  = (MultLoop_acc_1181_nl) + (MultLoop_acc_1180_nl)
      + (MultLoop_acc_1179_nl) + (MultLoop_acc_1178_nl);
  assign nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[639:632]));
  assign MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[647:640]));
  assign MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1177_nl = (readslicef_29_22_7((MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1177_nl = nl_MultLoop_acc_1177_nl[21:0];
  assign nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[655:648]));
  assign MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[663:656]));
  assign MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1176_nl = (readslicef_29_22_7((MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1176_nl = nl_MultLoop_acc_1176_nl[21:0];
  assign nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[671:664]));
  assign MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[679:672]));
  assign MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1175_nl = (readslicef_29_22_7((MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1175_nl = nl_MultLoop_acc_1175_nl[21:0];
  assign nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[687:680]));
  assign MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[695:688]));
  assign MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1174_nl = (readslicef_29_22_7((MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1174_nl = nl_MultLoop_acc_1174_nl[21:0];
  assign nl_MultLoop_acc_1255_itm_1  = (MultLoop_acc_1177_nl) + (MultLoop_acc_1176_nl)
      + (MultLoop_acc_1175_nl) + (MultLoop_acc_1174_nl);
  assign nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[703:696]));
  assign MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[711:704]));
  assign MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1173_nl = (readslicef_29_22_7((MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1173_nl = nl_MultLoop_acc_1173_nl[21:0];
  assign nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[719:712]));
  assign MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[727:720]));
  assign MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1172_nl = (readslicef_29_22_7((MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1172_nl = nl_MultLoop_acc_1172_nl[21:0];
  assign nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[735:728]));
  assign MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[743:736]));
  assign MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1171_nl = (readslicef_29_22_7((MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1171_nl = nl_MultLoop_acc_1171_nl[21:0];
  assign nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[751:744]));
  assign MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[759:752]));
  assign MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1170_nl = (readslicef_29_22_7((MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1170_nl = nl_MultLoop_acc_1170_nl[21:0];
  assign nl_MultLoop_acc_1254_itm_1  = (MultLoop_acc_1173_nl) + (MultLoop_acc_1172_nl)
      + (MultLoop_acc_1171_nl) + (MultLoop_acc_1170_nl);
  assign nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[767:760]));
  assign MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[775:768]));
  assign MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1169_nl = (readslicef_29_22_7((MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1169_nl = nl_MultLoop_acc_1169_nl[21:0];
  assign nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[783:776]));
  assign MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[791:784]));
  assign MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1168_nl = (readslicef_29_22_7((MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1168_nl = nl_MultLoop_acc_1168_nl[21:0];
  assign nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[799:792]));
  assign MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[807:800]));
  assign MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1167_nl = (readslicef_29_22_7((MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1167_nl = nl_MultLoop_acc_1167_nl[21:0];
  assign nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[815:808]));
  assign MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[823:816]));
  assign MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1166_nl = (readslicef_29_22_7((MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1166_nl = nl_MultLoop_acc_1166_nl[21:0];
  assign nl_MultLoop_acc_1253_itm_1  = (MultLoop_acc_1169_nl) + (MultLoop_acc_1168_nl)
      + (MultLoop_acc_1167_nl) + (MultLoop_acc_1166_nl);
  assign nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[831:824]));
  assign MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[839:832]));
  assign MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1165_nl = (readslicef_29_22_7((MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1165_nl = nl_MultLoop_acc_1165_nl[21:0];
  assign nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[847:840]));
  assign MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[855:848]));
  assign MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1164_nl = (readslicef_29_22_7((MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1164_nl = nl_MultLoop_acc_1164_nl[21:0];
  assign nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[863:856]));
  assign MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[871:864]));
  assign MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1163_nl = (readslicef_29_22_7((MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1163_nl = nl_MultLoop_acc_1163_nl[21:0];
  assign nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[879:872]));
  assign MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[887:880]));
  assign MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1162_nl = (readslicef_29_22_7((MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1162_nl = nl_MultLoop_acc_1162_nl[21:0];
  assign nl_MultLoop_acc_1252_itm_1  = (MultLoop_acc_1165_nl) + (MultLoop_acc_1164_nl)
      + (MultLoop_acc_1163_nl) + (MultLoop_acc_1162_nl);
  assign nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[895:888]));
  assign MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[903:896]));
  assign MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1161_nl = (readslicef_29_22_7((MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1161_nl = nl_MultLoop_acc_1161_nl[21:0];
  assign nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[911:904]));
  assign MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[919:912]));
  assign MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1160_nl = (readslicef_29_22_7((MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1160_nl = nl_MultLoop_acc_1160_nl[21:0];
  assign nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[927:920]));
  assign MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[935:928]));
  assign MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1159_nl = (readslicef_29_22_7((MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1159_nl = nl_MultLoop_acc_1159_nl[21:0];
  assign nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[943:936]));
  assign MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[951:944]));
  assign MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1158_nl = (readslicef_29_22_7((MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1158_nl = nl_MultLoop_acc_1158_nl[21:0];
  assign nl_MultLoop_acc_1251_itm_1  = (MultLoop_acc_1161_nl) + (MultLoop_acc_1160_nl)
      + (MultLoop_acc_1159_nl) + (MultLoop_acc_1158_nl);
  assign nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[959:952]));
  assign MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[967:960]));
  assign MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1157_nl = (readslicef_29_22_7((MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1157_nl = nl_MultLoop_acc_1157_nl[21:0];
  assign nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[975:968]));
  assign MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[983:976]));
  assign MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1156_nl = (readslicef_29_22_7((MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1156_nl = nl_MultLoop_acc_1156_nl[21:0];
  assign nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[991:984]));
  assign MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[999:992]));
  assign MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1155_nl = (readslicef_29_22_7((MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1155_nl = nl_MultLoop_acc_1155_nl[21:0];
  assign nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1007:1000]));
  assign MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1015:1008]));
  assign MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1154_nl = (readslicef_29_22_7((MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1154_nl = nl_MultLoop_acc_1154_nl[21:0];
  assign nl_MultLoop_acc_1250_itm_1  = (MultLoop_acc_1157_nl) + (MultLoop_acc_1156_nl)
      + (MultLoop_acc_1155_nl) + (MultLoop_acc_1154_nl);
  assign nl_MultLoop_acc_1288_nl = (MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[79:72]);
  assign MultLoop_acc_1288_nl = nl_MultLoop_acc_1288_nl[10:0];
  assign nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[9223:9216]));
  assign MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1090_nl = ({(MultLoop_acc_1288_nl) , (MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1090_nl = nl_MultLoop_acc_1090_nl[21:0];
  assign nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9231:9224]));
  assign MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9239:9232]));
  assign MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1089_nl = (readslicef_29_22_7((MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1089_nl = nl_MultLoop_acc_1089_nl[21:0];
  assign nl_MultLoop_acc_1122_nl = (MultLoop_acc_1090_nl) + (MultLoop_acc_1089_nl);
  assign MultLoop_acc_1122_nl = nl_MultLoop_acc_1122_nl[21:0];
  assign nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9247:9240]));
  assign MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9255:9248]));
  assign MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1088_nl = (readslicef_29_22_7((MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1088_nl = nl_MultLoop_acc_1088_nl[21:0];
  assign nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9263:9256]));
  assign MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9271:9264]));
  assign MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1087_nl = (readslicef_29_22_7((MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1087_nl = nl_MultLoop_acc_1087_nl[21:0];
  assign nl_MultLoop_acc_1121_nl = (MultLoop_acc_1088_nl) + (MultLoop_acc_1087_nl);
  assign MultLoop_acc_1121_nl = nl_MultLoop_acc_1121_nl[21:0];
  assign nl_MultLoop_acc_1138_itm_1  = (MultLoop_acc_1122_nl) + (MultLoop_acc_1121_nl);
  assign nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9279:9272]));
  assign MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9287:9280]));
  assign MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1086_nl = (readslicef_29_22_7((MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1086_nl = nl_MultLoop_acc_1086_nl[21:0];
  assign nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9295:9288]));
  assign MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9303:9296]));
  assign MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1085_nl = (readslicef_29_22_7((MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1085_nl = nl_MultLoop_acc_1085_nl[21:0];
  assign nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9311:9304]));
  assign MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9319:9312]));
  assign MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1084_nl = (readslicef_29_22_7((MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1084_nl = nl_MultLoop_acc_1084_nl[21:0];
  assign nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9327:9320]));
  assign MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9335:9328]));
  assign MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1083_nl = (readslicef_29_22_7((MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1083_nl = nl_MultLoop_acc_1083_nl[21:0];
  assign nl_MultLoop_acc_1137_itm_1  = (MultLoop_acc_1086_nl) + (MultLoop_acc_1085_nl)
      + (MultLoop_acc_1084_nl) + (MultLoop_acc_1083_nl);
  assign nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9343:9336]));
  assign MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9351:9344]));
  assign MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1082_nl = (readslicef_29_22_7((MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1082_nl = nl_MultLoop_acc_1082_nl[21:0];
  assign nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9359:9352]));
  assign MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9367:9360]));
  assign MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1081_nl = (readslicef_29_22_7((MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1081_nl = nl_MultLoop_acc_1081_nl[21:0];
  assign nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9375:9368]));
  assign MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9383:9376]));
  assign MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1080_nl = (readslicef_29_22_7((MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1080_nl = nl_MultLoop_acc_1080_nl[21:0];
  assign nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9391:9384]));
  assign MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9399:9392]));
  assign MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1079_nl = (readslicef_29_22_7((MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1079_nl = nl_MultLoop_acc_1079_nl[21:0];
  assign nl_MultLoop_acc_1136_itm_1  = (MultLoop_acc_1082_nl) + (MultLoop_acc_1081_nl)
      + (MultLoop_acc_1080_nl) + (MultLoop_acc_1079_nl);
  assign nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9407:9400]));
  assign MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9415:9408]));
  assign MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1078_nl = (readslicef_29_22_7((MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1078_nl = nl_MultLoop_acc_1078_nl[21:0];
  assign nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9423:9416]));
  assign MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9431:9424]));
  assign MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1077_nl = (readslicef_29_22_7((MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1077_nl = nl_MultLoop_acc_1077_nl[21:0];
  assign nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9439:9432]));
  assign MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9447:9440]));
  assign MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1076_nl = (readslicef_29_22_7((MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1076_nl = nl_MultLoop_acc_1076_nl[21:0];
  assign nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9455:9448]));
  assign MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9463:9456]));
  assign MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1075_nl = (readslicef_29_22_7((MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1075_nl = nl_MultLoop_acc_1075_nl[21:0];
  assign nl_MultLoop_acc_1135_itm_1  = (MultLoop_acc_1078_nl) + (MultLoop_acc_1077_nl)
      + (MultLoop_acc_1076_nl) + (MultLoop_acc_1075_nl);
  assign nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9471:9464]));
  assign MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9479:9472]));
  assign MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1074_nl = (readslicef_29_22_7((MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1074_nl = nl_MultLoop_acc_1074_nl[21:0];
  assign nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9487:9480]));
  assign MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9495:9488]));
  assign MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1073_nl = (readslicef_29_22_7((MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1073_nl = nl_MultLoop_acc_1073_nl[21:0];
  assign nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9503:9496]));
  assign MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9511:9504]));
  assign MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1072_nl = (readslicef_29_22_7((MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1072_nl = nl_MultLoop_acc_1072_nl[21:0];
  assign nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9519:9512]));
  assign MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9527:9520]));
  assign MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1071_nl = (readslicef_29_22_7((MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1071_nl = nl_MultLoop_acc_1071_nl[21:0];
  assign nl_MultLoop_acc_1134_itm_1  = (MultLoop_acc_1074_nl) + (MultLoop_acc_1073_nl)
      + (MultLoop_acc_1072_nl) + (MultLoop_acc_1071_nl);
  assign nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9535:9528]));
  assign MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9543:9536]));
  assign MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1070_nl = (readslicef_29_22_7((MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1070_nl = nl_MultLoop_acc_1070_nl[21:0];
  assign nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9551:9544]));
  assign MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9559:9552]));
  assign MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1069_nl = (readslicef_29_22_7((MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1069_nl = nl_MultLoop_acc_1069_nl[21:0];
  assign nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9567:9560]));
  assign MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9575:9568]));
  assign MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1068_nl = (readslicef_29_22_7((MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1068_nl = nl_MultLoop_acc_1068_nl[21:0];
  assign nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9583:9576]));
  assign MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9591:9584]));
  assign MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1067_nl = (readslicef_29_22_7((MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1067_nl = nl_MultLoop_acc_1067_nl[21:0];
  assign nl_MultLoop_acc_1133_itm_1  = (MultLoop_acc_1070_nl) + (MultLoop_acc_1069_nl)
      + (MultLoop_acc_1068_nl) + (MultLoop_acc_1067_nl);
  assign nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9599:9592]));
  assign MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9607:9600]));
  assign MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1066_nl = (readslicef_29_22_7((MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1066_nl = nl_MultLoop_acc_1066_nl[21:0];
  assign nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9615:9608]));
  assign MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9623:9616]));
  assign MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1065_nl = (readslicef_29_22_7((MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1065_nl = nl_MultLoop_acc_1065_nl[21:0];
  assign nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9631:9624]));
  assign MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9639:9632]));
  assign MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1064_nl = (readslicef_29_22_7((MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1064_nl = nl_MultLoop_acc_1064_nl[21:0];
  assign nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9647:9640]));
  assign MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9655:9648]));
  assign MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1063_nl = (readslicef_29_22_7((MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1063_nl = nl_MultLoop_acc_1063_nl[21:0];
  assign nl_MultLoop_acc_1132_itm_1  = (MultLoop_acc_1066_nl) + (MultLoop_acc_1065_nl)
      + (MultLoop_acc_1064_nl) + (MultLoop_acc_1063_nl);
  assign nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9663:9656]));
  assign MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9671:9664]));
  assign MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1062_nl = (readslicef_29_22_7((MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1062_nl = nl_MultLoop_acc_1062_nl[21:0];
  assign nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9679:9672]));
  assign MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9687:9680]));
  assign MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1061_nl = (readslicef_29_22_7((MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1061_nl = nl_MultLoop_acc_1061_nl[21:0];
  assign nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9695:9688]));
  assign MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9703:9696]));
  assign MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1060_nl = (readslicef_29_22_7((MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1060_nl = nl_MultLoop_acc_1060_nl[21:0];
  assign nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9711:9704]));
  assign MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9719:9712]));
  assign MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1059_nl = (readslicef_29_22_7((MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1059_nl = nl_MultLoop_acc_1059_nl[21:0];
  assign nl_MultLoop_acc_1131_itm_1  = (MultLoop_acc_1062_nl) + (MultLoop_acc_1061_nl)
      + (MultLoop_acc_1060_nl) + (MultLoop_acc_1059_nl);
  assign nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9727:9720]));
  assign MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9735:9728]));
  assign MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1058_nl = (readslicef_29_22_7((MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1058_nl = nl_MultLoop_acc_1058_nl[21:0];
  assign nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9743:9736]));
  assign MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9751:9744]));
  assign MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1057_nl = (readslicef_29_22_7((MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1057_nl = nl_MultLoop_acc_1057_nl[21:0];
  assign nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9759:9752]));
  assign MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9767:9760]));
  assign MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1056_nl = (readslicef_29_22_7((MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1056_nl = nl_MultLoop_acc_1056_nl[21:0];
  assign nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9775:9768]));
  assign MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9783:9776]));
  assign MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1055_nl = (readslicef_29_22_7((MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1055_nl = nl_MultLoop_acc_1055_nl[21:0];
  assign nl_MultLoop_acc_1130_itm_1  = (MultLoop_acc_1058_nl) + (MultLoop_acc_1057_nl)
      + (MultLoop_acc_1056_nl) + (MultLoop_acc_1055_nl);
  assign nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9791:9784]));
  assign MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9799:9792]));
  assign MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1054_nl = (readslicef_29_22_7((MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1054_nl = nl_MultLoop_acc_1054_nl[21:0];
  assign nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9807:9800]));
  assign MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9815:9808]));
  assign MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1053_nl = (readslicef_29_22_7((MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1053_nl = nl_MultLoop_acc_1053_nl[21:0];
  assign nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9823:9816]));
  assign MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9831:9824]));
  assign MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1052_nl = (readslicef_29_22_7((MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1052_nl = nl_MultLoop_acc_1052_nl[21:0];
  assign nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9839:9832]));
  assign MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9847:9840]));
  assign MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1051_nl = (readslicef_29_22_7((MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1051_nl = nl_MultLoop_acc_1051_nl[21:0];
  assign nl_MultLoop_acc_1129_itm_1  = (MultLoop_acc_1054_nl) + (MultLoop_acc_1053_nl)
      + (MultLoop_acc_1052_nl) + (MultLoop_acc_1051_nl);
  assign nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9855:9848]));
  assign MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9863:9856]));
  assign MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1050_nl = (readslicef_29_22_7((MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1050_nl = nl_MultLoop_acc_1050_nl[21:0];
  assign nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9871:9864]));
  assign MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9879:9872]));
  assign MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1049_nl = (readslicef_29_22_7((MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1049_nl = nl_MultLoop_acc_1049_nl[21:0];
  assign nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9887:9880]));
  assign MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9895:9888]));
  assign MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1048_nl = (readslicef_29_22_7((MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1048_nl = nl_MultLoop_acc_1048_nl[21:0];
  assign nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9903:9896]));
  assign MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9911:9904]));
  assign MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1047_nl = (readslicef_29_22_7((MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1047_nl = nl_MultLoop_acc_1047_nl[21:0];
  assign nl_MultLoop_acc_1128_itm_1  = (MultLoop_acc_1050_nl) + (MultLoop_acc_1049_nl)
      + (MultLoop_acc_1048_nl) + (MultLoop_acc_1047_nl);
  assign nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9919:9912]));
  assign MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9927:9920]));
  assign MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1046_nl = (readslicef_29_22_7((MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1046_nl = nl_MultLoop_acc_1046_nl[21:0];
  assign nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9935:9928]));
  assign MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9943:9936]));
  assign MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1045_nl = (readslicef_29_22_7((MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1045_nl = nl_MultLoop_acc_1045_nl[21:0];
  assign nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9951:9944]));
  assign MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9959:9952]));
  assign MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1044_nl = (readslicef_29_22_7((MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1044_nl = nl_MultLoop_acc_1044_nl[21:0];
  assign nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9967:9960]));
  assign MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9975:9968]));
  assign MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1043_nl = (readslicef_29_22_7((MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1043_nl = nl_MultLoop_acc_1043_nl[21:0];
  assign nl_MultLoop_acc_1127_itm_1  = (MultLoop_acc_1046_nl) + (MultLoop_acc_1045_nl)
      + (MultLoop_acc_1044_nl) + (MultLoop_acc_1043_nl);
  assign nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9983:9976]));
  assign MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9991:9984]));
  assign MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1042_nl = (readslicef_29_22_7((MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1042_nl = nl_MultLoop_acc_1042_nl[21:0];
  assign nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9999:9992]));
  assign MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10007:10000]));
  assign MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1041_nl = (readslicef_29_22_7((MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1041_nl = nl_MultLoop_acc_1041_nl[21:0];
  assign nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10015:10008]));
  assign MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10023:10016]));
  assign MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1040_nl = (readslicef_29_22_7((MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1040_nl = nl_MultLoop_acc_1040_nl[21:0];
  assign nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10031:10024]));
  assign MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10039:10032]));
  assign MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1039_nl = (readslicef_29_22_7((MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1039_nl = nl_MultLoop_acc_1039_nl[21:0];
  assign nl_MultLoop_acc_1126_itm_1  = (MultLoop_acc_1042_nl) + (MultLoop_acc_1041_nl)
      + (MultLoop_acc_1040_nl) + (MultLoop_acc_1039_nl);
  assign nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10047:10040]));
  assign MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10055:10048]));
  assign MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1038_nl = (readslicef_29_22_7((MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1038_nl = nl_MultLoop_acc_1038_nl[21:0];
  assign nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10063:10056]));
  assign MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10071:10064]));
  assign MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1037_nl = (readslicef_29_22_7((MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1037_nl = nl_MultLoop_acc_1037_nl[21:0];
  assign nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10079:10072]));
  assign MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10087:10080]));
  assign MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1036_nl = (readslicef_29_22_7((MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1036_nl = nl_MultLoop_acc_1036_nl[21:0];
  assign nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10095:10088]));
  assign MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10103:10096]));
  assign MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1035_nl = (readslicef_29_22_7((MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1035_nl = nl_MultLoop_acc_1035_nl[21:0];
  assign nl_MultLoop_acc_1125_itm_1  = (MultLoop_acc_1038_nl) + (MultLoop_acc_1037_nl)
      + (MultLoop_acc_1036_nl) + (MultLoop_acc_1035_nl);
  assign nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10111:10104]));
  assign MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10119:10112]));
  assign MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1034_nl = (readslicef_29_22_7((MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1034_nl = nl_MultLoop_acc_1034_nl[21:0];
  assign nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10127:10120]));
  assign MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10135:10128]));
  assign MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1033_nl = (readslicef_29_22_7((MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1033_nl = nl_MultLoop_acc_1033_nl[21:0];
  assign nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10143:10136]));
  assign MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10151:10144]));
  assign MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1032_nl = (readslicef_29_22_7((MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1032_nl = nl_MultLoop_acc_1032_nl[21:0];
  assign nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10159:10152]));
  assign MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10167:10160]));
  assign MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1031_nl = (readslicef_29_22_7((MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1031_nl = nl_MultLoop_acc_1031_nl[21:0];
  assign nl_MultLoop_acc_1124_itm_1  = (MultLoop_acc_1034_nl) + (MultLoop_acc_1033_nl)
      + (MultLoop_acc_1032_nl) + (MultLoop_acc_1031_nl);
  assign nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10175:10168]));
  assign MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10183:10176]));
  assign MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1030_nl = (readslicef_29_22_7((MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1030_nl = nl_MultLoop_acc_1030_nl[21:0];
  assign nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10191:10184]));
  assign MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10199:10192]));
  assign MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1029_nl = (readslicef_29_22_7((MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1029_nl = nl_MultLoop_acc_1029_nl[21:0];
  assign nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10207:10200]));
  assign MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10215:10208]));
  assign MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1028_nl = (readslicef_29_22_7((MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1028_nl = nl_MultLoop_acc_1028_nl[21:0];
  assign nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10223:10216]));
  assign MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10231:10224]));
  assign MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1027_nl = (readslicef_29_22_7((MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1027_nl = nl_MultLoop_acc_1027_nl[21:0];
  assign nl_MultLoop_acc_1123_itm_1  = (MultLoop_acc_1030_nl) + (MultLoop_acc_1029_nl)
      + (MultLoop_acc_1028_nl) + (MultLoop_acc_1027_nl);
  assign nl_MultLoop_acc_1287_nl = (MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[71:64]);
  assign MultLoop_acc_1287_nl = nl_MultLoop_acc_1287_nl[10:0];
  assign nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[8199:8192]));
  assign MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_963_nl = ({(MultLoop_acc_1287_nl) , (MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_963_nl = nl_MultLoop_acc_963_nl[21:0];
  assign nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8207:8200]));
  assign MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8215:8208]));
  assign MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_962_nl = (readslicef_29_22_7((MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_962_nl = nl_MultLoop_acc_962_nl[21:0];
  assign nl_MultLoop_acc_995_nl = (MultLoop_acc_963_nl) + (MultLoop_acc_962_nl);
  assign MultLoop_acc_995_nl = nl_MultLoop_acc_995_nl[21:0];
  assign nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8223:8216]));
  assign MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8231:8224]));
  assign MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_961_nl = (readslicef_29_22_7((MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_961_nl = nl_MultLoop_acc_961_nl[21:0];
  assign nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8239:8232]));
  assign MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8247:8240]));
  assign MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_960_nl = (readslicef_29_22_7((MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_960_nl = nl_MultLoop_acc_960_nl[21:0];
  assign nl_MultLoop_acc_994_nl = (MultLoop_acc_961_nl) + (MultLoop_acc_960_nl);
  assign MultLoop_acc_994_nl = nl_MultLoop_acc_994_nl[21:0];
  assign nl_MultLoop_acc_1011_itm_1  = (MultLoop_acc_995_nl) + (MultLoop_acc_994_nl);
  assign nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8255:8248]));
  assign MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8263:8256]));
  assign MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_959_nl = (readslicef_29_22_7((MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_959_nl = nl_MultLoop_acc_959_nl[21:0];
  assign nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8271:8264]));
  assign MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8279:8272]));
  assign MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_958_nl = (readslicef_29_22_7((MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_958_nl = nl_MultLoop_acc_958_nl[21:0];
  assign nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8287:8280]));
  assign MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8295:8288]));
  assign MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_957_nl = (readslicef_29_22_7((MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_957_nl = nl_MultLoop_acc_957_nl[21:0];
  assign nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8303:8296]));
  assign MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8311:8304]));
  assign MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_956_nl = (readslicef_29_22_7((MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_956_nl = nl_MultLoop_acc_956_nl[21:0];
  assign nl_MultLoop_acc_1010_itm_1  = (MultLoop_acc_959_nl) + (MultLoop_acc_958_nl)
      + (MultLoop_acc_957_nl) + (MultLoop_acc_956_nl);
  assign nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8319:8312]));
  assign MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8327:8320]));
  assign MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_955_nl = (readslicef_29_22_7((MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_955_nl = nl_MultLoop_acc_955_nl[21:0];
  assign nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8335:8328]));
  assign MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8343:8336]));
  assign MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_954_nl = (readslicef_29_22_7((MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_954_nl = nl_MultLoop_acc_954_nl[21:0];
  assign nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8351:8344]));
  assign MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8359:8352]));
  assign MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_953_nl = (readslicef_29_22_7((MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_953_nl = nl_MultLoop_acc_953_nl[21:0];
  assign nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8367:8360]));
  assign MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8375:8368]));
  assign MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_952_nl = (readslicef_29_22_7((MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_952_nl = nl_MultLoop_acc_952_nl[21:0];
  assign nl_MultLoop_acc_1009_itm_1  = (MultLoop_acc_955_nl) + (MultLoop_acc_954_nl)
      + (MultLoop_acc_953_nl) + (MultLoop_acc_952_nl);
  assign nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8383:8376]));
  assign MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8391:8384]));
  assign MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_951_nl = (readslicef_29_22_7((MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_951_nl = nl_MultLoop_acc_951_nl[21:0];
  assign nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8399:8392]));
  assign MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8407:8400]));
  assign MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_950_nl = (readslicef_29_22_7((MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_950_nl = nl_MultLoop_acc_950_nl[21:0];
  assign nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8415:8408]));
  assign MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8423:8416]));
  assign MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_949_nl = (readslicef_29_22_7((MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_949_nl = nl_MultLoop_acc_949_nl[21:0];
  assign nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8431:8424]));
  assign MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8439:8432]));
  assign MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_948_nl = (readslicef_29_22_7((MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_948_nl = nl_MultLoop_acc_948_nl[21:0];
  assign nl_MultLoop_acc_1008_itm_1  = (MultLoop_acc_951_nl) + (MultLoop_acc_950_nl)
      + (MultLoop_acc_949_nl) + (MultLoop_acc_948_nl);
  assign nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8447:8440]));
  assign MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8455:8448]));
  assign MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_947_nl = (readslicef_29_22_7((MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_947_nl = nl_MultLoop_acc_947_nl[21:0];
  assign nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8463:8456]));
  assign MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8471:8464]));
  assign MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_946_nl = (readslicef_29_22_7((MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_946_nl = nl_MultLoop_acc_946_nl[21:0];
  assign nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8479:8472]));
  assign MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8487:8480]));
  assign MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_945_nl = (readslicef_29_22_7((MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_945_nl = nl_MultLoop_acc_945_nl[21:0];
  assign nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8495:8488]));
  assign MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8503:8496]));
  assign MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_944_nl = (readslicef_29_22_7((MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_944_nl = nl_MultLoop_acc_944_nl[21:0];
  assign nl_MultLoop_acc_1007_itm_1  = (MultLoop_acc_947_nl) + (MultLoop_acc_946_nl)
      + (MultLoop_acc_945_nl) + (MultLoop_acc_944_nl);
  assign nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8511:8504]));
  assign MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8519:8512]));
  assign MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_943_nl = (readslicef_29_22_7((MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_943_nl = nl_MultLoop_acc_943_nl[21:0];
  assign nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8527:8520]));
  assign MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8535:8528]));
  assign MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_942_nl = (readslicef_29_22_7((MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_942_nl = nl_MultLoop_acc_942_nl[21:0];
  assign nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8543:8536]));
  assign MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8551:8544]));
  assign MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_941_nl = (readslicef_29_22_7((MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_941_nl = nl_MultLoop_acc_941_nl[21:0];
  assign nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8559:8552]));
  assign MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8567:8560]));
  assign MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_940_nl = (readslicef_29_22_7((MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_940_nl = nl_MultLoop_acc_940_nl[21:0];
  assign nl_MultLoop_acc_1006_itm_1  = (MultLoop_acc_943_nl) + (MultLoop_acc_942_nl)
      + (MultLoop_acc_941_nl) + (MultLoop_acc_940_nl);
  assign nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8575:8568]));
  assign MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8583:8576]));
  assign MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_939_nl = (readslicef_29_22_7((MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_939_nl = nl_MultLoop_acc_939_nl[21:0];
  assign nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8591:8584]));
  assign MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8599:8592]));
  assign MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_938_nl = (readslicef_29_22_7((MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_938_nl = nl_MultLoop_acc_938_nl[21:0];
  assign nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8607:8600]));
  assign MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8615:8608]));
  assign MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_937_nl = (readslicef_29_22_7((MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_937_nl = nl_MultLoop_acc_937_nl[21:0];
  assign nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8623:8616]));
  assign MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8631:8624]));
  assign MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_936_nl = (readslicef_29_22_7((MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_936_nl = nl_MultLoop_acc_936_nl[21:0];
  assign nl_MultLoop_acc_1005_itm_1  = (MultLoop_acc_939_nl) + (MultLoop_acc_938_nl)
      + (MultLoop_acc_937_nl) + (MultLoop_acc_936_nl);
  assign nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8639:8632]));
  assign MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8647:8640]));
  assign MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_935_nl = (readslicef_29_22_7((MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_935_nl = nl_MultLoop_acc_935_nl[21:0];
  assign nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8655:8648]));
  assign MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8663:8656]));
  assign MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_934_nl = (readslicef_29_22_7((MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_934_nl = nl_MultLoop_acc_934_nl[21:0];
  assign nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8671:8664]));
  assign MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8679:8672]));
  assign MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_933_nl = (readslicef_29_22_7((MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_933_nl = nl_MultLoop_acc_933_nl[21:0];
  assign nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8687:8680]));
  assign MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8695:8688]));
  assign MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_932_nl = (readslicef_29_22_7((MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_932_nl = nl_MultLoop_acc_932_nl[21:0];
  assign nl_MultLoop_acc_1004_itm_1  = (MultLoop_acc_935_nl) + (MultLoop_acc_934_nl)
      + (MultLoop_acc_933_nl) + (MultLoop_acc_932_nl);
  assign nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8703:8696]));
  assign MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8711:8704]));
  assign MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_931_nl = (readslicef_29_22_7((MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_931_nl = nl_MultLoop_acc_931_nl[21:0];
  assign nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8719:8712]));
  assign MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8727:8720]));
  assign MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_930_nl = (readslicef_29_22_7((MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_930_nl = nl_MultLoop_acc_930_nl[21:0];
  assign nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8735:8728]));
  assign MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8743:8736]));
  assign MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_929_nl = (readslicef_29_22_7((MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_929_nl = nl_MultLoop_acc_929_nl[21:0];
  assign nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8751:8744]));
  assign MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8759:8752]));
  assign MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_928_nl = (readslicef_29_22_7((MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_928_nl = nl_MultLoop_acc_928_nl[21:0];
  assign nl_MultLoop_acc_1003_itm_1  = (MultLoop_acc_931_nl) + (MultLoop_acc_930_nl)
      + (MultLoop_acc_929_nl) + (MultLoop_acc_928_nl);
  assign nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8767:8760]));
  assign MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8775:8768]));
  assign MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_927_nl = (readslicef_29_22_7((MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_927_nl = nl_MultLoop_acc_927_nl[21:0];
  assign nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8783:8776]));
  assign MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8791:8784]));
  assign MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_926_nl = (readslicef_29_22_7((MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_926_nl = nl_MultLoop_acc_926_nl[21:0];
  assign nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8799:8792]));
  assign MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8807:8800]));
  assign MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_925_nl = (readslicef_29_22_7((MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_925_nl = nl_MultLoop_acc_925_nl[21:0];
  assign nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8815:8808]));
  assign MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8823:8816]));
  assign MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_924_nl = (readslicef_29_22_7((MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_924_nl = nl_MultLoop_acc_924_nl[21:0];
  assign nl_MultLoop_acc_1002_itm_1  = (MultLoop_acc_927_nl) + (MultLoop_acc_926_nl)
      + (MultLoop_acc_925_nl) + (MultLoop_acc_924_nl);
  assign nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8831:8824]));
  assign MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8839:8832]));
  assign MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_923_nl = (readslicef_29_22_7((MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_923_nl = nl_MultLoop_acc_923_nl[21:0];
  assign nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8847:8840]));
  assign MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8855:8848]));
  assign MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_922_nl = (readslicef_29_22_7((MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_922_nl = nl_MultLoop_acc_922_nl[21:0];
  assign nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8863:8856]));
  assign MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8871:8864]));
  assign MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_921_nl = (readslicef_29_22_7((MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_921_nl = nl_MultLoop_acc_921_nl[21:0];
  assign nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8879:8872]));
  assign MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8887:8880]));
  assign MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_920_nl = (readslicef_29_22_7((MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_920_nl = nl_MultLoop_acc_920_nl[21:0];
  assign nl_MultLoop_acc_1001_itm_1  = (MultLoop_acc_923_nl) + (MultLoop_acc_922_nl)
      + (MultLoop_acc_921_nl) + (MultLoop_acc_920_nl);
  assign nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8895:8888]));
  assign MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8903:8896]));
  assign MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_919_nl = (readslicef_29_22_7((MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_919_nl = nl_MultLoop_acc_919_nl[21:0];
  assign nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8911:8904]));
  assign MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8919:8912]));
  assign MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_918_nl = (readslicef_29_22_7((MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_918_nl = nl_MultLoop_acc_918_nl[21:0];
  assign nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8927:8920]));
  assign MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8935:8928]));
  assign MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_917_nl = (readslicef_29_22_7((MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_917_nl = nl_MultLoop_acc_917_nl[21:0];
  assign nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8943:8936]));
  assign MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8951:8944]));
  assign MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_916_nl = (readslicef_29_22_7((MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_916_nl = nl_MultLoop_acc_916_nl[21:0];
  assign nl_MultLoop_acc_1000_itm_1  = (MultLoop_acc_919_nl) + (MultLoop_acc_918_nl)
      + (MultLoop_acc_917_nl) + (MultLoop_acc_916_nl);
  assign nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8959:8952]));
  assign MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8967:8960]));
  assign MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_915_nl = (readslicef_29_22_7((MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_915_nl = nl_MultLoop_acc_915_nl[21:0];
  assign nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8975:8968]));
  assign MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8983:8976]));
  assign MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_914_nl = (readslicef_29_22_7((MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_914_nl = nl_MultLoop_acc_914_nl[21:0];
  assign nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8991:8984]));
  assign MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8999:8992]));
  assign MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_913_nl = (readslicef_29_22_7((MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_913_nl = nl_MultLoop_acc_913_nl[21:0];
  assign nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9007:9000]));
  assign MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9015:9008]));
  assign MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_912_nl = (readslicef_29_22_7((MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_912_nl = nl_MultLoop_acc_912_nl[21:0];
  assign nl_MultLoop_acc_999_itm_1  = (MultLoop_acc_915_nl) + (MultLoop_acc_914_nl)
      + (MultLoop_acc_913_nl) + (MultLoop_acc_912_nl);
  assign nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9023:9016]));
  assign MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9031:9024]));
  assign MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_911_nl = (readslicef_29_22_7((MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_911_nl = nl_MultLoop_acc_911_nl[21:0];
  assign nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9039:9032]));
  assign MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9047:9040]));
  assign MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_910_nl = (readslicef_29_22_7((MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_910_nl = nl_MultLoop_acc_910_nl[21:0];
  assign nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9055:9048]));
  assign MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9063:9056]));
  assign MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_909_nl = (readslicef_29_22_7((MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_909_nl = nl_MultLoop_acc_909_nl[21:0];
  assign nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9071:9064]));
  assign MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9079:9072]));
  assign MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_908_nl = (readslicef_29_22_7((MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_908_nl = nl_MultLoop_acc_908_nl[21:0];
  assign nl_MultLoop_acc_998_itm_1  = (MultLoop_acc_911_nl) + (MultLoop_acc_910_nl)
      + (MultLoop_acc_909_nl) + (MultLoop_acc_908_nl);
  assign nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9087:9080]));
  assign MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9095:9088]));
  assign MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_907_nl = (readslicef_29_22_7((MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_907_nl = nl_MultLoop_acc_907_nl[21:0];
  assign nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9103:9096]));
  assign MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9111:9104]));
  assign MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_906_nl = (readslicef_29_22_7((MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_906_nl = nl_MultLoop_acc_906_nl[21:0];
  assign nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9119:9112]));
  assign MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9127:9120]));
  assign MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_905_nl = (readslicef_29_22_7((MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_905_nl = nl_MultLoop_acc_905_nl[21:0];
  assign nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9135:9128]));
  assign MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9143:9136]));
  assign MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_904_nl = (readslicef_29_22_7((MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_904_nl = nl_MultLoop_acc_904_nl[21:0];
  assign nl_MultLoop_acc_997_itm_1  = (MultLoop_acc_907_nl) + (MultLoop_acc_906_nl)
      + (MultLoop_acc_905_nl) + (MultLoop_acc_904_nl);
  assign nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9151:9144]));
  assign MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9159:9152]));
  assign MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_903_nl = (readslicef_29_22_7((MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_903_nl = nl_MultLoop_acc_903_nl[21:0];
  assign nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9167:9160]));
  assign MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9175:9168]));
  assign MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_902_nl = (readslicef_29_22_7((MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_902_nl = nl_MultLoop_acc_902_nl[21:0];
  assign nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9183:9176]));
  assign MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9191:9184]));
  assign MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_901_nl = (readslicef_29_22_7((MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_901_nl = nl_MultLoop_acc_901_nl[21:0];
  assign nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9199:9192]));
  assign MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9207:9200]));
  assign MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_900_nl = (readslicef_29_22_7((MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_900_nl = nl_MultLoop_acc_900_nl[21:0];
  assign nl_MultLoop_acc_996_itm_1  = (MultLoop_acc_903_nl) + (MultLoop_acc_902_nl)
      + (MultLoop_acc_901_nl) + (MultLoop_acc_900_nl);
  assign nl_MultLoop_acc_1286_nl = (MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[63:56]);
  assign MultLoop_acc_1286_nl = nl_MultLoop_acc_1286_nl[10:0];
  assign nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[7175:7168]));
  assign MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_836_nl = ({(MultLoop_acc_1286_nl) , (MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_836_nl = nl_MultLoop_acc_836_nl[21:0];
  assign nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7183:7176]));
  assign MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7191:7184]));
  assign MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_835_nl = (readslicef_29_22_7((MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_835_nl = nl_MultLoop_acc_835_nl[21:0];
  assign nl_MultLoop_acc_868_nl = (MultLoop_acc_836_nl) + (MultLoop_acc_835_nl);
  assign MultLoop_acc_868_nl = nl_MultLoop_acc_868_nl[21:0];
  assign nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7199:7192]));
  assign MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7207:7200]));
  assign MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_834_nl = (readslicef_29_22_7((MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_834_nl = nl_MultLoop_acc_834_nl[21:0];
  assign nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7215:7208]));
  assign MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7223:7216]));
  assign MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_833_nl = (readslicef_29_22_7((MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_833_nl = nl_MultLoop_acc_833_nl[21:0];
  assign nl_MultLoop_acc_867_nl = (MultLoop_acc_834_nl) + (MultLoop_acc_833_nl);
  assign MultLoop_acc_867_nl = nl_MultLoop_acc_867_nl[21:0];
  assign nl_MultLoop_acc_884_itm_1  = (MultLoop_acc_868_nl) + (MultLoop_acc_867_nl);
  assign nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7231:7224]));
  assign MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7239:7232]));
  assign MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_832_nl = (readslicef_29_22_7((MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_832_nl = nl_MultLoop_acc_832_nl[21:0];
  assign nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7247:7240]));
  assign MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7255:7248]));
  assign MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_831_nl = (readslicef_29_22_7((MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_831_nl = nl_MultLoop_acc_831_nl[21:0];
  assign nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7263:7256]));
  assign MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7271:7264]));
  assign MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_830_nl = (readslicef_29_22_7((MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_830_nl = nl_MultLoop_acc_830_nl[21:0];
  assign nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7279:7272]));
  assign MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7287:7280]));
  assign MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_829_nl = (readslicef_29_22_7((MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_829_nl = nl_MultLoop_acc_829_nl[21:0];
  assign nl_MultLoop_acc_883_itm_1  = (MultLoop_acc_832_nl) + (MultLoop_acc_831_nl)
      + (MultLoop_acc_830_nl) + (MultLoop_acc_829_nl);
  assign nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7295:7288]));
  assign MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7303:7296]));
  assign MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_828_nl = (readslicef_29_22_7((MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_828_nl = nl_MultLoop_acc_828_nl[21:0];
  assign nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7311:7304]));
  assign MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7319:7312]));
  assign MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_827_nl = (readslicef_29_22_7((MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_827_nl = nl_MultLoop_acc_827_nl[21:0];
  assign nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7327:7320]));
  assign MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7335:7328]));
  assign MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_826_nl = (readslicef_29_22_7((MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_826_nl = nl_MultLoop_acc_826_nl[21:0];
  assign nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7343:7336]));
  assign MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7351:7344]));
  assign MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_825_nl = (readslicef_29_22_7((MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_825_nl = nl_MultLoop_acc_825_nl[21:0];
  assign nl_MultLoop_acc_882_itm_1  = (MultLoop_acc_828_nl) + (MultLoop_acc_827_nl)
      + (MultLoop_acc_826_nl) + (MultLoop_acc_825_nl);
  assign nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7359:7352]));
  assign MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7367:7360]));
  assign MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_824_nl = (readslicef_29_22_7((MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_824_nl = nl_MultLoop_acc_824_nl[21:0];
  assign nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7375:7368]));
  assign MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7383:7376]));
  assign MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_823_nl = (readslicef_29_22_7((MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_823_nl = nl_MultLoop_acc_823_nl[21:0];
  assign nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7391:7384]));
  assign MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7399:7392]));
  assign MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_822_nl = (readslicef_29_22_7((MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_822_nl = nl_MultLoop_acc_822_nl[21:0];
  assign nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7407:7400]));
  assign MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7415:7408]));
  assign MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_821_nl = (readslicef_29_22_7((MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_821_nl = nl_MultLoop_acc_821_nl[21:0];
  assign nl_MultLoop_acc_881_itm_1  = (MultLoop_acc_824_nl) + (MultLoop_acc_823_nl)
      + (MultLoop_acc_822_nl) + (MultLoop_acc_821_nl);
  assign nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7423:7416]));
  assign MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7431:7424]));
  assign MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_820_nl = (readslicef_29_22_7((MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_820_nl = nl_MultLoop_acc_820_nl[21:0];
  assign nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7439:7432]));
  assign MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7447:7440]));
  assign MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_819_nl = (readslicef_29_22_7((MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_819_nl = nl_MultLoop_acc_819_nl[21:0];
  assign nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7455:7448]));
  assign MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7463:7456]));
  assign MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_818_nl = (readslicef_29_22_7((MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_818_nl = nl_MultLoop_acc_818_nl[21:0];
  assign nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7471:7464]));
  assign MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7479:7472]));
  assign MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_817_nl = (readslicef_29_22_7((MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_817_nl = nl_MultLoop_acc_817_nl[21:0];
  assign nl_MultLoop_acc_880_itm_1  = (MultLoop_acc_820_nl) + (MultLoop_acc_819_nl)
      + (MultLoop_acc_818_nl) + (MultLoop_acc_817_nl);
  assign nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7487:7480]));
  assign MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7495:7488]));
  assign MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_816_nl = (readslicef_29_22_7((MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_816_nl = nl_MultLoop_acc_816_nl[21:0];
  assign nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7503:7496]));
  assign MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7511:7504]));
  assign MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_815_nl = (readslicef_29_22_7((MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_815_nl = nl_MultLoop_acc_815_nl[21:0];
  assign nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7519:7512]));
  assign MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7527:7520]));
  assign MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_814_nl = (readslicef_29_22_7((MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_814_nl = nl_MultLoop_acc_814_nl[21:0];
  assign nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7535:7528]));
  assign MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7543:7536]));
  assign MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_813_nl = (readslicef_29_22_7((MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_813_nl = nl_MultLoop_acc_813_nl[21:0];
  assign nl_MultLoop_acc_879_itm_1  = (MultLoop_acc_816_nl) + (MultLoop_acc_815_nl)
      + (MultLoop_acc_814_nl) + (MultLoop_acc_813_nl);
  assign nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7551:7544]));
  assign MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7559:7552]));
  assign MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_812_nl = (readslicef_29_22_7((MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_812_nl = nl_MultLoop_acc_812_nl[21:0];
  assign nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7567:7560]));
  assign MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7575:7568]));
  assign MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_811_nl = (readslicef_29_22_7((MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_811_nl = nl_MultLoop_acc_811_nl[21:0];
  assign nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7583:7576]));
  assign MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7591:7584]));
  assign MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_810_nl = (readslicef_29_22_7((MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_810_nl = nl_MultLoop_acc_810_nl[21:0];
  assign nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7599:7592]));
  assign MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7607:7600]));
  assign MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_809_nl = (readslicef_29_22_7((MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_809_nl = nl_MultLoop_acc_809_nl[21:0];
  assign nl_MultLoop_acc_878_itm_1  = (MultLoop_acc_812_nl) + (MultLoop_acc_811_nl)
      + (MultLoop_acc_810_nl) + (MultLoop_acc_809_nl);
  assign nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7615:7608]));
  assign MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7623:7616]));
  assign MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_808_nl = (readslicef_29_22_7((MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_808_nl = nl_MultLoop_acc_808_nl[21:0];
  assign nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7631:7624]));
  assign MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7639:7632]));
  assign MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_807_nl = (readslicef_29_22_7((MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_807_nl = nl_MultLoop_acc_807_nl[21:0];
  assign nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7647:7640]));
  assign MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7655:7648]));
  assign MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_806_nl = (readslicef_29_22_7((MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_806_nl = nl_MultLoop_acc_806_nl[21:0];
  assign nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7663:7656]));
  assign MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7671:7664]));
  assign MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_805_nl = (readslicef_29_22_7((MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_805_nl = nl_MultLoop_acc_805_nl[21:0];
  assign nl_MultLoop_acc_877_itm_1  = (MultLoop_acc_808_nl) + (MultLoop_acc_807_nl)
      + (MultLoop_acc_806_nl) + (MultLoop_acc_805_nl);
  assign nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7679:7672]));
  assign MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7687:7680]));
  assign MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_804_nl = (readslicef_29_22_7((MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_804_nl = nl_MultLoop_acc_804_nl[21:0];
  assign nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7695:7688]));
  assign MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7703:7696]));
  assign MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_803_nl = (readslicef_29_22_7((MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_803_nl = nl_MultLoop_acc_803_nl[21:0];
  assign nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7711:7704]));
  assign MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7719:7712]));
  assign MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_802_nl = (readslicef_29_22_7((MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_802_nl = nl_MultLoop_acc_802_nl[21:0];
  assign nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7727:7720]));
  assign MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7735:7728]));
  assign MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_801_nl = (readslicef_29_22_7((MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_801_nl = nl_MultLoop_acc_801_nl[21:0];
  assign nl_MultLoop_acc_876_itm_1  = (MultLoop_acc_804_nl) + (MultLoop_acc_803_nl)
      + (MultLoop_acc_802_nl) + (MultLoop_acc_801_nl);
  assign nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7743:7736]));
  assign MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7751:7744]));
  assign MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_800_nl = (readslicef_29_22_7((MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_800_nl = nl_MultLoop_acc_800_nl[21:0];
  assign nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7759:7752]));
  assign MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7767:7760]));
  assign MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_799_nl = (readslicef_29_22_7((MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_799_nl = nl_MultLoop_acc_799_nl[21:0];
  assign nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7775:7768]));
  assign MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7783:7776]));
  assign MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_798_nl = (readslicef_29_22_7((MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_798_nl = nl_MultLoop_acc_798_nl[21:0];
  assign nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7791:7784]));
  assign MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7799:7792]));
  assign MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_797_nl = (readslicef_29_22_7((MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_797_nl = nl_MultLoop_acc_797_nl[21:0];
  assign nl_MultLoop_acc_875_itm_1  = (MultLoop_acc_800_nl) + (MultLoop_acc_799_nl)
      + (MultLoop_acc_798_nl) + (MultLoop_acc_797_nl);
  assign nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7807:7800]));
  assign MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7815:7808]));
  assign MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_796_nl = (readslicef_29_22_7((MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_796_nl = nl_MultLoop_acc_796_nl[21:0];
  assign nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7823:7816]));
  assign MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7831:7824]));
  assign MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_795_nl = (readslicef_29_22_7((MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_795_nl = nl_MultLoop_acc_795_nl[21:0];
  assign nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7839:7832]));
  assign MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7847:7840]));
  assign MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_794_nl = (readslicef_29_22_7((MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_794_nl = nl_MultLoop_acc_794_nl[21:0];
  assign nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7855:7848]));
  assign MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7863:7856]));
  assign MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_793_nl = (readslicef_29_22_7((MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_793_nl = nl_MultLoop_acc_793_nl[21:0];
  assign nl_MultLoop_acc_874_itm_1  = (MultLoop_acc_796_nl) + (MultLoop_acc_795_nl)
      + (MultLoop_acc_794_nl) + (MultLoop_acc_793_nl);
  assign nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7871:7864]));
  assign MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7879:7872]));
  assign MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_792_nl = (readslicef_29_22_7((MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_792_nl = nl_MultLoop_acc_792_nl[21:0];
  assign nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7887:7880]));
  assign MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7895:7888]));
  assign MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_791_nl = (readslicef_29_22_7((MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_791_nl = nl_MultLoop_acc_791_nl[21:0];
  assign nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7903:7896]));
  assign MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7911:7904]));
  assign MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_790_nl = (readslicef_29_22_7((MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_790_nl = nl_MultLoop_acc_790_nl[21:0];
  assign nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7919:7912]));
  assign MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7927:7920]));
  assign MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_789_nl = (readslicef_29_22_7((MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_789_nl = nl_MultLoop_acc_789_nl[21:0];
  assign nl_MultLoop_acc_873_itm_1  = (MultLoop_acc_792_nl) + (MultLoop_acc_791_nl)
      + (MultLoop_acc_790_nl) + (MultLoop_acc_789_nl);
  assign nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7935:7928]));
  assign MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7943:7936]));
  assign MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_788_nl = (readslicef_29_22_7((MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_788_nl = nl_MultLoop_acc_788_nl[21:0];
  assign nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7951:7944]));
  assign MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7959:7952]));
  assign MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_787_nl = (readslicef_29_22_7((MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_787_nl = nl_MultLoop_acc_787_nl[21:0];
  assign nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7967:7960]));
  assign MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7975:7968]));
  assign MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_786_nl = (readslicef_29_22_7((MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_786_nl = nl_MultLoop_acc_786_nl[21:0];
  assign nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7983:7976]));
  assign MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7991:7984]));
  assign MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_785_nl = (readslicef_29_22_7((MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_785_nl = nl_MultLoop_acc_785_nl[21:0];
  assign nl_MultLoop_acc_872_itm_1  = (MultLoop_acc_788_nl) + (MultLoop_acc_787_nl)
      + (MultLoop_acc_786_nl) + (MultLoop_acc_785_nl);
  assign nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7999:7992]));
  assign MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8007:8000]));
  assign MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_784_nl = (readslicef_29_22_7((MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_784_nl = nl_MultLoop_acc_784_nl[21:0];
  assign nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8015:8008]));
  assign MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8023:8016]));
  assign MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_783_nl = (readslicef_29_22_7((MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_783_nl = nl_MultLoop_acc_783_nl[21:0];
  assign nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8031:8024]));
  assign MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8039:8032]));
  assign MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_782_nl = (readslicef_29_22_7((MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_782_nl = nl_MultLoop_acc_782_nl[21:0];
  assign nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8047:8040]));
  assign MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8055:8048]));
  assign MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_781_nl = (readslicef_29_22_7((MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_781_nl = nl_MultLoop_acc_781_nl[21:0];
  assign nl_MultLoop_acc_871_itm_1  = (MultLoop_acc_784_nl) + (MultLoop_acc_783_nl)
      + (MultLoop_acc_782_nl) + (MultLoop_acc_781_nl);
  assign nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8063:8056]));
  assign MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8071:8064]));
  assign MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_780_nl = (readslicef_29_22_7((MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_780_nl = nl_MultLoop_acc_780_nl[21:0];
  assign nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8079:8072]));
  assign MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8087:8080]));
  assign MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_779_nl = (readslicef_29_22_7((MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_779_nl = nl_MultLoop_acc_779_nl[21:0];
  assign nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8095:8088]));
  assign MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8103:8096]));
  assign MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_778_nl = (readslicef_29_22_7((MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_778_nl = nl_MultLoop_acc_778_nl[21:0];
  assign nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8111:8104]));
  assign MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8119:8112]));
  assign MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_777_nl = (readslicef_29_22_7((MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_777_nl = nl_MultLoop_acc_777_nl[21:0];
  assign nl_MultLoop_acc_870_itm_1  = (MultLoop_acc_780_nl) + (MultLoop_acc_779_nl)
      + (MultLoop_acc_778_nl) + (MultLoop_acc_777_nl);
  assign nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8127:8120]));
  assign MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8135:8128]));
  assign MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_776_nl = (readslicef_29_22_7((MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_776_nl = nl_MultLoop_acc_776_nl[21:0];
  assign nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8143:8136]));
  assign MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8151:8144]));
  assign MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_775_nl = (readslicef_29_22_7((MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_775_nl = nl_MultLoop_acc_775_nl[21:0];
  assign nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8159:8152]));
  assign MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8167:8160]));
  assign MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_774_nl = (readslicef_29_22_7((MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_774_nl = nl_MultLoop_acc_774_nl[21:0];
  assign nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8175:8168]));
  assign MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8183:8176]));
  assign MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_773_nl = (readslicef_29_22_7((MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_773_nl = nl_MultLoop_acc_773_nl[21:0];
  assign nl_MultLoop_acc_869_itm_1  = (MultLoop_acc_776_nl) + (MultLoop_acc_775_nl)
      + (MultLoop_acc_774_nl) + (MultLoop_acc_773_nl);
  assign nl_MultLoop_acc_1285_nl = (MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[55:48]);
  assign MultLoop_acc_1285_nl = nl_MultLoop_acc_1285_nl[10:0];
  assign nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[6151:6144]));
  assign MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_709_nl = ({(MultLoop_acc_1285_nl) , (MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_709_nl = nl_MultLoop_acc_709_nl[21:0];
  assign nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6159:6152]));
  assign MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6167:6160]));
  assign MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_708_nl = (readslicef_29_22_7((MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_708_nl = nl_MultLoop_acc_708_nl[21:0];
  assign nl_MultLoop_acc_741_nl = (MultLoop_acc_709_nl) + (MultLoop_acc_708_nl);
  assign MultLoop_acc_741_nl = nl_MultLoop_acc_741_nl[21:0];
  assign nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6175:6168]));
  assign MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6183:6176]));
  assign MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_707_nl = (readslicef_29_22_7((MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_707_nl = nl_MultLoop_acc_707_nl[21:0];
  assign nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6191:6184]));
  assign MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6199:6192]));
  assign MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_706_nl = (readslicef_29_22_7((MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_706_nl = nl_MultLoop_acc_706_nl[21:0];
  assign nl_MultLoop_acc_740_nl = (MultLoop_acc_707_nl) + (MultLoop_acc_706_nl);
  assign MultLoop_acc_740_nl = nl_MultLoop_acc_740_nl[21:0];
  assign nl_MultLoop_acc_757_itm_1  = (MultLoop_acc_741_nl) + (MultLoop_acc_740_nl);
  assign nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6207:6200]));
  assign MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6215:6208]));
  assign MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_705_nl = (readslicef_29_22_7((MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_705_nl = nl_MultLoop_acc_705_nl[21:0];
  assign nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6223:6216]));
  assign MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6231:6224]));
  assign MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_704_nl = (readslicef_29_22_7((MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_704_nl = nl_MultLoop_acc_704_nl[21:0];
  assign nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6239:6232]));
  assign MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6247:6240]));
  assign MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_703_nl = (readslicef_29_22_7((MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_703_nl = nl_MultLoop_acc_703_nl[21:0];
  assign nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6255:6248]));
  assign MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6263:6256]));
  assign MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_702_nl = (readslicef_29_22_7((MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_702_nl = nl_MultLoop_acc_702_nl[21:0];
  assign nl_MultLoop_acc_756_itm_1  = (MultLoop_acc_705_nl) + (MultLoop_acc_704_nl)
      + (MultLoop_acc_703_nl) + (MultLoop_acc_702_nl);
  assign nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6271:6264]));
  assign MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6279:6272]));
  assign MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_701_nl = (readslicef_29_22_7((MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_701_nl = nl_MultLoop_acc_701_nl[21:0];
  assign nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6287:6280]));
  assign MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6295:6288]));
  assign MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_700_nl = (readslicef_29_22_7((MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_700_nl = nl_MultLoop_acc_700_nl[21:0];
  assign nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6303:6296]));
  assign MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6311:6304]));
  assign MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_699_nl = (readslicef_29_22_7((MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_699_nl = nl_MultLoop_acc_699_nl[21:0];
  assign nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6319:6312]));
  assign MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6327:6320]));
  assign MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_698_nl = (readslicef_29_22_7((MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_698_nl = nl_MultLoop_acc_698_nl[21:0];
  assign nl_MultLoop_acc_755_itm_1  = (MultLoop_acc_701_nl) + (MultLoop_acc_700_nl)
      + (MultLoop_acc_699_nl) + (MultLoop_acc_698_nl);
  assign nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6335:6328]));
  assign MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6343:6336]));
  assign MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_697_nl = (readslicef_29_22_7((MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_697_nl = nl_MultLoop_acc_697_nl[21:0];
  assign nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6351:6344]));
  assign MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6359:6352]));
  assign MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_696_nl = (readslicef_29_22_7((MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_696_nl = nl_MultLoop_acc_696_nl[21:0];
  assign nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6367:6360]));
  assign MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6375:6368]));
  assign MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_695_nl = (readslicef_29_22_7((MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_695_nl = nl_MultLoop_acc_695_nl[21:0];
  assign nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6383:6376]));
  assign MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6391:6384]));
  assign MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_694_nl = (readslicef_29_22_7((MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_694_nl = nl_MultLoop_acc_694_nl[21:0];
  assign nl_MultLoop_acc_754_itm_1  = (MultLoop_acc_697_nl) + (MultLoop_acc_696_nl)
      + (MultLoop_acc_695_nl) + (MultLoop_acc_694_nl);
  assign nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6399:6392]));
  assign MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6407:6400]));
  assign MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_693_nl = (readslicef_29_22_7((MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_693_nl = nl_MultLoop_acc_693_nl[21:0];
  assign nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6415:6408]));
  assign MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6423:6416]));
  assign MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_692_nl = (readslicef_29_22_7((MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_692_nl = nl_MultLoop_acc_692_nl[21:0];
  assign nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6431:6424]));
  assign MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6439:6432]));
  assign MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_691_nl = (readslicef_29_22_7((MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_691_nl = nl_MultLoop_acc_691_nl[21:0];
  assign nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6447:6440]));
  assign MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6455:6448]));
  assign MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_690_nl = (readslicef_29_22_7((MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_690_nl = nl_MultLoop_acc_690_nl[21:0];
  assign nl_MultLoop_acc_753_itm_1  = (MultLoop_acc_693_nl) + (MultLoop_acc_692_nl)
      + (MultLoop_acc_691_nl) + (MultLoop_acc_690_nl);
  assign nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6463:6456]));
  assign MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6471:6464]));
  assign MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_689_nl = (readslicef_29_22_7((MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_689_nl = nl_MultLoop_acc_689_nl[21:0];
  assign nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6479:6472]));
  assign MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6487:6480]));
  assign MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_688_nl = (readslicef_29_22_7((MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_688_nl = nl_MultLoop_acc_688_nl[21:0];
  assign nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6495:6488]));
  assign MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6503:6496]));
  assign MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_687_nl = (readslicef_29_22_7((MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_687_nl = nl_MultLoop_acc_687_nl[21:0];
  assign nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6511:6504]));
  assign MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6519:6512]));
  assign MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_686_nl = (readslicef_29_22_7((MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_686_nl = nl_MultLoop_acc_686_nl[21:0];
  assign nl_MultLoop_acc_752_itm_1  = (MultLoop_acc_689_nl) + (MultLoop_acc_688_nl)
      + (MultLoop_acc_687_nl) + (MultLoop_acc_686_nl);
  assign nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6527:6520]));
  assign MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6535:6528]));
  assign MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_685_nl = (readslicef_29_22_7((MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_685_nl = nl_MultLoop_acc_685_nl[21:0];
  assign nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6543:6536]));
  assign MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6551:6544]));
  assign MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_684_nl = (readslicef_29_22_7((MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_684_nl = nl_MultLoop_acc_684_nl[21:0];
  assign nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6559:6552]));
  assign MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6567:6560]));
  assign MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_683_nl = (readslicef_29_22_7((MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_683_nl = nl_MultLoop_acc_683_nl[21:0];
  assign nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6575:6568]));
  assign MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6583:6576]));
  assign MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_682_nl = (readslicef_29_22_7((MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_682_nl = nl_MultLoop_acc_682_nl[21:0];
  assign nl_MultLoop_acc_751_itm_1  = (MultLoop_acc_685_nl) + (MultLoop_acc_684_nl)
      + (MultLoop_acc_683_nl) + (MultLoop_acc_682_nl);
  assign nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6591:6584]));
  assign MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6599:6592]));
  assign MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_681_nl = (readslicef_29_22_7((MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_681_nl = nl_MultLoop_acc_681_nl[21:0];
  assign nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6607:6600]));
  assign MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6615:6608]));
  assign MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_680_nl = (readslicef_29_22_7((MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_680_nl = nl_MultLoop_acc_680_nl[21:0];
  assign nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6623:6616]));
  assign MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6631:6624]));
  assign MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_679_nl = (readslicef_29_22_7((MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_679_nl = nl_MultLoop_acc_679_nl[21:0];
  assign nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6639:6632]));
  assign MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6647:6640]));
  assign MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_678_nl = (readslicef_29_22_7((MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_678_nl = nl_MultLoop_acc_678_nl[21:0];
  assign nl_MultLoop_acc_750_itm_1  = (MultLoop_acc_681_nl) + (MultLoop_acc_680_nl)
      + (MultLoop_acc_679_nl) + (MultLoop_acc_678_nl);
  assign nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6655:6648]));
  assign MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6663:6656]));
  assign MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_677_nl = (readslicef_29_22_7((MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_677_nl = nl_MultLoop_acc_677_nl[21:0];
  assign nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6671:6664]));
  assign MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6679:6672]));
  assign MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_676_nl = (readslicef_29_22_7((MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_676_nl = nl_MultLoop_acc_676_nl[21:0];
  assign nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6687:6680]));
  assign MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6695:6688]));
  assign MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_675_nl = (readslicef_29_22_7((MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_675_nl = nl_MultLoop_acc_675_nl[21:0];
  assign nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6703:6696]));
  assign MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6711:6704]));
  assign MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_674_nl = (readslicef_29_22_7((MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_674_nl = nl_MultLoop_acc_674_nl[21:0];
  assign nl_MultLoop_acc_749_itm_1  = (MultLoop_acc_677_nl) + (MultLoop_acc_676_nl)
      + (MultLoop_acc_675_nl) + (MultLoop_acc_674_nl);
  assign nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6719:6712]));
  assign MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6727:6720]));
  assign MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_673_nl = (readslicef_29_22_7((MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_673_nl = nl_MultLoop_acc_673_nl[21:0];
  assign nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6735:6728]));
  assign MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6743:6736]));
  assign MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_672_nl = (readslicef_29_22_7((MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_672_nl = nl_MultLoop_acc_672_nl[21:0];
  assign nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6751:6744]));
  assign MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6759:6752]));
  assign MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_671_nl = (readslicef_29_22_7((MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_671_nl = nl_MultLoop_acc_671_nl[21:0];
  assign nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6767:6760]));
  assign MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6775:6768]));
  assign MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_670_nl = (readslicef_29_22_7((MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_670_nl = nl_MultLoop_acc_670_nl[21:0];
  assign nl_MultLoop_acc_748_itm_1  = (MultLoop_acc_673_nl) + (MultLoop_acc_672_nl)
      + (MultLoop_acc_671_nl) + (MultLoop_acc_670_nl);
  assign nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6783:6776]));
  assign MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6791:6784]));
  assign MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_669_nl = (readslicef_29_22_7((MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_669_nl = nl_MultLoop_acc_669_nl[21:0];
  assign nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6799:6792]));
  assign MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6807:6800]));
  assign MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_668_nl = (readslicef_29_22_7((MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_668_nl = nl_MultLoop_acc_668_nl[21:0];
  assign nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6815:6808]));
  assign MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6823:6816]));
  assign MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_667_nl = (readslicef_29_22_7((MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_667_nl = nl_MultLoop_acc_667_nl[21:0];
  assign nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6831:6824]));
  assign MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6839:6832]));
  assign MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_666_nl = (readslicef_29_22_7((MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_666_nl = nl_MultLoop_acc_666_nl[21:0];
  assign nl_MultLoop_acc_747_itm_1  = (MultLoop_acc_669_nl) + (MultLoop_acc_668_nl)
      + (MultLoop_acc_667_nl) + (MultLoop_acc_666_nl);
  assign nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6847:6840]));
  assign MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6855:6848]));
  assign MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_665_nl = (readslicef_29_22_7((MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_665_nl = nl_MultLoop_acc_665_nl[21:0];
  assign nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6863:6856]));
  assign MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6871:6864]));
  assign MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_664_nl = (readslicef_29_22_7((MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_664_nl = nl_MultLoop_acc_664_nl[21:0];
  assign nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6879:6872]));
  assign MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6887:6880]));
  assign MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_663_nl = (readslicef_29_22_7((MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_663_nl = nl_MultLoop_acc_663_nl[21:0];
  assign nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6895:6888]));
  assign MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6903:6896]));
  assign MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_662_nl = (readslicef_29_22_7((MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_662_nl = nl_MultLoop_acc_662_nl[21:0];
  assign nl_MultLoop_acc_746_itm_1  = (MultLoop_acc_665_nl) + (MultLoop_acc_664_nl)
      + (MultLoop_acc_663_nl) + (MultLoop_acc_662_nl);
  assign nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6911:6904]));
  assign MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6919:6912]));
  assign MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_661_nl = (readslicef_29_22_7((MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_661_nl = nl_MultLoop_acc_661_nl[21:0];
  assign nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6927:6920]));
  assign MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6935:6928]));
  assign MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_660_nl = (readslicef_29_22_7((MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_660_nl = nl_MultLoop_acc_660_nl[21:0];
  assign nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6943:6936]));
  assign MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6951:6944]));
  assign MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_659_nl = (readslicef_29_22_7((MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_659_nl = nl_MultLoop_acc_659_nl[21:0];
  assign nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6959:6952]));
  assign MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6967:6960]));
  assign MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_658_nl = (readslicef_29_22_7((MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_658_nl = nl_MultLoop_acc_658_nl[21:0];
  assign nl_MultLoop_acc_745_itm_1  = (MultLoop_acc_661_nl) + (MultLoop_acc_660_nl)
      + (MultLoop_acc_659_nl) + (MultLoop_acc_658_nl);
  assign nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6975:6968]));
  assign MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6983:6976]));
  assign MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_657_nl = (readslicef_29_22_7((MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_657_nl = nl_MultLoop_acc_657_nl[21:0];
  assign nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6991:6984]));
  assign MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6999:6992]));
  assign MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_656_nl = (readslicef_29_22_7((MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_656_nl = nl_MultLoop_acc_656_nl[21:0];
  assign nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7007:7000]));
  assign MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7015:7008]));
  assign MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_655_nl = (readslicef_29_22_7((MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_655_nl = nl_MultLoop_acc_655_nl[21:0];
  assign nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7023:7016]));
  assign MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7031:7024]));
  assign MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_654_nl = (readslicef_29_22_7((MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_654_nl = nl_MultLoop_acc_654_nl[21:0];
  assign nl_MultLoop_acc_744_itm_1  = (MultLoop_acc_657_nl) + (MultLoop_acc_656_nl)
      + (MultLoop_acc_655_nl) + (MultLoop_acc_654_nl);
  assign nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7039:7032]));
  assign MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7047:7040]));
  assign MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_653_nl = (readslicef_29_22_7((MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_653_nl = nl_MultLoop_acc_653_nl[21:0];
  assign nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7055:7048]));
  assign MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7063:7056]));
  assign MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_652_nl = (readslicef_29_22_7((MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_652_nl = nl_MultLoop_acc_652_nl[21:0];
  assign nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7071:7064]));
  assign MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7079:7072]));
  assign MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_651_nl = (readslicef_29_22_7((MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_651_nl = nl_MultLoop_acc_651_nl[21:0];
  assign nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7087:7080]));
  assign MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7095:7088]));
  assign MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_650_nl = (readslicef_29_22_7((MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_650_nl = nl_MultLoop_acc_650_nl[21:0];
  assign nl_MultLoop_acc_743_itm_1  = (MultLoop_acc_653_nl) + (MultLoop_acc_652_nl)
      + (MultLoop_acc_651_nl) + (MultLoop_acc_650_nl);
  assign nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7103:7096]));
  assign MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7111:7104]));
  assign MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_649_nl = (readslicef_29_22_7((MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_649_nl = nl_MultLoop_acc_649_nl[21:0];
  assign nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7119:7112]));
  assign MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7127:7120]));
  assign MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_648_nl = (readslicef_29_22_7((MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_648_nl = nl_MultLoop_acc_648_nl[21:0];
  assign nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7135:7128]));
  assign MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7143:7136]));
  assign MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_647_nl = (readslicef_29_22_7((MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_647_nl = nl_MultLoop_acc_647_nl[21:0];
  assign nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7151:7144]));
  assign MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7159:7152]));
  assign MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_646_nl = (readslicef_29_22_7((MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_646_nl = nl_MultLoop_acc_646_nl[21:0];
  assign nl_MultLoop_acc_742_itm_1  = (MultLoop_acc_649_nl) + (MultLoop_acc_648_nl)
      + (MultLoop_acc_647_nl) + (MultLoop_acc_646_nl);
  assign nl_MultLoop_acc_1284_nl = (MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[47:40]);
  assign MultLoop_acc_1284_nl = nl_MultLoop_acc_1284_nl[10:0];
  assign nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[5127:5120]));
  assign MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_582_nl = ({(MultLoop_acc_1284_nl) , (MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_582_nl = nl_MultLoop_acc_582_nl[21:0];
  assign nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5135:5128]));
  assign MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5143:5136]));
  assign MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_581_nl = (readslicef_29_22_7((MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_581_nl = nl_MultLoop_acc_581_nl[21:0];
  assign nl_MultLoop_acc_614_nl = (MultLoop_acc_582_nl) + (MultLoop_acc_581_nl);
  assign MultLoop_acc_614_nl = nl_MultLoop_acc_614_nl[21:0];
  assign nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5151:5144]));
  assign MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5159:5152]));
  assign MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_580_nl = (readslicef_29_22_7((MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_580_nl = nl_MultLoop_acc_580_nl[21:0];
  assign nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5167:5160]));
  assign MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5175:5168]));
  assign MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_579_nl = (readslicef_29_22_7((MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_579_nl = nl_MultLoop_acc_579_nl[21:0];
  assign nl_MultLoop_acc_613_nl = (MultLoop_acc_580_nl) + (MultLoop_acc_579_nl);
  assign MultLoop_acc_613_nl = nl_MultLoop_acc_613_nl[21:0];
  assign nl_MultLoop_acc_630_itm_1  = (MultLoop_acc_614_nl) + (MultLoop_acc_613_nl);
  assign nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5183:5176]));
  assign MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5191:5184]));
  assign MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_578_nl = (readslicef_29_22_7((MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_578_nl = nl_MultLoop_acc_578_nl[21:0];
  assign nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5199:5192]));
  assign MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5207:5200]));
  assign MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_577_nl = (readslicef_29_22_7((MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_577_nl = nl_MultLoop_acc_577_nl[21:0];
  assign nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5215:5208]));
  assign MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5223:5216]));
  assign MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_576_nl = (readslicef_29_22_7((MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_576_nl = nl_MultLoop_acc_576_nl[21:0];
  assign nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5231:5224]));
  assign MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5239:5232]));
  assign MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_575_nl = (readslicef_29_22_7((MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_575_nl = nl_MultLoop_acc_575_nl[21:0];
  assign nl_MultLoop_acc_629_itm_1  = (MultLoop_acc_578_nl) + (MultLoop_acc_577_nl)
      + (MultLoop_acc_576_nl) + (MultLoop_acc_575_nl);
  assign nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5247:5240]));
  assign MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5255:5248]));
  assign MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_574_nl = (readslicef_29_22_7((MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_574_nl = nl_MultLoop_acc_574_nl[21:0];
  assign nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5263:5256]));
  assign MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5271:5264]));
  assign MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_573_nl = (readslicef_29_22_7((MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_573_nl = nl_MultLoop_acc_573_nl[21:0];
  assign nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5279:5272]));
  assign MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5287:5280]));
  assign MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_572_nl = (readslicef_29_22_7((MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_572_nl = nl_MultLoop_acc_572_nl[21:0];
  assign nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5295:5288]));
  assign MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5303:5296]));
  assign MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_571_nl = (readslicef_29_22_7((MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_571_nl = nl_MultLoop_acc_571_nl[21:0];
  assign nl_MultLoop_acc_628_itm_1  = (MultLoop_acc_574_nl) + (MultLoop_acc_573_nl)
      + (MultLoop_acc_572_nl) + (MultLoop_acc_571_nl);
  assign nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5311:5304]));
  assign MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5319:5312]));
  assign MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_570_nl = (readslicef_29_22_7((MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_570_nl = nl_MultLoop_acc_570_nl[21:0];
  assign nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5327:5320]));
  assign MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5335:5328]));
  assign MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_569_nl = (readslicef_29_22_7((MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_569_nl = nl_MultLoop_acc_569_nl[21:0];
  assign nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5343:5336]));
  assign MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5351:5344]));
  assign MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_568_nl = (readslicef_29_22_7((MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_568_nl = nl_MultLoop_acc_568_nl[21:0];
  assign nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5359:5352]));
  assign MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5367:5360]));
  assign MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_567_nl = (readslicef_29_22_7((MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_567_nl = nl_MultLoop_acc_567_nl[21:0];
  assign nl_MultLoop_acc_627_itm_1  = (MultLoop_acc_570_nl) + (MultLoop_acc_569_nl)
      + (MultLoop_acc_568_nl) + (MultLoop_acc_567_nl);
  assign nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5375:5368]));
  assign MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5383:5376]));
  assign MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_566_nl = (readslicef_29_22_7((MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_566_nl = nl_MultLoop_acc_566_nl[21:0];
  assign nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5391:5384]));
  assign MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5399:5392]));
  assign MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_565_nl = (readslicef_29_22_7((MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_565_nl = nl_MultLoop_acc_565_nl[21:0];
  assign nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5407:5400]));
  assign MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5415:5408]));
  assign MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_564_nl = (readslicef_29_22_7((MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_564_nl = nl_MultLoop_acc_564_nl[21:0];
  assign nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5423:5416]));
  assign MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5431:5424]));
  assign MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_563_nl = (readslicef_29_22_7((MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_563_nl = nl_MultLoop_acc_563_nl[21:0];
  assign nl_MultLoop_acc_626_itm_1  = (MultLoop_acc_566_nl) + (MultLoop_acc_565_nl)
      + (MultLoop_acc_564_nl) + (MultLoop_acc_563_nl);
  assign nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5439:5432]));
  assign MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5447:5440]));
  assign MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_562_nl = (readslicef_29_22_7((MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_562_nl = nl_MultLoop_acc_562_nl[21:0];
  assign nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5455:5448]));
  assign MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5463:5456]));
  assign MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_561_nl = (readslicef_29_22_7((MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_561_nl = nl_MultLoop_acc_561_nl[21:0];
  assign nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5471:5464]));
  assign MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5479:5472]));
  assign MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_560_nl = (readslicef_29_22_7((MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_560_nl = nl_MultLoop_acc_560_nl[21:0];
  assign nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5487:5480]));
  assign MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5495:5488]));
  assign MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_559_nl = (readslicef_29_22_7((MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_559_nl = nl_MultLoop_acc_559_nl[21:0];
  assign nl_MultLoop_acc_625_itm_1  = (MultLoop_acc_562_nl) + (MultLoop_acc_561_nl)
      + (MultLoop_acc_560_nl) + (MultLoop_acc_559_nl);
  assign nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5503:5496]));
  assign MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5511:5504]));
  assign MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_558_nl = (readslicef_29_22_7((MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_558_nl = nl_MultLoop_acc_558_nl[21:0];
  assign nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5519:5512]));
  assign MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5527:5520]));
  assign MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_557_nl = (readslicef_29_22_7((MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_557_nl = nl_MultLoop_acc_557_nl[21:0];
  assign nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5535:5528]));
  assign MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5543:5536]));
  assign MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_556_nl = (readslicef_29_22_7((MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_556_nl = nl_MultLoop_acc_556_nl[21:0];
  assign nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5551:5544]));
  assign MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5559:5552]));
  assign MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_555_nl = (readslicef_29_22_7((MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_555_nl = nl_MultLoop_acc_555_nl[21:0];
  assign nl_MultLoop_acc_624_itm_1  = (MultLoop_acc_558_nl) + (MultLoop_acc_557_nl)
      + (MultLoop_acc_556_nl) + (MultLoop_acc_555_nl);
  assign nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5567:5560]));
  assign MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5575:5568]));
  assign MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_554_nl = (readslicef_29_22_7((MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_554_nl = nl_MultLoop_acc_554_nl[21:0];
  assign nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5583:5576]));
  assign MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5591:5584]));
  assign MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_553_nl = (readslicef_29_22_7((MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_553_nl = nl_MultLoop_acc_553_nl[21:0];
  assign nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5599:5592]));
  assign MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5607:5600]));
  assign MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_552_nl = (readslicef_29_22_7((MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_552_nl = nl_MultLoop_acc_552_nl[21:0];
  assign nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5615:5608]));
  assign MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5623:5616]));
  assign MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_551_nl = (readslicef_29_22_7((MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_551_nl = nl_MultLoop_acc_551_nl[21:0];
  assign nl_MultLoop_acc_623_itm_1  = (MultLoop_acc_554_nl) + (MultLoop_acc_553_nl)
      + (MultLoop_acc_552_nl) + (MultLoop_acc_551_nl);
  assign nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5631:5624]));
  assign MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5639:5632]));
  assign MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_550_nl = (readslicef_29_22_7((MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_550_nl = nl_MultLoop_acc_550_nl[21:0];
  assign nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5647:5640]));
  assign MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5655:5648]));
  assign MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_549_nl = (readslicef_29_22_7((MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_549_nl = nl_MultLoop_acc_549_nl[21:0];
  assign nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5663:5656]));
  assign MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5671:5664]));
  assign MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_548_nl = (readslicef_29_22_7((MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_548_nl = nl_MultLoop_acc_548_nl[21:0];
  assign nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5679:5672]));
  assign MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5687:5680]));
  assign MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_547_nl = (readslicef_29_22_7((MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_547_nl = nl_MultLoop_acc_547_nl[21:0];
  assign nl_MultLoop_acc_622_itm_1  = (MultLoop_acc_550_nl) + (MultLoop_acc_549_nl)
      + (MultLoop_acc_548_nl) + (MultLoop_acc_547_nl);
  assign nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5695:5688]));
  assign MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5703:5696]));
  assign MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_546_nl = (readslicef_29_22_7((MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_546_nl = nl_MultLoop_acc_546_nl[21:0];
  assign nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5711:5704]));
  assign MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5719:5712]));
  assign MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_545_nl = (readslicef_29_22_7((MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_545_nl = nl_MultLoop_acc_545_nl[21:0];
  assign nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5727:5720]));
  assign MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5735:5728]));
  assign MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_544_nl = (readslicef_29_22_7((MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_544_nl = nl_MultLoop_acc_544_nl[21:0];
  assign nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5743:5736]));
  assign MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5751:5744]));
  assign MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_543_nl = (readslicef_29_22_7((MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_543_nl = nl_MultLoop_acc_543_nl[21:0];
  assign nl_MultLoop_acc_621_itm_1  = (MultLoop_acc_546_nl) + (MultLoop_acc_545_nl)
      + (MultLoop_acc_544_nl) + (MultLoop_acc_543_nl);
  assign nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5759:5752]));
  assign MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5767:5760]));
  assign MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_542_nl = (readslicef_29_22_7((MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_542_nl = nl_MultLoop_acc_542_nl[21:0];
  assign nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5775:5768]));
  assign MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5783:5776]));
  assign MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_541_nl = (readslicef_29_22_7((MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_541_nl = nl_MultLoop_acc_541_nl[21:0];
  assign nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5791:5784]));
  assign MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5799:5792]));
  assign MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_540_nl = (readslicef_29_22_7((MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_540_nl = nl_MultLoop_acc_540_nl[21:0];
  assign nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5807:5800]));
  assign MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5815:5808]));
  assign MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_539_nl = (readslicef_29_22_7((MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_539_nl = nl_MultLoop_acc_539_nl[21:0];
  assign nl_MultLoop_acc_620_itm_1  = (MultLoop_acc_542_nl) + (MultLoop_acc_541_nl)
      + (MultLoop_acc_540_nl) + (MultLoop_acc_539_nl);
  assign nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5823:5816]));
  assign MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5831:5824]));
  assign MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_538_nl = (readslicef_29_22_7((MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_538_nl = nl_MultLoop_acc_538_nl[21:0];
  assign nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5839:5832]));
  assign MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5847:5840]));
  assign MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_537_nl = (readslicef_29_22_7((MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_537_nl = nl_MultLoop_acc_537_nl[21:0];
  assign nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5855:5848]));
  assign MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5863:5856]));
  assign MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_536_nl = (readslicef_29_22_7((MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_536_nl = nl_MultLoop_acc_536_nl[21:0];
  assign nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5871:5864]));
  assign MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5879:5872]));
  assign MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_535_nl = (readslicef_29_22_7((MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_535_nl = nl_MultLoop_acc_535_nl[21:0];
  assign nl_MultLoop_acc_619_itm_1  = (MultLoop_acc_538_nl) + (MultLoop_acc_537_nl)
      + (MultLoop_acc_536_nl) + (MultLoop_acc_535_nl);
  assign nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5887:5880]));
  assign MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5895:5888]));
  assign MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_534_nl = (readslicef_29_22_7((MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_534_nl = nl_MultLoop_acc_534_nl[21:0];
  assign nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5903:5896]));
  assign MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5911:5904]));
  assign MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_533_nl = (readslicef_29_22_7((MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_533_nl = nl_MultLoop_acc_533_nl[21:0];
  assign nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5919:5912]));
  assign MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5927:5920]));
  assign MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_532_nl = (readslicef_29_22_7((MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_532_nl = nl_MultLoop_acc_532_nl[21:0];
  assign nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5935:5928]));
  assign MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5943:5936]));
  assign MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_531_nl = (readslicef_29_22_7((MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_531_nl = nl_MultLoop_acc_531_nl[21:0];
  assign nl_MultLoop_acc_618_itm_1  = (MultLoop_acc_534_nl) + (MultLoop_acc_533_nl)
      + (MultLoop_acc_532_nl) + (MultLoop_acc_531_nl);
  assign nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5951:5944]));
  assign MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5959:5952]));
  assign MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_530_nl = (readslicef_29_22_7((MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_530_nl = nl_MultLoop_acc_530_nl[21:0];
  assign nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5967:5960]));
  assign MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5975:5968]));
  assign MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_529_nl = (readslicef_29_22_7((MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_529_nl = nl_MultLoop_acc_529_nl[21:0];
  assign nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5983:5976]));
  assign MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5991:5984]));
  assign MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_528_nl = (readslicef_29_22_7((MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_528_nl = nl_MultLoop_acc_528_nl[21:0];
  assign nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5999:5992]));
  assign MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6007:6000]));
  assign MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_527_nl = (readslicef_29_22_7((MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_527_nl = nl_MultLoop_acc_527_nl[21:0];
  assign nl_MultLoop_acc_617_itm_1  = (MultLoop_acc_530_nl) + (MultLoop_acc_529_nl)
      + (MultLoop_acc_528_nl) + (MultLoop_acc_527_nl);
  assign nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6015:6008]));
  assign MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6023:6016]));
  assign MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_526_nl = (readslicef_29_22_7((MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_526_nl = nl_MultLoop_acc_526_nl[21:0];
  assign nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6031:6024]));
  assign MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6039:6032]));
  assign MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_525_nl = (readslicef_29_22_7((MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_525_nl = nl_MultLoop_acc_525_nl[21:0];
  assign nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6047:6040]));
  assign MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6055:6048]));
  assign MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_524_nl = (readslicef_29_22_7((MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_524_nl = nl_MultLoop_acc_524_nl[21:0];
  assign nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6063:6056]));
  assign MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6071:6064]));
  assign MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_523_nl = (readslicef_29_22_7((MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_523_nl = nl_MultLoop_acc_523_nl[21:0];
  assign nl_MultLoop_acc_616_itm_1  = (MultLoop_acc_526_nl) + (MultLoop_acc_525_nl)
      + (MultLoop_acc_524_nl) + (MultLoop_acc_523_nl);
  assign nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6079:6072]));
  assign MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6087:6080]));
  assign MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_522_nl = (readslicef_29_22_7((MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_522_nl = nl_MultLoop_acc_522_nl[21:0];
  assign nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6095:6088]));
  assign MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6103:6096]));
  assign MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_521_nl = (readslicef_29_22_7((MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_521_nl = nl_MultLoop_acc_521_nl[21:0];
  assign nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6111:6104]));
  assign MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6119:6112]));
  assign MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_520_nl = (readslicef_29_22_7((MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_520_nl = nl_MultLoop_acc_520_nl[21:0];
  assign nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6127:6120]));
  assign MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6135:6128]));
  assign MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_519_nl = (readslicef_29_22_7((MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_519_nl = nl_MultLoop_acc_519_nl[21:0];
  assign nl_MultLoop_acc_615_itm_1  = (MultLoop_acc_522_nl) + (MultLoop_acc_521_nl)
      + (MultLoop_acc_520_nl) + (MultLoop_acc_519_nl);
  assign nl_MultLoop_acc_1283_nl = (MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[39:32]);
  assign MultLoop_acc_1283_nl = nl_MultLoop_acc_1283_nl[10:0];
  assign nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[4103:4096]));
  assign MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_455_nl = ({(MultLoop_acc_1283_nl) , (MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_455_nl = nl_MultLoop_acc_455_nl[21:0];
  assign nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4111:4104]));
  assign MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4119:4112]));
  assign MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_454_nl = (readslicef_29_22_7((MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_454_nl = nl_MultLoop_acc_454_nl[21:0];
  assign nl_MultLoop_acc_487_nl = (MultLoop_acc_455_nl) + (MultLoop_acc_454_nl);
  assign MultLoop_acc_487_nl = nl_MultLoop_acc_487_nl[21:0];
  assign nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4127:4120]));
  assign MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4135:4128]));
  assign MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_453_nl = (readslicef_29_22_7((MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_453_nl = nl_MultLoop_acc_453_nl[21:0];
  assign nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4143:4136]));
  assign MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4151:4144]));
  assign MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_452_nl = (readslicef_29_22_7((MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_452_nl = nl_MultLoop_acc_452_nl[21:0];
  assign nl_MultLoop_acc_486_nl = (MultLoop_acc_453_nl) + (MultLoop_acc_452_nl);
  assign MultLoop_acc_486_nl = nl_MultLoop_acc_486_nl[21:0];
  assign nl_MultLoop_acc_503_itm_1  = (MultLoop_acc_487_nl) + (MultLoop_acc_486_nl);
  assign nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4159:4152]));
  assign MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4167:4160]));
  assign MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_451_nl = (readslicef_29_22_7((MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_451_nl = nl_MultLoop_acc_451_nl[21:0];
  assign nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4175:4168]));
  assign MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4183:4176]));
  assign MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_450_nl = (readslicef_29_22_7((MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_450_nl = nl_MultLoop_acc_450_nl[21:0];
  assign nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4191:4184]));
  assign MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4199:4192]));
  assign MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_449_nl = (readslicef_29_22_7((MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_449_nl = nl_MultLoop_acc_449_nl[21:0];
  assign nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4207:4200]));
  assign MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4215:4208]));
  assign MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_448_nl = (readslicef_29_22_7((MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_448_nl = nl_MultLoop_acc_448_nl[21:0];
  assign nl_MultLoop_acc_502_itm_1  = (MultLoop_acc_451_nl) + (MultLoop_acc_450_nl)
      + (MultLoop_acc_449_nl) + (MultLoop_acc_448_nl);
  assign nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4223:4216]));
  assign MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4231:4224]));
  assign MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_447_nl = (readslicef_29_22_7((MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_447_nl = nl_MultLoop_acc_447_nl[21:0];
  assign nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4239:4232]));
  assign MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4247:4240]));
  assign MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_446_nl = (readslicef_29_22_7((MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_446_nl = nl_MultLoop_acc_446_nl[21:0];
  assign nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4255:4248]));
  assign MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4263:4256]));
  assign MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_445_nl = (readslicef_29_22_7((MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_445_nl = nl_MultLoop_acc_445_nl[21:0];
  assign nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4271:4264]));
  assign MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4279:4272]));
  assign MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_444_nl = (readslicef_29_22_7((MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_444_nl = nl_MultLoop_acc_444_nl[21:0];
  assign nl_MultLoop_acc_501_itm_1  = (MultLoop_acc_447_nl) + (MultLoop_acc_446_nl)
      + (MultLoop_acc_445_nl) + (MultLoop_acc_444_nl);
  assign nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4287:4280]));
  assign MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4295:4288]));
  assign MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_443_nl = (readslicef_29_22_7((MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_443_nl = nl_MultLoop_acc_443_nl[21:0];
  assign nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4303:4296]));
  assign MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4311:4304]));
  assign MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_442_nl = (readslicef_29_22_7((MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_442_nl = nl_MultLoop_acc_442_nl[21:0];
  assign nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4319:4312]));
  assign MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4327:4320]));
  assign MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_441_nl = (readslicef_29_22_7((MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_441_nl = nl_MultLoop_acc_441_nl[21:0];
  assign nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4335:4328]));
  assign MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4343:4336]));
  assign MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_440_nl = (readslicef_29_22_7((MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_440_nl = nl_MultLoop_acc_440_nl[21:0];
  assign nl_MultLoop_acc_500_itm_1  = (MultLoop_acc_443_nl) + (MultLoop_acc_442_nl)
      + (MultLoop_acc_441_nl) + (MultLoop_acc_440_nl);
  assign nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4351:4344]));
  assign MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4359:4352]));
  assign MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_439_nl = (readslicef_29_22_7((MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_439_nl = nl_MultLoop_acc_439_nl[21:0];
  assign nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4367:4360]));
  assign MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4375:4368]));
  assign MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_438_nl = (readslicef_29_22_7((MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_438_nl = nl_MultLoop_acc_438_nl[21:0];
  assign nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4383:4376]));
  assign MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4391:4384]));
  assign MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_437_nl = (readslicef_29_22_7((MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_437_nl = nl_MultLoop_acc_437_nl[21:0];
  assign nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4399:4392]));
  assign MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4407:4400]));
  assign MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_436_nl = (readslicef_29_22_7((MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_436_nl = nl_MultLoop_acc_436_nl[21:0];
  assign nl_MultLoop_acc_499_itm_1  = (MultLoop_acc_439_nl) + (MultLoop_acc_438_nl)
      + (MultLoop_acc_437_nl) + (MultLoop_acc_436_nl);
  assign nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4415:4408]));
  assign MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4423:4416]));
  assign MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_435_nl = (readslicef_29_22_7((MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_435_nl = nl_MultLoop_acc_435_nl[21:0];
  assign nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4431:4424]));
  assign MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4439:4432]));
  assign MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_434_nl = (readslicef_29_22_7((MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_434_nl = nl_MultLoop_acc_434_nl[21:0];
  assign nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4447:4440]));
  assign MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4455:4448]));
  assign MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_433_nl = (readslicef_29_22_7((MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_433_nl = nl_MultLoop_acc_433_nl[21:0];
  assign nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4463:4456]));
  assign MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4471:4464]));
  assign MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_432_nl = (readslicef_29_22_7((MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_432_nl = nl_MultLoop_acc_432_nl[21:0];
  assign nl_MultLoop_acc_498_itm_1  = (MultLoop_acc_435_nl) + (MultLoop_acc_434_nl)
      + (MultLoop_acc_433_nl) + (MultLoop_acc_432_nl);
  assign nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4479:4472]));
  assign MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4487:4480]));
  assign MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_431_nl = (readslicef_29_22_7((MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_431_nl = nl_MultLoop_acc_431_nl[21:0];
  assign nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4495:4488]));
  assign MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4503:4496]));
  assign MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_430_nl = (readslicef_29_22_7((MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_430_nl = nl_MultLoop_acc_430_nl[21:0];
  assign nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4511:4504]));
  assign MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4519:4512]));
  assign MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_429_nl = (readslicef_29_22_7((MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_429_nl = nl_MultLoop_acc_429_nl[21:0];
  assign nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4527:4520]));
  assign MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4535:4528]));
  assign MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_428_nl = (readslicef_29_22_7((MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_428_nl = nl_MultLoop_acc_428_nl[21:0];
  assign nl_MultLoop_acc_497_itm_1  = (MultLoop_acc_431_nl) + (MultLoop_acc_430_nl)
      + (MultLoop_acc_429_nl) + (MultLoop_acc_428_nl);
  assign nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4543:4536]));
  assign MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4551:4544]));
  assign MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_427_nl = (readslicef_29_22_7((MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_427_nl = nl_MultLoop_acc_427_nl[21:0];
  assign nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4559:4552]));
  assign MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4567:4560]));
  assign MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_426_nl = (readslicef_29_22_7((MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_426_nl = nl_MultLoop_acc_426_nl[21:0];
  assign nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4575:4568]));
  assign MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4583:4576]));
  assign MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_425_nl = (readslicef_29_22_7((MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_425_nl = nl_MultLoop_acc_425_nl[21:0];
  assign nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4591:4584]));
  assign MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4599:4592]));
  assign MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_424_nl = (readslicef_29_22_7((MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_424_nl = nl_MultLoop_acc_424_nl[21:0];
  assign nl_MultLoop_acc_496_itm_1  = (MultLoop_acc_427_nl) + (MultLoop_acc_426_nl)
      + (MultLoop_acc_425_nl) + (MultLoop_acc_424_nl);
  assign nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4607:4600]));
  assign MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4615:4608]));
  assign MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_423_nl = (readslicef_29_22_7((MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_423_nl = nl_MultLoop_acc_423_nl[21:0];
  assign nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4623:4616]));
  assign MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4631:4624]));
  assign MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_422_nl = (readslicef_29_22_7((MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_422_nl = nl_MultLoop_acc_422_nl[21:0];
  assign nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4639:4632]));
  assign MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4647:4640]));
  assign MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_421_nl = (readslicef_29_22_7((MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_421_nl = nl_MultLoop_acc_421_nl[21:0];
  assign nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4655:4648]));
  assign MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4663:4656]));
  assign MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_420_nl = (readslicef_29_22_7((MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_420_nl = nl_MultLoop_acc_420_nl[21:0];
  assign nl_MultLoop_acc_495_itm_1  = (MultLoop_acc_423_nl) + (MultLoop_acc_422_nl)
      + (MultLoop_acc_421_nl) + (MultLoop_acc_420_nl);
  assign nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4671:4664]));
  assign MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4679:4672]));
  assign MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_419_nl = (readslicef_29_22_7((MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_419_nl = nl_MultLoop_acc_419_nl[21:0];
  assign nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4687:4680]));
  assign MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4695:4688]));
  assign MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_418_nl = (readslicef_29_22_7((MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_418_nl = nl_MultLoop_acc_418_nl[21:0];
  assign nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4703:4696]));
  assign MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4711:4704]));
  assign MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_417_nl = (readslicef_29_22_7((MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_417_nl = nl_MultLoop_acc_417_nl[21:0];
  assign nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4719:4712]));
  assign MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4727:4720]));
  assign MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_416_nl = (readslicef_29_22_7((MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_416_nl = nl_MultLoop_acc_416_nl[21:0];
  assign nl_MultLoop_acc_494_itm_1  = (MultLoop_acc_419_nl) + (MultLoop_acc_418_nl)
      + (MultLoop_acc_417_nl) + (MultLoop_acc_416_nl);
  assign nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4735:4728]));
  assign MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4743:4736]));
  assign MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_415_nl = (readslicef_29_22_7((MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_415_nl = nl_MultLoop_acc_415_nl[21:0];
  assign nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4751:4744]));
  assign MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4759:4752]));
  assign MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_414_nl = (readslicef_29_22_7((MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_414_nl = nl_MultLoop_acc_414_nl[21:0];
  assign nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4767:4760]));
  assign MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4775:4768]));
  assign MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_413_nl = (readslicef_29_22_7((MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_413_nl = nl_MultLoop_acc_413_nl[21:0];
  assign nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4783:4776]));
  assign MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4791:4784]));
  assign MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_412_nl = (readslicef_29_22_7((MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_412_nl = nl_MultLoop_acc_412_nl[21:0];
  assign nl_MultLoop_acc_493_itm_1  = (MultLoop_acc_415_nl) + (MultLoop_acc_414_nl)
      + (MultLoop_acc_413_nl) + (MultLoop_acc_412_nl);
  assign nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4799:4792]));
  assign MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4807:4800]));
  assign MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_411_nl = (readslicef_29_22_7((MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_411_nl = nl_MultLoop_acc_411_nl[21:0];
  assign nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4815:4808]));
  assign MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4823:4816]));
  assign MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_410_nl = (readslicef_29_22_7((MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_410_nl = nl_MultLoop_acc_410_nl[21:0];
  assign nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4831:4824]));
  assign MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4839:4832]));
  assign MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_409_nl = (readslicef_29_22_7((MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_409_nl = nl_MultLoop_acc_409_nl[21:0];
  assign nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4847:4840]));
  assign MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4855:4848]));
  assign MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_408_nl = (readslicef_29_22_7((MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_408_nl = nl_MultLoop_acc_408_nl[21:0];
  assign nl_MultLoop_acc_492_itm_1  = (MultLoop_acc_411_nl) + (MultLoop_acc_410_nl)
      + (MultLoop_acc_409_nl) + (MultLoop_acc_408_nl);
  assign nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4863:4856]));
  assign MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4871:4864]));
  assign MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_407_nl = (readslicef_29_22_7((MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_407_nl = nl_MultLoop_acc_407_nl[21:0];
  assign nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4879:4872]));
  assign MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4887:4880]));
  assign MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_406_nl = (readslicef_29_22_7((MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_406_nl = nl_MultLoop_acc_406_nl[21:0];
  assign nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4895:4888]));
  assign MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4903:4896]));
  assign MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_405_nl = (readslicef_29_22_7((MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_405_nl = nl_MultLoop_acc_405_nl[21:0];
  assign nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4911:4904]));
  assign MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4919:4912]));
  assign MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_404_nl = (readslicef_29_22_7((MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_404_nl = nl_MultLoop_acc_404_nl[21:0];
  assign nl_MultLoop_acc_491_itm_1  = (MultLoop_acc_407_nl) + (MultLoop_acc_406_nl)
      + (MultLoop_acc_405_nl) + (MultLoop_acc_404_nl);
  assign nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4927:4920]));
  assign MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4935:4928]));
  assign MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_403_nl = (readslicef_29_22_7((MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_403_nl = nl_MultLoop_acc_403_nl[21:0];
  assign nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4943:4936]));
  assign MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4951:4944]));
  assign MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_402_nl = (readslicef_29_22_7((MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_402_nl = nl_MultLoop_acc_402_nl[21:0];
  assign nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4959:4952]));
  assign MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4967:4960]));
  assign MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_401_nl = (readslicef_29_22_7((MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_401_nl = nl_MultLoop_acc_401_nl[21:0];
  assign nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4975:4968]));
  assign MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4983:4976]));
  assign MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_400_nl = (readslicef_29_22_7((MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_400_nl = nl_MultLoop_acc_400_nl[21:0];
  assign nl_MultLoop_acc_490_itm_1  = (MultLoop_acc_403_nl) + (MultLoop_acc_402_nl)
      + (MultLoop_acc_401_nl) + (MultLoop_acc_400_nl);
  assign nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4991:4984]));
  assign MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4999:4992]));
  assign MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_399_nl = (readslicef_29_22_7((MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_399_nl = nl_MultLoop_acc_399_nl[21:0];
  assign nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5007:5000]));
  assign MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5015:5008]));
  assign MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_398_nl = (readslicef_29_22_7((MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_398_nl = nl_MultLoop_acc_398_nl[21:0];
  assign nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5023:5016]));
  assign MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5031:5024]));
  assign MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_397_nl = (readslicef_29_22_7((MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_397_nl = nl_MultLoop_acc_397_nl[21:0];
  assign nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5039:5032]));
  assign MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5047:5040]));
  assign MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_396_nl = (readslicef_29_22_7((MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_396_nl = nl_MultLoop_acc_396_nl[21:0];
  assign nl_MultLoop_acc_489_itm_1  = (MultLoop_acc_399_nl) + (MultLoop_acc_398_nl)
      + (MultLoop_acc_397_nl) + (MultLoop_acc_396_nl);
  assign nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5055:5048]));
  assign MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5063:5056]));
  assign MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_395_nl = (readslicef_29_22_7((MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_395_nl = nl_MultLoop_acc_395_nl[21:0];
  assign nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5071:5064]));
  assign MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5079:5072]));
  assign MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_394_nl = (readslicef_29_22_7((MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_394_nl = nl_MultLoop_acc_394_nl[21:0];
  assign nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5087:5080]));
  assign MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5095:5088]));
  assign MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_393_nl = (readslicef_29_22_7((MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_393_nl = nl_MultLoop_acc_393_nl[21:0];
  assign nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5103:5096]));
  assign MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5111:5104]));
  assign MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_392_nl = (readslicef_29_22_7((MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_392_nl = nl_MultLoop_acc_392_nl[21:0];
  assign nl_MultLoop_acc_488_itm_1  = (MultLoop_acc_395_nl) + (MultLoop_acc_394_nl)
      + (MultLoop_acc_393_nl) + (MultLoop_acc_392_nl);
  assign nl_MultLoop_acc_1282_nl = (MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[31:24]);
  assign MultLoop_acc_1282_nl = nl_MultLoop_acc_1282_nl[10:0];
  assign nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[3079:3072]));
  assign MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_328_nl = ({(MultLoop_acc_1282_nl) , (MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_328_nl = nl_MultLoop_acc_328_nl[21:0];
  assign nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3087:3080]));
  assign MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3095:3088]));
  assign MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_327_nl = (readslicef_29_22_7((MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_327_nl = nl_MultLoop_acc_327_nl[21:0];
  assign nl_MultLoop_acc_360_nl = (MultLoop_acc_328_nl) + (MultLoop_acc_327_nl);
  assign MultLoop_acc_360_nl = nl_MultLoop_acc_360_nl[21:0];
  assign nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3103:3096]));
  assign MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3111:3104]));
  assign MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_326_nl = (readslicef_29_22_7((MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_326_nl = nl_MultLoop_acc_326_nl[21:0];
  assign nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3119:3112]));
  assign MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3127:3120]));
  assign MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_325_nl = (readslicef_29_22_7((MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_325_nl = nl_MultLoop_acc_325_nl[21:0];
  assign nl_MultLoop_acc_359_nl = (MultLoop_acc_326_nl) + (MultLoop_acc_325_nl);
  assign MultLoop_acc_359_nl = nl_MultLoop_acc_359_nl[21:0];
  assign nl_MultLoop_acc_376_itm_1  = (MultLoop_acc_360_nl) + (MultLoop_acc_359_nl);
  assign nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3135:3128]));
  assign MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3143:3136]));
  assign MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_324_nl = (readslicef_29_22_7((MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_324_nl = nl_MultLoop_acc_324_nl[21:0];
  assign nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3151:3144]));
  assign MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3159:3152]));
  assign MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_323_nl = (readslicef_29_22_7((MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_323_nl = nl_MultLoop_acc_323_nl[21:0];
  assign nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3167:3160]));
  assign MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3175:3168]));
  assign MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_322_nl = (readslicef_29_22_7((MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_322_nl = nl_MultLoop_acc_322_nl[21:0];
  assign nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3183:3176]));
  assign MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3191:3184]));
  assign MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_321_nl = (readslicef_29_22_7((MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_321_nl = nl_MultLoop_acc_321_nl[21:0];
  assign nl_MultLoop_acc_375_itm_1  = (MultLoop_acc_324_nl) + (MultLoop_acc_323_nl)
      + (MultLoop_acc_322_nl) + (MultLoop_acc_321_nl);
  assign nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3199:3192]));
  assign MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3207:3200]));
  assign MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_320_nl = (readslicef_29_22_7((MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_320_nl = nl_MultLoop_acc_320_nl[21:0];
  assign nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3215:3208]));
  assign MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3223:3216]));
  assign MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_319_nl = (readslicef_29_22_7((MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_319_nl = nl_MultLoop_acc_319_nl[21:0];
  assign nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3231:3224]));
  assign MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3239:3232]));
  assign MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_318_nl = (readslicef_29_22_7((MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_318_nl = nl_MultLoop_acc_318_nl[21:0];
  assign nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3247:3240]));
  assign MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3255:3248]));
  assign MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_317_nl = (readslicef_29_22_7((MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_317_nl = nl_MultLoop_acc_317_nl[21:0];
  assign nl_MultLoop_acc_374_itm_1  = (MultLoop_acc_320_nl) + (MultLoop_acc_319_nl)
      + (MultLoop_acc_318_nl) + (MultLoop_acc_317_nl);
  assign nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3263:3256]));
  assign MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3271:3264]));
  assign MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_316_nl = (readslicef_29_22_7((MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_316_nl = nl_MultLoop_acc_316_nl[21:0];
  assign nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3279:3272]));
  assign MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3287:3280]));
  assign MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_315_nl = (readslicef_29_22_7((MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_315_nl = nl_MultLoop_acc_315_nl[21:0];
  assign nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3295:3288]));
  assign MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3303:3296]));
  assign MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_314_nl = (readslicef_29_22_7((MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_314_nl = nl_MultLoop_acc_314_nl[21:0];
  assign nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3311:3304]));
  assign MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3319:3312]));
  assign MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_313_nl = (readslicef_29_22_7((MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_313_nl = nl_MultLoop_acc_313_nl[21:0];
  assign nl_MultLoop_acc_373_itm_1  = (MultLoop_acc_316_nl) + (MultLoop_acc_315_nl)
      + (MultLoop_acc_314_nl) + (MultLoop_acc_313_nl);
  assign nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3327:3320]));
  assign MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3335:3328]));
  assign MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_312_nl = (readslicef_29_22_7((MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_312_nl = nl_MultLoop_acc_312_nl[21:0];
  assign nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3343:3336]));
  assign MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3351:3344]));
  assign MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_311_nl = (readslicef_29_22_7((MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_311_nl = nl_MultLoop_acc_311_nl[21:0];
  assign nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3359:3352]));
  assign MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3367:3360]));
  assign MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_310_nl = (readslicef_29_22_7((MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[21:0];
  assign nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3375:3368]));
  assign MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3383:3376]));
  assign MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_309_nl = (readslicef_29_22_7((MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_309_nl = nl_MultLoop_acc_309_nl[21:0];
  assign nl_MultLoop_acc_372_itm_1  = (MultLoop_acc_312_nl) + (MultLoop_acc_311_nl)
      + (MultLoop_acc_310_nl) + (MultLoop_acc_309_nl);
  assign nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3391:3384]));
  assign MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3399:3392]));
  assign MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_308_nl = (readslicef_29_22_7((MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_308_nl = nl_MultLoop_acc_308_nl[21:0];
  assign nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3407:3400]));
  assign MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3415:3408]));
  assign MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_307_nl = (readslicef_29_22_7((MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[21:0];
  assign nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3423:3416]));
  assign MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3431:3424]));
  assign MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_306_nl = (readslicef_29_22_7((MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_306_nl = nl_MultLoop_acc_306_nl[21:0];
  assign nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3439:3432]));
  assign MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3447:3440]));
  assign MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_305_nl = (readslicef_29_22_7((MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_305_nl = nl_MultLoop_acc_305_nl[21:0];
  assign nl_MultLoop_acc_371_itm_1  = (MultLoop_acc_308_nl) + (MultLoop_acc_307_nl)
      + (MultLoop_acc_306_nl) + (MultLoop_acc_305_nl);
  assign nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3455:3448]));
  assign MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3463:3456]));
  assign MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_304_nl = (readslicef_29_22_7((MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[21:0];
  assign nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3471:3464]));
  assign MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3479:3472]));
  assign MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_303_nl = (readslicef_29_22_7((MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_303_nl = nl_MultLoop_acc_303_nl[21:0];
  assign nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3487:3480]));
  assign MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3495:3488]));
  assign MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_302_nl = (readslicef_29_22_7((MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_302_nl = nl_MultLoop_acc_302_nl[21:0];
  assign nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3503:3496]));
  assign MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3511:3504]));
  assign MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_301_nl = (readslicef_29_22_7((MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_301_nl = nl_MultLoop_acc_301_nl[21:0];
  assign nl_MultLoop_acc_370_itm_1  = (MultLoop_acc_304_nl) + (MultLoop_acc_303_nl)
      + (MultLoop_acc_302_nl) + (MultLoop_acc_301_nl);
  assign nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3519:3512]));
  assign MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3527:3520]));
  assign MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_300_nl = (readslicef_29_22_7((MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_300_nl = nl_MultLoop_acc_300_nl[21:0];
  assign nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3535:3528]));
  assign MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3543:3536]));
  assign MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_299_nl = (readslicef_29_22_7((MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_299_nl = nl_MultLoop_acc_299_nl[21:0];
  assign nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3551:3544]));
  assign MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3559:3552]));
  assign MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_298_nl = (readslicef_29_22_7((MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_298_nl = nl_MultLoop_acc_298_nl[21:0];
  assign nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3567:3560]));
  assign MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3575:3568]));
  assign MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_297_nl = (readslicef_29_22_7((MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_297_nl = nl_MultLoop_acc_297_nl[21:0];
  assign nl_MultLoop_acc_369_itm_1  = (MultLoop_acc_300_nl) + (MultLoop_acc_299_nl)
      + (MultLoop_acc_298_nl) + (MultLoop_acc_297_nl);
  assign nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3583:3576]));
  assign MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3591:3584]));
  assign MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_296_nl = (readslicef_29_22_7((MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_296_nl = nl_MultLoop_acc_296_nl[21:0];
  assign nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3599:3592]));
  assign MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3607:3600]));
  assign MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_295_nl = (readslicef_29_22_7((MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_295_nl = nl_MultLoop_acc_295_nl[21:0];
  assign nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3615:3608]));
  assign MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3623:3616]));
  assign MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_294_nl = (readslicef_29_22_7((MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_294_nl = nl_MultLoop_acc_294_nl[21:0];
  assign nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3631:3624]));
  assign MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3639:3632]));
  assign MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_293_nl = (readslicef_29_22_7((MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_293_nl = nl_MultLoop_acc_293_nl[21:0];
  assign nl_MultLoop_acc_368_itm_1  = (MultLoop_acc_296_nl) + (MultLoop_acc_295_nl)
      + (MultLoop_acc_294_nl) + (MultLoop_acc_293_nl);
  assign nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3647:3640]));
  assign MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3655:3648]));
  assign MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_292_nl = (readslicef_29_22_7((MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_292_nl = nl_MultLoop_acc_292_nl[21:0];
  assign nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3663:3656]));
  assign MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3671:3664]));
  assign MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_291_nl = (readslicef_29_22_7((MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_291_nl = nl_MultLoop_acc_291_nl[21:0];
  assign nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3679:3672]));
  assign MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3687:3680]));
  assign MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_290_nl = (readslicef_29_22_7((MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_290_nl = nl_MultLoop_acc_290_nl[21:0];
  assign nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3695:3688]));
  assign MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3703:3696]));
  assign MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_289_nl = (readslicef_29_22_7((MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_289_nl = nl_MultLoop_acc_289_nl[21:0];
  assign nl_MultLoop_acc_367_itm_1  = (MultLoop_acc_292_nl) + (MultLoop_acc_291_nl)
      + (MultLoop_acc_290_nl) + (MultLoop_acc_289_nl);
  assign nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3711:3704]));
  assign MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3719:3712]));
  assign MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_288_nl = (readslicef_29_22_7((MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_288_nl = nl_MultLoop_acc_288_nl[21:0];
  assign nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3727:3720]));
  assign MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3735:3728]));
  assign MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_287_nl = (readslicef_29_22_7((MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_287_nl = nl_MultLoop_acc_287_nl[21:0];
  assign nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3743:3736]));
  assign MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3751:3744]));
  assign MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_286_nl = (readslicef_29_22_7((MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_286_nl = nl_MultLoop_acc_286_nl[21:0];
  assign nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3759:3752]));
  assign MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3767:3760]));
  assign MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_285_nl = (readslicef_29_22_7((MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_285_nl = nl_MultLoop_acc_285_nl[21:0];
  assign nl_MultLoop_acc_366_itm_1  = (MultLoop_acc_288_nl) + (MultLoop_acc_287_nl)
      + (MultLoop_acc_286_nl) + (MultLoop_acc_285_nl);
  assign nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3775:3768]));
  assign MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3783:3776]));
  assign MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_284_nl = (readslicef_29_22_7((MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_284_nl = nl_MultLoop_acc_284_nl[21:0];
  assign nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3791:3784]));
  assign MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3799:3792]));
  assign MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_283_nl = (readslicef_29_22_7((MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_283_nl = nl_MultLoop_acc_283_nl[21:0];
  assign nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3807:3800]));
  assign MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3815:3808]));
  assign MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_282_nl = (readslicef_29_22_7((MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_282_nl = nl_MultLoop_acc_282_nl[21:0];
  assign nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3823:3816]));
  assign MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3831:3824]));
  assign MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_281_nl = (readslicef_29_22_7((MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_281_nl = nl_MultLoop_acc_281_nl[21:0];
  assign nl_MultLoop_acc_365_itm_1  = (MultLoop_acc_284_nl) + (MultLoop_acc_283_nl)
      + (MultLoop_acc_282_nl) + (MultLoop_acc_281_nl);
  assign nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3839:3832]));
  assign MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3847:3840]));
  assign MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_280_nl = (readslicef_29_22_7((MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_280_nl = nl_MultLoop_acc_280_nl[21:0];
  assign nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3855:3848]));
  assign MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3863:3856]));
  assign MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_279_nl = (readslicef_29_22_7((MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_279_nl = nl_MultLoop_acc_279_nl[21:0];
  assign nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3871:3864]));
  assign MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3879:3872]));
  assign MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_278_nl = (readslicef_29_22_7((MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_278_nl = nl_MultLoop_acc_278_nl[21:0];
  assign nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3887:3880]));
  assign MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3895:3888]));
  assign MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_277_nl = (readslicef_29_22_7((MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_277_nl = nl_MultLoop_acc_277_nl[21:0];
  assign nl_MultLoop_acc_364_itm_1  = (MultLoop_acc_280_nl) + (MultLoop_acc_279_nl)
      + (MultLoop_acc_278_nl) + (MultLoop_acc_277_nl);
  assign nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3903:3896]));
  assign MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3911:3904]));
  assign MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_276_nl = (readslicef_29_22_7((MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_276_nl = nl_MultLoop_acc_276_nl[21:0];
  assign nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3919:3912]));
  assign MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3927:3920]));
  assign MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_275_nl = (readslicef_29_22_7((MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_275_nl = nl_MultLoop_acc_275_nl[21:0];
  assign nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3935:3928]));
  assign MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3943:3936]));
  assign MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_274_nl = (readslicef_29_22_7((MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_274_nl = nl_MultLoop_acc_274_nl[21:0];
  assign nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3951:3944]));
  assign MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3959:3952]));
  assign MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_273_nl = (readslicef_29_22_7((MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_273_nl = nl_MultLoop_acc_273_nl[21:0];
  assign nl_MultLoop_acc_363_itm_1  = (MultLoop_acc_276_nl) + (MultLoop_acc_275_nl)
      + (MultLoop_acc_274_nl) + (MultLoop_acc_273_nl);
  assign nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3967:3960]));
  assign MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3975:3968]));
  assign MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_272_nl = (readslicef_29_22_7((MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_272_nl = nl_MultLoop_acc_272_nl[21:0];
  assign nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3983:3976]));
  assign MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3991:3984]));
  assign MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_271_nl = (readslicef_29_22_7((MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[21:0];
  assign nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3999:3992]));
  assign MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4007:4000]));
  assign MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_270_nl = (readslicef_29_22_7((MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[21:0];
  assign nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4015:4008]));
  assign MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4023:4016]));
  assign MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_269_nl = (readslicef_29_22_7((MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_269_nl = nl_MultLoop_acc_269_nl[21:0];
  assign nl_MultLoop_acc_362_itm_1  = (MultLoop_acc_272_nl) + (MultLoop_acc_271_nl)
      + (MultLoop_acc_270_nl) + (MultLoop_acc_269_nl);
  assign nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4031:4024]));
  assign MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4039:4032]));
  assign MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_268_nl = (readslicef_29_22_7((MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_268_nl = nl_MultLoop_acc_268_nl[21:0];
  assign nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4047:4040]));
  assign MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4055:4048]));
  assign MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_267_nl = (readslicef_29_22_7((MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_267_nl = nl_MultLoop_acc_267_nl[21:0];
  assign nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4063:4056]));
  assign MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4071:4064]));
  assign MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_266_nl = (readslicef_29_22_7((MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_266_nl = nl_MultLoop_acc_266_nl[21:0];
  assign nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4079:4072]));
  assign MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4087:4080]));
  assign MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_265_nl = (readslicef_29_22_7((MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_265_nl = nl_MultLoop_acc_265_nl[21:0];
  assign nl_MultLoop_acc_361_itm_1  = (MultLoop_acc_268_nl) + (MultLoop_acc_267_nl)
      + (MultLoop_acc_266_nl) + (MultLoop_acc_265_nl);
  assign nl_MultLoop_acc_1281_nl = (MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[23:16]);
  assign MultLoop_acc_1281_nl = nl_MultLoop_acc_1281_nl[10:0];
  assign nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[2055:2048]));
  assign MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_201_nl = ({(MultLoop_acc_1281_nl) , (MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_201_nl = nl_MultLoop_acc_201_nl[21:0];
  assign nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2063:2056]));
  assign MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2071:2064]));
  assign MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_200_nl = (readslicef_29_22_7((MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_200_nl = nl_MultLoop_acc_200_nl[21:0];
  assign nl_MultLoop_acc_233_nl = (MultLoop_acc_201_nl) + (MultLoop_acc_200_nl);
  assign MultLoop_acc_233_nl = nl_MultLoop_acc_233_nl[21:0];
  assign nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2079:2072]));
  assign MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2087:2080]));
  assign MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_199_nl = (readslicef_29_22_7((MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_199_nl = nl_MultLoop_acc_199_nl[21:0];
  assign nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2095:2088]));
  assign MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2103:2096]));
  assign MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_198_nl = (readslicef_29_22_7((MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_198_nl = nl_MultLoop_acc_198_nl[21:0];
  assign nl_MultLoop_acc_232_nl = (MultLoop_acc_199_nl) + (MultLoop_acc_198_nl);
  assign MultLoop_acc_232_nl = nl_MultLoop_acc_232_nl[21:0];
  assign nl_MultLoop_acc_249_itm_1  = (MultLoop_acc_233_nl) + (MultLoop_acc_232_nl);
  assign nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2111:2104]));
  assign MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2119:2112]));
  assign MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_197_nl = (readslicef_29_22_7((MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_197_nl = nl_MultLoop_acc_197_nl[21:0];
  assign nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2127:2120]));
  assign MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2135:2128]));
  assign MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_196_nl = (readslicef_29_22_7((MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_196_nl = nl_MultLoop_acc_196_nl[21:0];
  assign nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2143:2136]));
  assign MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2151:2144]));
  assign MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_195_nl = (readslicef_29_22_7((MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_195_nl = nl_MultLoop_acc_195_nl[21:0];
  assign nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2159:2152]));
  assign MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2167:2160]));
  assign MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_194_nl = (readslicef_29_22_7((MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_194_nl = nl_MultLoop_acc_194_nl[21:0];
  assign nl_MultLoop_acc_248_itm_1  = (MultLoop_acc_197_nl) + (MultLoop_acc_196_nl)
      + (MultLoop_acc_195_nl) + (MultLoop_acc_194_nl);
  assign nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2175:2168]));
  assign MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2183:2176]));
  assign MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_193_nl = (readslicef_29_22_7((MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_193_nl = nl_MultLoop_acc_193_nl[21:0];
  assign nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2191:2184]));
  assign MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2199:2192]));
  assign MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_192_nl = (readslicef_29_22_7((MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_192_nl = nl_MultLoop_acc_192_nl[21:0];
  assign nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2207:2200]));
  assign MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2215:2208]));
  assign MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_191_nl = (readslicef_29_22_7((MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_191_nl = nl_MultLoop_acc_191_nl[21:0];
  assign nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2223:2216]));
  assign MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2231:2224]));
  assign MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_190_nl = (readslicef_29_22_7((MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_190_nl = nl_MultLoop_acc_190_nl[21:0];
  assign nl_MultLoop_acc_247_itm_1  = (MultLoop_acc_193_nl) + (MultLoop_acc_192_nl)
      + (MultLoop_acc_191_nl) + (MultLoop_acc_190_nl);
  assign nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2239:2232]));
  assign MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2247:2240]));
  assign MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_189_nl = (readslicef_29_22_7((MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_189_nl = nl_MultLoop_acc_189_nl[21:0];
  assign nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2255:2248]));
  assign MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2263:2256]));
  assign MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_188_nl = (readslicef_29_22_7((MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_188_nl = nl_MultLoop_acc_188_nl[21:0];
  assign nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2271:2264]));
  assign MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2279:2272]));
  assign MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_187_nl = (readslicef_29_22_7((MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_187_nl = nl_MultLoop_acc_187_nl[21:0];
  assign nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2287:2280]));
  assign MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2295:2288]));
  assign MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_186_nl = (readslicef_29_22_7((MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_186_nl = nl_MultLoop_acc_186_nl[21:0];
  assign nl_MultLoop_acc_246_itm_1  = (MultLoop_acc_189_nl) + (MultLoop_acc_188_nl)
      + (MultLoop_acc_187_nl) + (MultLoop_acc_186_nl);
  assign nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2303:2296]));
  assign MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2311:2304]));
  assign MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_185_nl = (readslicef_29_22_7((MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_185_nl = nl_MultLoop_acc_185_nl[21:0];
  assign nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2319:2312]));
  assign MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2327:2320]));
  assign MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_184_nl = (readslicef_29_22_7((MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_184_nl = nl_MultLoop_acc_184_nl[21:0];
  assign nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2335:2328]));
  assign MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2343:2336]));
  assign MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_183_nl = (readslicef_29_22_7((MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_183_nl = nl_MultLoop_acc_183_nl[21:0];
  assign nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2351:2344]));
  assign MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2359:2352]));
  assign MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_182_nl = (readslicef_29_22_7((MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_182_nl = nl_MultLoop_acc_182_nl[21:0];
  assign nl_MultLoop_acc_245_itm_1  = (MultLoop_acc_185_nl) + (MultLoop_acc_184_nl)
      + (MultLoop_acc_183_nl) + (MultLoop_acc_182_nl);
  assign nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2367:2360]));
  assign MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2375:2368]));
  assign MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_181_nl = (readslicef_29_22_7((MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_181_nl = nl_MultLoop_acc_181_nl[21:0];
  assign nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2383:2376]));
  assign MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2391:2384]));
  assign MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_180_nl = (readslicef_29_22_7((MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_180_nl = nl_MultLoop_acc_180_nl[21:0];
  assign nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2399:2392]));
  assign MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2407:2400]));
  assign MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_179_nl = (readslicef_29_22_7((MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_179_nl = nl_MultLoop_acc_179_nl[21:0];
  assign nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2415:2408]));
  assign MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2423:2416]));
  assign MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_178_nl = (readslicef_29_22_7((MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_178_nl = nl_MultLoop_acc_178_nl[21:0];
  assign nl_MultLoop_acc_244_itm_1  = (MultLoop_acc_181_nl) + (MultLoop_acc_180_nl)
      + (MultLoop_acc_179_nl) + (MultLoop_acc_178_nl);
  assign nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2431:2424]));
  assign MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2439:2432]));
  assign MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_177_nl = (readslicef_29_22_7((MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_177_nl = nl_MultLoop_acc_177_nl[21:0];
  assign nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2447:2440]));
  assign MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2455:2448]));
  assign MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_176_nl = (readslicef_29_22_7((MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_176_nl = nl_MultLoop_acc_176_nl[21:0];
  assign nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2463:2456]));
  assign MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2471:2464]));
  assign MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_175_nl = (readslicef_29_22_7((MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_175_nl = nl_MultLoop_acc_175_nl[21:0];
  assign nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2479:2472]));
  assign MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2487:2480]));
  assign MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_174_nl = (readslicef_29_22_7((MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_174_nl = nl_MultLoop_acc_174_nl[21:0];
  assign nl_MultLoop_acc_243_itm_1  = (MultLoop_acc_177_nl) + (MultLoop_acc_176_nl)
      + (MultLoop_acc_175_nl) + (MultLoop_acc_174_nl);
  assign nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2495:2488]));
  assign MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2503:2496]));
  assign MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_173_nl = (readslicef_29_22_7((MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_173_nl = nl_MultLoop_acc_173_nl[21:0];
  assign nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2511:2504]));
  assign MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2519:2512]));
  assign MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_172_nl = (readslicef_29_22_7((MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_172_nl = nl_MultLoop_acc_172_nl[21:0];
  assign nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2527:2520]));
  assign MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2535:2528]));
  assign MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_171_nl = (readslicef_29_22_7((MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_171_nl = nl_MultLoop_acc_171_nl[21:0];
  assign nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2543:2536]));
  assign MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2551:2544]));
  assign MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_170_nl = (readslicef_29_22_7((MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_170_nl = nl_MultLoop_acc_170_nl[21:0];
  assign nl_MultLoop_acc_242_itm_1  = (MultLoop_acc_173_nl) + (MultLoop_acc_172_nl)
      + (MultLoop_acc_171_nl) + (MultLoop_acc_170_nl);
  assign nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2559:2552]));
  assign MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2567:2560]));
  assign MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_169_nl = (readslicef_29_22_7((MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_169_nl = nl_MultLoop_acc_169_nl[21:0];
  assign nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2575:2568]));
  assign MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2583:2576]));
  assign MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_168_nl = (readslicef_29_22_7((MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_168_nl = nl_MultLoop_acc_168_nl[21:0];
  assign nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2591:2584]));
  assign MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2599:2592]));
  assign MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_167_nl = (readslicef_29_22_7((MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_167_nl = nl_MultLoop_acc_167_nl[21:0];
  assign nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2607:2600]));
  assign MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2615:2608]));
  assign MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_166_nl = (readslicef_29_22_7((MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_166_nl = nl_MultLoop_acc_166_nl[21:0];
  assign nl_MultLoop_acc_241_itm_1  = (MultLoop_acc_169_nl) + (MultLoop_acc_168_nl)
      + (MultLoop_acc_167_nl) + (MultLoop_acc_166_nl);
  assign nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2623:2616]));
  assign MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2631:2624]));
  assign MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_165_nl = (readslicef_29_22_7((MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[21:0];
  assign nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2639:2632]));
  assign MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2647:2640]));
  assign MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_164_nl = (readslicef_29_22_7((MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_164_nl = nl_MultLoop_acc_164_nl[21:0];
  assign nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2655:2648]));
  assign MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2663:2656]));
  assign MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_163_nl = (readslicef_29_22_7((MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_163_nl = nl_MultLoop_acc_163_nl[21:0];
  assign nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2671:2664]));
  assign MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2679:2672]));
  assign MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_162_nl = (readslicef_29_22_7((MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_162_nl = nl_MultLoop_acc_162_nl[21:0];
  assign nl_MultLoop_acc_240_itm_1  = (MultLoop_acc_165_nl) + (MultLoop_acc_164_nl)
      + (MultLoop_acc_163_nl) + (MultLoop_acc_162_nl);
  assign nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2687:2680]));
  assign MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2695:2688]));
  assign MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_161_nl = (readslicef_29_22_7((MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_161_nl = nl_MultLoop_acc_161_nl[21:0];
  assign nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2703:2696]));
  assign MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2711:2704]));
  assign MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_160_nl = (readslicef_29_22_7((MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_160_nl = nl_MultLoop_acc_160_nl[21:0];
  assign nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2719:2712]));
  assign MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2727:2720]));
  assign MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_159_nl = (readslicef_29_22_7((MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[21:0];
  assign nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2735:2728]));
  assign MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2743:2736]));
  assign MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_158_nl = (readslicef_29_22_7((MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[21:0];
  assign nl_MultLoop_acc_239_itm_1  = (MultLoop_acc_161_nl) + (MultLoop_acc_160_nl)
      + (MultLoop_acc_159_nl) + (MultLoop_acc_158_nl);
  assign nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2751:2744]));
  assign MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2759:2752]));
  assign MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_157_nl = (readslicef_29_22_7((MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_157_nl = nl_MultLoop_acc_157_nl[21:0];
  assign nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2767:2760]));
  assign MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2775:2768]));
  assign MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_156_nl = (readslicef_29_22_7((MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_156_nl = nl_MultLoop_acc_156_nl[21:0];
  assign nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2783:2776]));
  assign MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2791:2784]));
  assign MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_155_nl = (readslicef_29_22_7((MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_155_nl = nl_MultLoop_acc_155_nl[21:0];
  assign nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2799:2792]));
  assign MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2807:2800]));
  assign MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_154_nl = (readslicef_29_22_7((MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_154_nl = nl_MultLoop_acc_154_nl[21:0];
  assign nl_MultLoop_acc_238_itm_1  = (MultLoop_acc_157_nl) + (MultLoop_acc_156_nl)
      + (MultLoop_acc_155_nl) + (MultLoop_acc_154_nl);
  assign nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2815:2808]));
  assign MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2823:2816]));
  assign MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_153_nl = (readslicef_29_22_7((MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_153_nl = nl_MultLoop_acc_153_nl[21:0];
  assign nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2831:2824]));
  assign MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2839:2832]));
  assign MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_152_nl = (readslicef_29_22_7((MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_152_nl = nl_MultLoop_acc_152_nl[21:0];
  assign nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2847:2840]));
  assign MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2855:2848]));
  assign MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_151_nl = (readslicef_29_22_7((MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_151_nl = nl_MultLoop_acc_151_nl[21:0];
  assign nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2863:2856]));
  assign MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2871:2864]));
  assign MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_150_nl = (readslicef_29_22_7((MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_150_nl = nl_MultLoop_acc_150_nl[21:0];
  assign nl_MultLoop_acc_237_itm_1  = (MultLoop_acc_153_nl) + (MultLoop_acc_152_nl)
      + (MultLoop_acc_151_nl) + (MultLoop_acc_150_nl);
  assign nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2879:2872]));
  assign MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2887:2880]));
  assign MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_149_nl = (readslicef_29_22_7((MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_149_nl = nl_MultLoop_acc_149_nl[21:0];
  assign nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2895:2888]));
  assign MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2903:2896]));
  assign MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_148_nl = (readslicef_29_22_7((MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_148_nl = nl_MultLoop_acc_148_nl[21:0];
  assign nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2911:2904]));
  assign MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2919:2912]));
  assign MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_147_nl = (readslicef_29_22_7((MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_147_nl = nl_MultLoop_acc_147_nl[21:0];
  assign nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2927:2920]));
  assign MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2935:2928]));
  assign MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_146_nl = (readslicef_29_22_7((MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_146_nl = nl_MultLoop_acc_146_nl[21:0];
  assign nl_MultLoop_acc_236_itm_1  = (MultLoop_acc_149_nl) + (MultLoop_acc_148_nl)
      + (MultLoop_acc_147_nl) + (MultLoop_acc_146_nl);
  assign nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2943:2936]));
  assign MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2951:2944]));
  assign MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_145_nl = (readslicef_29_22_7((MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_145_nl = nl_MultLoop_acc_145_nl[21:0];
  assign nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2959:2952]));
  assign MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2967:2960]));
  assign MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_144_nl = (readslicef_29_22_7((MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_144_nl = nl_MultLoop_acc_144_nl[21:0];
  assign nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2975:2968]));
  assign MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2983:2976]));
  assign MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_143_nl = (readslicef_29_22_7((MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[21:0];
  assign nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2991:2984]));
  assign MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2999:2992]));
  assign MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_142_nl = (readslicef_29_22_7((MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_142_nl = nl_MultLoop_acc_142_nl[21:0];
  assign nl_MultLoop_acc_235_itm_1  = (MultLoop_acc_145_nl) + (MultLoop_acc_144_nl)
      + (MultLoop_acc_143_nl) + (MultLoop_acc_142_nl);
  assign nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3007:3000]));
  assign MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3015:3008]));
  assign MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_141_nl = (readslicef_29_22_7((MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_141_nl = nl_MultLoop_acc_141_nl[21:0];
  assign nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3023:3016]));
  assign MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3031:3024]));
  assign MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_140_nl = (readslicef_29_22_7((MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_140_nl = nl_MultLoop_acc_140_nl[21:0];
  assign nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3039:3032]));
  assign MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3047:3040]));
  assign MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_139_nl = (readslicef_29_22_7((MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_139_nl = nl_MultLoop_acc_139_nl[21:0];
  assign nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3055:3048]));
  assign MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3063:3056]));
  assign MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_138_nl = (readslicef_29_22_7((MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_138_nl = nl_MultLoop_acc_138_nl[21:0];
  assign nl_MultLoop_acc_234_itm_1  = (MultLoop_acc_141_nl) + (MultLoop_acc_140_nl)
      + (MultLoop_acc_139_nl) + (MultLoop_acc_138_nl);
  assign nl_MultLoop_acc_1280_nl = (MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2s_8_11(b4_rsci_idat_mxwt[15:8]);
  assign MultLoop_acc_1280_nl = nl_MultLoop_acc_1280_nl[10:0];
  assign nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[1031:1024]));
  assign MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_106_nl = ({(MultLoop_acc_1280_nl) , (MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_106_nl = nl_MultLoop_acc_106_nl[21:0];
  assign nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1039:1032]));
  assign MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1047:1040]));
  assign MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_73_nl = (readslicef_29_22_7((MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[21:0];
  assign nl_MultLoop_acc_122_nl = (MultLoop_acc_106_nl) + (MultLoop_acc_73_nl);
  assign MultLoop_acc_122_nl = nl_MultLoop_acc_122_nl[21:0];
  assign nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1055:1048]));
  assign MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1063:1056]));
  assign MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_72_nl = (readslicef_29_22_7((MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_72_nl = nl_MultLoop_acc_72_nl[21:0];
  assign nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1071:1064]));
  assign MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1079:1072]));
  assign MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_71_nl = (readslicef_29_22_7((MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_71_nl = nl_MultLoop_acc_71_nl[21:0];
  assign nl_MultLoop_acc_105_nl = (MultLoop_acc_72_nl) + (MultLoop_acc_71_nl);
  assign MultLoop_acc_105_nl = nl_MultLoop_acc_105_nl[21:0];
  assign nl_MultLoop_acc_130_itm_1  = (MultLoop_acc_122_nl) + (MultLoop_acc_105_nl);
  assign nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1087:1080]));
  assign MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1095:1088]));
  assign MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_70_nl = (readslicef_29_22_7((MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_70_nl = nl_MultLoop_acc_70_nl[21:0];
  assign nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1103:1096]));
  assign MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1111:1104]));
  assign MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_69_nl = (readslicef_29_22_7((MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_69_nl = nl_MultLoop_acc_69_nl[21:0];
  assign nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1119:1112]));
  assign MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1127:1120]));
  assign MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_68_nl = (readslicef_29_22_7((MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_68_nl = nl_MultLoop_acc_68_nl[21:0];
  assign nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1135:1128]));
  assign MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1143:1136]));
  assign MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_67_nl = (readslicef_29_22_7((MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_67_nl = nl_MultLoop_acc_67_nl[21:0];
  assign nl_MultLoop_acc_121_itm_1  = (MultLoop_acc_70_nl) + (MultLoop_acc_69_nl)
      + (MultLoop_acc_68_nl) + (MultLoop_acc_67_nl);
  assign nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1151:1144]));
  assign MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1159:1152]));
  assign MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_66_nl = (readslicef_29_22_7((MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_66_nl = nl_MultLoop_acc_66_nl[21:0];
  assign nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1167:1160]));
  assign MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1175:1168]));
  assign MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_65_nl = (readslicef_29_22_7((MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[21:0];
  assign nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1183:1176]));
  assign MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1191:1184]));
  assign MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_64_nl = (readslicef_29_22_7((MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_64_nl = nl_MultLoop_acc_64_nl[21:0];
  assign nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1199:1192]));
  assign MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1207:1200]));
  assign MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_63_nl = (readslicef_29_22_7((MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_63_nl = nl_MultLoop_acc_63_nl[21:0];
  assign nl_MultLoop_acc_120_itm_1  = (MultLoop_acc_66_nl) + (MultLoop_acc_65_nl)
      + (MultLoop_acc_64_nl) + (MultLoop_acc_63_nl);
  assign nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1215:1208]));
  assign MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1223:1216]));
  assign MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_62_nl = (readslicef_29_22_7((MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_62_nl = nl_MultLoop_acc_62_nl[21:0];
  assign nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1231:1224]));
  assign MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1239:1232]));
  assign MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_61_nl = (readslicef_29_22_7((MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_61_nl = nl_MultLoop_acc_61_nl[21:0];
  assign nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1247:1240]));
  assign MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1255:1248]));
  assign MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_60_nl = (readslicef_29_22_7((MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_60_nl = nl_MultLoop_acc_60_nl[21:0];
  assign nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1263:1256]));
  assign MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1271:1264]));
  assign MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_59_nl = (readslicef_29_22_7((MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_59_nl = nl_MultLoop_acc_59_nl[21:0];
  assign nl_MultLoop_acc_119_itm_1  = (MultLoop_acc_62_nl) + (MultLoop_acc_61_nl)
      + (MultLoop_acc_60_nl) + (MultLoop_acc_59_nl);
  assign nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1279:1272]));
  assign MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1287:1280]));
  assign MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_58_nl = (readslicef_29_22_7((MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_58_nl = nl_MultLoop_acc_58_nl[21:0];
  assign nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1295:1288]));
  assign MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1303:1296]));
  assign MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_57_nl = (readslicef_29_22_7((MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_57_nl = nl_MultLoop_acc_57_nl[21:0];
  assign nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1311:1304]));
  assign MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1319:1312]));
  assign MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_56_nl = (readslicef_29_22_7((MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_56_nl = nl_MultLoop_acc_56_nl[21:0];
  assign nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1327:1320]));
  assign MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1335:1328]));
  assign MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_55_nl = (readslicef_29_22_7((MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_55_nl = nl_MultLoop_acc_55_nl[21:0];
  assign nl_MultLoop_acc_118_itm_1  = (MultLoop_acc_58_nl) + (MultLoop_acc_57_nl)
      + (MultLoop_acc_56_nl) + (MultLoop_acc_55_nl);
  assign nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1343:1336]));
  assign MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1351:1344]));
  assign MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_54_nl = (readslicef_29_22_7((MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_54_nl = nl_MultLoop_acc_54_nl[21:0];
  assign nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1359:1352]));
  assign MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1367:1360]));
  assign MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_53_nl = (readslicef_29_22_7((MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[21:0];
  assign nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1375:1368]));
  assign MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1383:1376]));
  assign MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_52_nl = (readslicef_29_22_7((MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_52_nl = nl_MultLoop_acc_52_nl[21:0];
  assign nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1391:1384]));
  assign MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1399:1392]));
  assign MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_51_nl = (readslicef_29_22_7((MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_51_nl = nl_MultLoop_acc_51_nl[21:0];
  assign nl_MultLoop_acc_117_itm_1  = (MultLoop_acc_54_nl) + (MultLoop_acc_53_nl)
      + (MultLoop_acc_52_nl) + (MultLoop_acc_51_nl);
  assign nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1407:1400]));
  assign MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1415:1408]));
  assign MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_50_nl = (readslicef_29_22_7((MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_50_nl = nl_MultLoop_acc_50_nl[21:0];
  assign nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1423:1416]));
  assign MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1431:1424]));
  assign MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_49_nl = (readslicef_29_22_7((MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_49_nl = nl_MultLoop_acc_49_nl[21:0];
  assign nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1439:1432]));
  assign MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1447:1440]));
  assign MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_48_nl = (readslicef_29_22_7((MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_48_nl = nl_MultLoop_acc_48_nl[21:0];
  assign nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1455:1448]));
  assign MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1463:1456]));
  assign MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_47_nl = (readslicef_29_22_7((MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_47_nl = nl_MultLoop_acc_47_nl[21:0];
  assign nl_MultLoop_acc_116_itm_1  = (MultLoop_acc_50_nl) + (MultLoop_acc_49_nl)
      + (MultLoop_acc_48_nl) + (MultLoop_acc_47_nl);
  assign nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1471:1464]));
  assign MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1479:1472]));
  assign MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_46_nl = (readslicef_29_22_7((MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_46_nl = nl_MultLoop_acc_46_nl[21:0];
  assign nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1487:1480]));
  assign MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1495:1488]));
  assign MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_45_nl = (readslicef_29_22_7((MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[21:0];
  assign nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1503:1496]));
  assign MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1511:1504]));
  assign MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_44_nl = (readslicef_29_22_7((MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_44_nl = nl_MultLoop_acc_44_nl[21:0];
  assign nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1519:1512]));
  assign MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1527:1520]));
  assign MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_43_nl = (readslicef_29_22_7((MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_43_nl = nl_MultLoop_acc_43_nl[21:0];
  assign nl_MultLoop_acc_115_itm_1  = (MultLoop_acc_46_nl) + (MultLoop_acc_45_nl)
      + (MultLoop_acc_44_nl) + (MultLoop_acc_43_nl);
  assign nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1535:1528]));
  assign MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1543:1536]));
  assign MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_42_nl = (readslicef_29_22_7((MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[21:0];
  assign nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1551:1544]));
  assign MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1559:1552]));
  assign MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_41_nl = (readslicef_29_22_7((MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_41_nl = nl_MultLoop_acc_41_nl[21:0];
  assign nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1567:1560]));
  assign MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1575:1568]));
  assign MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_40_nl = (readslicef_29_22_7((MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_40_nl = nl_MultLoop_acc_40_nl[21:0];
  assign nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1583:1576]));
  assign MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1591:1584]));
  assign MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_39_nl = (readslicef_29_22_7((MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_39_nl = nl_MultLoop_acc_39_nl[21:0];
  assign nl_MultLoop_acc_114_itm_1  = (MultLoop_acc_42_nl) + (MultLoop_acc_41_nl)
      + (MultLoop_acc_40_nl) + (MultLoop_acc_39_nl);
  assign nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1599:1592]));
  assign MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1607:1600]));
  assign MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_38_nl = (readslicef_29_22_7((MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_38_nl = nl_MultLoop_acc_38_nl[21:0];
  assign nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1615:1608]));
  assign MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1623:1616]));
  assign MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_37_nl = (readslicef_29_22_7((MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_37_nl = nl_MultLoop_acc_37_nl[21:0];
  assign nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1631:1624]));
  assign MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1639:1632]));
  assign MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_36_nl = (readslicef_29_22_7((MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_36_nl = nl_MultLoop_acc_36_nl[21:0];
  assign nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1647:1640]));
  assign MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1655:1648]));
  assign MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_35_nl = (readslicef_29_22_7((MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_35_nl = nl_MultLoop_acc_35_nl[21:0];
  assign nl_MultLoop_acc_113_itm_1  = (MultLoop_acc_38_nl) + (MultLoop_acc_37_nl)
      + (MultLoop_acc_36_nl) + (MultLoop_acc_35_nl);
  assign nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1663:1656]));
  assign MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1671:1664]));
  assign MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_34_nl = (readslicef_29_22_7((MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_34_nl = nl_MultLoop_acc_34_nl[21:0];
  assign nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1679:1672]));
  assign MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1687:1680]));
  assign MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_33_nl = (readslicef_29_22_7((MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_33_nl = nl_MultLoop_acc_33_nl[21:0];
  assign nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1695:1688]));
  assign MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1703:1696]));
  assign MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_32_nl = (readslicef_29_22_7((MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_32_nl = nl_MultLoop_acc_32_nl[21:0];
  assign nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1711:1704]));
  assign MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1719:1712]));
  assign MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_31_nl = (readslicef_29_22_7((MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_31_nl = nl_MultLoop_acc_31_nl[21:0];
  assign nl_MultLoop_acc_112_itm_1  = (MultLoop_acc_34_nl) + (MultLoop_acc_33_nl)
      + (MultLoop_acc_32_nl) + (MultLoop_acc_31_nl);
  assign nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1727:1720]));
  assign MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1735:1728]));
  assign MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_30_nl = (readslicef_29_22_7((MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_30_nl = nl_MultLoop_acc_30_nl[21:0];
  assign nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1743:1736]));
  assign MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1751:1744]));
  assign MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_29_nl = (readslicef_29_22_7((MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_29_nl = nl_MultLoop_acc_29_nl[21:0];
  assign nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1759:1752]));
  assign MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1767:1760]));
  assign MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_28_nl = (readslicef_29_22_7((MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_28_nl = nl_MultLoop_acc_28_nl[21:0];
  assign nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1775:1768]));
  assign MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1783:1776]));
  assign MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_27_nl = (readslicef_29_22_7((MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_27_nl = nl_MultLoop_acc_27_nl[21:0];
  assign nl_MultLoop_acc_111_itm_1  = (MultLoop_acc_30_nl) + (MultLoop_acc_29_nl)
      + (MultLoop_acc_28_nl) + (MultLoop_acc_27_nl);
  assign nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1791:1784]));
  assign MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1799:1792]));
  assign MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_26_nl = (readslicef_29_22_7((MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_26_nl = nl_MultLoop_acc_26_nl[21:0];
  assign nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1807:1800]));
  assign MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1815:1808]));
  assign MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_25_nl = (readslicef_29_22_7((MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_25_nl = nl_MultLoop_acc_25_nl[21:0];
  assign nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1823:1816]));
  assign MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1831:1824]));
  assign MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_24_nl = (readslicef_29_22_7((MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_24_nl = nl_MultLoop_acc_24_nl[21:0];
  assign nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1839:1832]));
  assign MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1847:1840]));
  assign MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_23_nl = (readslicef_29_22_7((MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_23_nl = nl_MultLoop_acc_23_nl[21:0];
  assign nl_MultLoop_acc_110_itm_1  = (MultLoop_acc_26_nl) + (MultLoop_acc_25_nl)
      + (MultLoop_acc_24_nl) + (MultLoop_acc_23_nl);
  assign nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1855:1848]));
  assign MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1863:1856]));
  assign MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_22_nl = (readslicef_29_22_7((MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_22_nl = nl_MultLoop_acc_22_nl[21:0];
  assign nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1871:1864]));
  assign MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1879:1872]));
  assign MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_21_nl = (readslicef_29_22_7((MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[21:0];
  assign nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1887:1880]));
  assign MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1895:1888]));
  assign MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_20_nl = (readslicef_29_22_7((MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_20_nl = nl_MultLoop_acc_20_nl[21:0];
  assign nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1903:1896]));
  assign MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1911:1904]));
  assign MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_19_nl = (readslicef_29_22_7((MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_19_nl = nl_MultLoop_acc_19_nl[21:0];
  assign nl_MultLoop_acc_109_itm_1  = (MultLoop_acc_22_nl) + (MultLoop_acc_21_nl)
      + (MultLoop_acc_20_nl) + (MultLoop_acc_19_nl);
  assign nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1919:1912]));
  assign MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1927:1920]));
  assign MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_18_nl = (readslicef_29_22_7((MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[21:0];
  assign nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1935:1928]));
  assign MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1943:1936]));
  assign MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_17_nl = (readslicef_29_22_7((MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_17_nl = nl_MultLoop_acc_17_nl[21:0];
  assign nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1951:1944]));
  assign MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1959:1952]));
  assign MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_16_nl = (readslicef_29_22_7((MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_16_nl = nl_MultLoop_acc_16_nl[21:0];
  assign nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1967:1960]));
  assign MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1975:1968]));
  assign MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_15_nl = (readslicef_29_22_7((MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_15_nl = nl_MultLoop_acc_15_nl[21:0];
  assign nl_MultLoop_acc_108_itm_1  = (MultLoop_acc_18_nl) + (MultLoop_acc_17_nl)
      + (MultLoop_acc_16_nl) + (MultLoop_acc_15_nl);
  assign nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1983:1976]));
  assign MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1991:1984]));
  assign MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_14_nl = (readslicef_29_22_7((MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[21:0];
  assign nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1999:1992]));
  assign MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2007:2000]));
  assign MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_13_nl = (readslicef_29_22_7((MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_13_nl = nl_MultLoop_acc_13_nl[21:0];
  assign nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2015:2008]));
  assign MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2023:2016]));
  assign MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_12_nl = (readslicef_29_22_7((MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_12_nl = nl_MultLoop_acc_12_nl[21:0];
  assign nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2031:2024]));
  assign MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2039:2032]));
  assign MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_11_nl = (readslicef_29_22_7((MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_11_nl = nl_MultLoop_acc_11_nl[21:0];
  assign nl_MultLoop_acc_107_itm_1  = (MultLoop_acc_14_nl) + (MultLoop_acc_13_nl)
      + (MultLoop_acc_12_nl) + (MultLoop_acc_11_nl);

  function automatic [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_23_1_22;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 22;
    readslicef_23_1_22 = tmp[0:0];
  end
  endfunction


  function automatic [21:0] readslicef_29_22_7;
    input [28:0] vector;
    reg [28:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_29_22_7 = tmp[21:0];
  end
  endfunction


  function automatic [20:0] readslicef_30_21_9;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_30_21_9 = tmp[20:0];
  end
  endfunction


  function automatic [9:0] conv_s2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_8_11 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_11 = {{3{vector[7]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [29:0] conv_s2u_30_30 ;
    input [29:0]  vector ;
  begin
    conv_s2u_30_30 = vector;
  end
  endfunction


  function automatic [21:0] conv_u2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_u2s_21_22 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10
// ------------------------------------------------------------------


module econ_4x4_d10 (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_triosy_lz, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_triosy_lz, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld, w2_rsc_triosy_lz, b2_rsc_dat,
      b2_rsc_vld, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_triosy_lz, b4_rsc_dat,
      b4_rsc_vld, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_triosy_lz;
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  econ_4x4_d10_core econ_4x4_d10_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz)
    );
endmodule



