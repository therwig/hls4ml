
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_vld_v1 (dat, vld, idat, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             vld;
  input  [width-1:0] idat;
  input              ivld;

  wire   [width-1:0] dat;
  wire               vld;

  assign dat = idat;
  assign vld = ivld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/nnet__relu_layer6_t_result_t_relu_config7__2ad7de4a814a089becf633139a3e7ec975ef_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:07:48 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer6_t_result_t_relu_config7_core
// ------------------------------------------------------------------


module nnet_relu_layer6_t_result_t_relu_config7_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [53:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [53:0] data_rsci_idat;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;

  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [53:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18 , 1'b0
      , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd20),
  .width(32'sd54)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd21),
  .width(32'sd54)) res_rsci (
      .d(nl_res_rsci_d[53:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer6_t_result_t_relu_config7
// ------------------------------------------------------------------


module nnet_relu_layer6_t_result_t_relu_config7 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [53:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer6_t_result_t_relu_config7_core nnet_relu_layer6_t_result_t_relu_config7_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_layer5_t_layer6_t_config6__04a4dab5ef72864301f0c122ebf62e1a90e4_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:07:55 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer5_t_layer6_t_config6_core
// ------------------------------------------------------------------


module nnet_dense_large_layer5_t_layer6_t_config6_core (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input [323:0] weights_rsc_dat;
  input [53:0] biases_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [107:0] data_rsci_idat;
  wire [323:0] weights_rsci_idat;
  wire [53:0] biases_rsci_idat;
  reg [17:0] res_rsci_d_53_36;
  wire [18:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [18:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [18:0] nl_res_rsci_d_17_0;

  wire[17:0] MultLoop_acc_8_nl;
  wire[18:0] nl_MultLoop_acc_8_nl;
  wire[17:0] MultLoop_acc_6_nl;
  wire[18:0] nl_MultLoop_acc_6_nl;
  wire[27:0] MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_5_nl;
  wire[18:0] nl_MultLoop_acc_5_nl;
  wire[27:0] MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_7_nl;
  wire[18:0] nl_MultLoop_acc_7_nl;
  wire[17:0] MultLoop_acc_4_nl;
  wire[18:0] nl_MultLoop_acc_4_nl;
  wire[27:0] MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_18_nl;
  wire[18:0] nl_MultLoop_acc_18_nl;
  wire[17:0] MultLoop_acc_16_nl;
  wire[18:0] nl_MultLoop_acc_16_nl;
  wire[27:0] MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_15_nl;
  wire[18:0] nl_MultLoop_acc_15_nl;
  wire[27:0] MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_17_nl;
  wire[18:0] nl_MultLoop_acc_17_nl;
  wire[17:0] MultLoop_acc_14_nl;
  wire[18:0] nl_MultLoop_acc_14_nl;
  wire[27:0] MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_13_nl;
  wire[18:0] nl_MultLoop_acc_13_nl;
  wire[17:0] MultLoop_acc_11_nl;
  wire[18:0] nl_MultLoop_acc_11_nl;
  wire[27:0] MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_10_nl;
  wire[18:0] nl_MultLoop_acc_10_nl;
  wire[27:0] MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_12_nl;
  wire[18:0] nl_MultLoop_acc_12_nl;
  wire[17:0] MultLoop_acc_9_nl;
  wire[18:0] nl_MultLoop_acc_9_nl;
  wire[27:0] MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [53:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_53_36 , res_rsci_d_35_18 , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd15),
  .width(32'sd108)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd16),
  .width(32'sd54)) res_rsci (
      .d(nl_res_rsci_d[53:0]),
      .z(res_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd17),
  .width(32'sd324)) weights_rsci (
      .dat(weights_rsc_dat),
      .idat(weights_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd18),
  .width(32'sd54)) biases_rsci (
      .dat(biases_rsc_dat),
      .idat(biases_rsci_idat)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_53_36 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
    end
  end
  assign nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[233:216]));
  assign MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[251:234]));
  assign MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_6_nl = (readslicef_28_18_10((MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_6_nl = nl_MultLoop_acc_6_nl[17:0];
  assign nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[269:252]));
  assign MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[287:270]));
  assign MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_5_nl = (readslicef_28_18_10((MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_5_nl = nl_MultLoop_acc_5_nl[17:0];
  assign nl_MultLoop_acc_8_nl = (MultLoop_acc_6_nl) + (MultLoop_acc_5_nl);
  assign MultLoop_acc_8_nl = nl_MultLoop_acc_8_nl[17:0];
  assign nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[305:288]));
  assign MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[323:306]));
  assign MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_4_nl = (readslicef_28_18_10((MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_4_nl = nl_MultLoop_acc_4_nl[17:0];
  assign nl_MultLoop_acc_7_nl = (MultLoop_acc_4_nl) + (biases_rsci_idat[53:36]);
  assign MultLoop_acc_7_nl = nl_MultLoop_acc_7_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_8_nl) + (MultLoop_acc_7_nl);
  assign nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[17:0]));
  assign MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[35:18]));
  assign MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_16_nl = (readslicef_28_18_10((MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_16_nl = nl_MultLoop_acc_16_nl[17:0];
  assign nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[53:36]));
  assign MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[71:54]));
  assign MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_15_nl = (readslicef_28_18_10((MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_15_nl = nl_MultLoop_acc_15_nl[17:0];
  assign nl_MultLoop_acc_18_nl = (MultLoop_acc_16_nl) + (MultLoop_acc_15_nl);
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[17:0];
  assign nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[89:72]));
  assign MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[107:90]));
  assign MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_14_nl = (readslicef_28_18_10((MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[17:0];
  assign nl_MultLoop_acc_17_nl = (MultLoop_acc_14_nl) + (biases_rsci_idat[17:0]);
  assign MultLoop_acc_17_nl = nl_MultLoop_acc_17_nl[17:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_18_nl) + (MultLoop_acc_17_nl);
  assign nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[125:108]));
  assign MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[143:126]));
  assign MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_11_nl = (readslicef_28_18_10((MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_11_nl = nl_MultLoop_acc_11_nl[17:0];
  assign nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[161:144]));
  assign MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[179:162]));
  assign MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_10_nl = (readslicef_28_18_10((MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_10_nl = nl_MultLoop_acc_10_nl[17:0];
  assign nl_MultLoop_acc_13_nl = (MultLoop_acc_11_nl) + (MultLoop_acc_10_nl);
  assign MultLoop_acc_13_nl = nl_MultLoop_acc_13_nl[17:0];
  assign nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[197:180]));
  assign MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[215:198]));
  assign MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_9_nl = (readslicef_28_18_10((MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_9_nl = nl_MultLoop_acc_9_nl[17:0];
  assign nl_MultLoop_acc_12_nl = (MultLoop_acc_9_nl) + (biases_rsci_idat[35:18]);
  assign MultLoop_acc_12_nl = nl_MultLoop_acc_12_nl[17:0];
  assign nl_res_rsci_d_35_18  = (MultLoop_acc_13_nl) + (MultLoop_acc_12_nl);

  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer5_t_layer6_t_config6
// ------------------------------------------------------------------


module nnet_dense_large_layer5_t_layer6_t_config6 (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input [323:0] weights_rsc_dat;
  input [53:0] biases_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_layer5_t_layer6_t_config6_core nnet_dense_large_layer5_t_layer6_t_config6_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .weights_rsc_dat(weights_rsc_dat),
      .biases_rsc_dat(biases_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__relu_layer4_t_layer5_t_relu_config5__9ce8b1180adac085c5d066ac8295b58a9071_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:08:02 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer4_t_layer5_t_relu_config5_core
// ------------------------------------------------------------------


module nnet_relu_layer4_t_layer5_t_relu_config5_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [107:0] data_rsci_idat;
  reg [16:0] res_rsci_d_106_90;
  reg [16:0] res_rsci_d_88_72;
  reg [16:0] res_rsci_d_70_54;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;

  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [107:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_106_90 , 1'b0 , res_rsci_d_88_72 , 1'b0
      , res_rsci_d_70_54 , 1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18 , 1'b0
      , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd13),
  .width(32'sd108)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd14),
  .width(32'sd108)) res_rsci (
      .d(nl_res_rsci_d[107:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_106_90 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
      res_rsci_d_88_72 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_70_54 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_106_90 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[106:90]),
          (readslicef_19_1_18((for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_88_72 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[88:72]),
          (readslicef_19_1_18((for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_70_54 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[70:54]),
          (readslicef_19_1_18((for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[107:90]);
  assign for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[89:72]);
  assign for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[71:54]);
  assign for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer4_t_layer5_t_relu_config5
// ------------------------------------------------------------------


module nnet_relu_layer4_t_layer5_t_relu_config5 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer4_t_layer5_t_relu_config5_core nnet_relu_layer4_t_layer5_t_relu_config5_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_layer3_t_layer4_t_config4__1cb780709f2603aadeb311c7716f7c8c155f2_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:08:16 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4_core
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4_core (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input [2591:0] weights_rsc_dat;
  input [107:0] biases_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [431:0] data_rsci_idat;
  wire [2591:0] weights_rsci_idat;
  wire [107:0] biases_rsci_idat;
  reg [17:0] res_rsci_d_107_90;
  wire [18:0] nl_res_rsci_d_107_90;
  reg [17:0] res_rsci_d_89_72;
  wire [18:0] nl_res_rsci_d_89_72;
  reg [17:0] res_rsci_d_71_54;
  wire [18:0] nl_res_rsci_d_71_54;
  reg [17:0] res_rsci_d_53_36;
  wire [18:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [18:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [18:0] nl_res_rsci_d_17_0;

  wire[17:0] MultLoop_acc_41_nl;
  wire[20:0] nl_MultLoop_acc_41_nl;
  wire[17:0] MultLoop_acc_23_nl;
  wire[18:0] nl_MultLoop_acc_23_nl;
  wire[27:0] MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_22_nl;
  wire[18:0] nl_MultLoop_acc_22_nl;
  wire[27:0] MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_27_nl;
  wire[18:0] nl_MultLoop_acc_27_nl;
  wire[27:0] MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_26_nl;
  wire[18:0] nl_MultLoop_acc_26_nl;
  wire[27:0] MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_25_nl;
  wire[18:0] nl_MultLoop_acc_25_nl;
  wire[27:0] MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_24_nl;
  wire[18:0] nl_MultLoop_acc_24_nl;
  wire[27:0] MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_21_nl;
  wire[18:0] nl_MultLoop_acc_21_nl;
  wire[27:0] MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_20_nl;
  wire[18:0] nl_MultLoop_acc_20_nl;
  wire[27:0] MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_40_nl;
  wire[19:0] nl_MultLoop_acc_40_nl;
  wire[17:0] MultLoop_acc_31_nl;
  wire[18:0] nl_MultLoop_acc_31_nl;
  wire[17:0] MultLoop_acc_19_nl;
  wire[18:0] nl_MultLoop_acc_19_nl;
  wire[27:0] MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_30_nl;
  wire[18:0] nl_MultLoop_acc_30_nl;
  wire[27:0] MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_29_nl;
  wire[18:0] nl_MultLoop_acc_29_nl;
  wire[27:0] MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_28_nl;
  wire[18:0] nl_MultLoop_acc_28_nl;
  wire[27:0] MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_156_nl;
  wire[20:0] nl_MultLoop_acc_156_nl;
  wire[17:0] MultLoop_acc_138_nl;
  wire[18:0] nl_MultLoop_acc_138_nl;
  wire[27:0] MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_137_nl;
  wire[18:0] nl_MultLoop_acc_137_nl;
  wire[27:0] MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_142_nl;
  wire[18:0] nl_MultLoop_acc_142_nl;
  wire[27:0] MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_141_nl;
  wire[18:0] nl_MultLoop_acc_141_nl;
  wire[27:0] MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_140_nl;
  wire[18:0] nl_MultLoop_acc_140_nl;
  wire[27:0] MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_139_nl;
  wire[18:0] nl_MultLoop_acc_139_nl;
  wire[27:0] MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_136_nl;
  wire[18:0] nl_MultLoop_acc_136_nl;
  wire[27:0] MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_135_nl;
  wire[18:0] nl_MultLoop_acc_135_nl;
  wire[27:0] MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_155_nl;
  wire[19:0] nl_MultLoop_acc_155_nl;
  wire[17:0] MultLoop_acc_146_nl;
  wire[18:0] nl_MultLoop_acc_146_nl;
  wire[17:0] MultLoop_acc_134_nl;
  wire[18:0] nl_MultLoop_acc_134_nl;
  wire[27:0] MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_145_nl;
  wire[18:0] nl_MultLoop_acc_145_nl;
  wire[27:0] MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_144_nl;
  wire[18:0] nl_MultLoop_acc_144_nl;
  wire[27:0] MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_143_nl;
  wire[18:0] nl_MultLoop_acc_143_nl;
  wire[27:0] MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_64_nl;
  wire[20:0] nl_MultLoop_acc_64_nl;
  wire[17:0] MultLoop_acc_46_nl;
  wire[18:0] nl_MultLoop_acc_46_nl;
  wire[27:0] MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_45_nl;
  wire[18:0] nl_MultLoop_acc_45_nl;
  wire[27:0] MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_50_nl;
  wire[18:0] nl_MultLoop_acc_50_nl;
  wire[27:0] MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_49_nl;
  wire[18:0] nl_MultLoop_acc_49_nl;
  wire[27:0] MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_48_nl;
  wire[18:0] nl_MultLoop_acc_48_nl;
  wire[27:0] MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_47_nl;
  wire[18:0] nl_MultLoop_acc_47_nl;
  wire[27:0] MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_44_nl;
  wire[18:0] nl_MultLoop_acc_44_nl;
  wire[27:0] MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_43_nl;
  wire[18:0] nl_MultLoop_acc_43_nl;
  wire[27:0] MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_63_nl;
  wire[19:0] nl_MultLoop_acc_63_nl;
  wire[17:0] MultLoop_acc_54_nl;
  wire[18:0] nl_MultLoop_acc_54_nl;
  wire[17:0] MultLoop_acc_42_nl;
  wire[18:0] nl_MultLoop_acc_42_nl;
  wire[27:0] MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_53_nl;
  wire[18:0] nl_MultLoop_acc_53_nl;
  wire[27:0] MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_52_nl;
  wire[18:0] nl_MultLoop_acc_52_nl;
  wire[27:0] MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_51_nl;
  wire[18:0] nl_MultLoop_acc_51_nl;
  wire[27:0] MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_133_nl;
  wire[20:0] nl_MultLoop_acc_133_nl;
  wire[17:0] MultLoop_acc_115_nl;
  wire[18:0] nl_MultLoop_acc_115_nl;
  wire[27:0] MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_114_nl;
  wire[18:0] nl_MultLoop_acc_114_nl;
  wire[27:0] MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_119_nl;
  wire[18:0] nl_MultLoop_acc_119_nl;
  wire[27:0] MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_118_nl;
  wire[18:0] nl_MultLoop_acc_118_nl;
  wire[27:0] MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_117_nl;
  wire[18:0] nl_MultLoop_acc_117_nl;
  wire[27:0] MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_116_nl;
  wire[18:0] nl_MultLoop_acc_116_nl;
  wire[27:0] MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_113_nl;
  wire[18:0] nl_MultLoop_acc_113_nl;
  wire[27:0] MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_112_nl;
  wire[18:0] nl_MultLoop_acc_112_nl;
  wire[27:0] MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_132_nl;
  wire[19:0] nl_MultLoop_acc_132_nl;
  wire[17:0] MultLoop_acc_123_nl;
  wire[18:0] nl_MultLoop_acc_123_nl;
  wire[17:0] MultLoop_acc_111_nl;
  wire[18:0] nl_MultLoop_acc_111_nl;
  wire[27:0] MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_122_nl;
  wire[18:0] nl_MultLoop_acc_122_nl;
  wire[27:0] MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_121_nl;
  wire[18:0] nl_MultLoop_acc_121_nl;
  wire[27:0] MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_120_nl;
  wire[18:0] nl_MultLoop_acc_120_nl;
  wire[27:0] MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_87_nl;
  wire[20:0] nl_MultLoop_acc_87_nl;
  wire[17:0] MultLoop_acc_69_nl;
  wire[18:0] nl_MultLoop_acc_69_nl;
  wire[27:0] MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_68_nl;
  wire[18:0] nl_MultLoop_acc_68_nl;
  wire[27:0] MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_73_nl;
  wire[18:0] nl_MultLoop_acc_73_nl;
  wire[27:0] MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_72_nl;
  wire[18:0] nl_MultLoop_acc_72_nl;
  wire[27:0] MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_71_nl;
  wire[18:0] nl_MultLoop_acc_71_nl;
  wire[27:0] MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_70_nl;
  wire[18:0] nl_MultLoop_acc_70_nl;
  wire[27:0] MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_67_nl;
  wire[18:0] nl_MultLoop_acc_67_nl;
  wire[27:0] MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_66_nl;
  wire[18:0] nl_MultLoop_acc_66_nl;
  wire[27:0] MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_86_nl;
  wire[19:0] nl_MultLoop_acc_86_nl;
  wire[17:0] MultLoop_acc_77_nl;
  wire[18:0] nl_MultLoop_acc_77_nl;
  wire[17:0] MultLoop_acc_65_nl;
  wire[18:0] nl_MultLoop_acc_65_nl;
  wire[27:0] MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_76_nl;
  wire[18:0] nl_MultLoop_acc_76_nl;
  wire[27:0] MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_75_nl;
  wire[18:0] nl_MultLoop_acc_75_nl;
  wire[27:0] MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_74_nl;
  wire[18:0] nl_MultLoop_acc_74_nl;
  wire[27:0] MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_110_nl;
  wire[20:0] nl_MultLoop_acc_110_nl;
  wire[17:0] MultLoop_acc_92_nl;
  wire[18:0] nl_MultLoop_acc_92_nl;
  wire[27:0] MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_91_nl;
  wire[18:0] nl_MultLoop_acc_91_nl;
  wire[27:0] MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_96_nl;
  wire[18:0] nl_MultLoop_acc_96_nl;
  wire[27:0] MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_95_nl;
  wire[18:0] nl_MultLoop_acc_95_nl;
  wire[27:0] MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_94_nl;
  wire[18:0] nl_MultLoop_acc_94_nl;
  wire[27:0] MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_93_nl;
  wire[18:0] nl_MultLoop_acc_93_nl;
  wire[27:0] MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_90_nl;
  wire[18:0] nl_MultLoop_acc_90_nl;
  wire[27:0] MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_89_nl;
  wire[18:0] nl_MultLoop_acc_89_nl;
  wire[27:0] MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_109_nl;
  wire[19:0] nl_MultLoop_acc_109_nl;
  wire[17:0] MultLoop_acc_100_nl;
  wire[18:0] nl_MultLoop_acc_100_nl;
  wire[17:0] MultLoop_acc_88_nl;
  wire[18:0] nl_MultLoop_acc_88_nl;
  wire[27:0] MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_99_nl;
  wire[18:0] nl_MultLoop_acc_99_nl;
  wire[27:0] MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_98_nl;
  wire[18:0] nl_MultLoop_acc_98_nl;
  wire[27:0] MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_97_nl;
  wire[18:0] nl_MultLoop_acc_97_nl;
  wire[27:0] MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [107:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_107_90 , res_rsci_d_89_72 , res_rsci_d_71_54
      , res_rsci_d_53_36 , res_rsci_d_35_18 , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd432)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd108)) res_rsci (
      .d(nl_res_rsci_d[107:0]),
      .z(res_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd10),
  .width(32'sd2592)) weights_rsci (
      .dat(weights_rsc_dat),
      .idat(weights_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd108)) biases_rsci (
      .dat(biases_rsc_dat),
      .idat(biases_rsci_idat)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_107_90 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_89_72 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
      res_rsci_d_71_54 <= 18'b000000000000000000;
      res_rsci_d_53_36 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_107_90 <= nl_res_rsci_d_107_90[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_89_72 <= nl_res_rsci_d_89_72[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
      res_rsci_d_71_54 <= nl_res_rsci_d_71_54[17:0];
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
    end
  end
  assign nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[2429:2412]));
  assign MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[2447:2430]));
  assign MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_23_nl = (readslicef_28_18_10((MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_23_nl = nl_MultLoop_acc_23_nl[17:0];
  assign nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[2465:2448]));
  assign MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[2483:2466]));
  assign MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_22_nl = (readslicef_28_18_10((MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_22_nl = nl_MultLoop_acc_22_nl[17:0];
  assign nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[2285:2268]));
  assign MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[2303:2286]));
  assign MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_27_nl = (readslicef_28_18_10((MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_27_nl = nl_MultLoop_acc_27_nl[17:0];
  assign nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[2321:2304]));
  assign MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[2339:2322]));
  assign MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_26_nl = (readslicef_28_18_10((MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_26_nl = nl_MultLoop_acc_26_nl[17:0];
  assign nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[2357:2340]));
  assign MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[2375:2358]));
  assign MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_25_nl = (readslicef_28_18_10((MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_25_nl = nl_MultLoop_acc_25_nl[17:0];
  assign nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[2393:2376]));
  assign MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[2411:2394]));
  assign MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_24_nl = (readslicef_28_18_10((MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_24_nl = nl_MultLoop_acc_24_nl[17:0];
  assign nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[2501:2484]));
  assign MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[2519:2502]));
  assign MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_21_nl = (readslicef_28_18_10((MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[17:0];
  assign nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[2537:2520]));
  assign MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[2555:2538]));
  assign MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_20_nl = (readslicef_28_18_10((MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_20_nl = nl_MultLoop_acc_20_nl[17:0];
  assign nl_MultLoop_acc_41_nl = (MultLoop_acc_23_nl) + (MultLoop_acc_22_nl) + (MultLoop_acc_27_nl)
      + (MultLoop_acc_26_nl) + (MultLoop_acc_25_nl) + (MultLoop_acc_24_nl) + (MultLoop_acc_21_nl)
      + (MultLoop_acc_20_nl);
  assign MultLoop_acc_41_nl = nl_MultLoop_acc_41_nl[17:0];
  assign nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[2573:2556]));
  assign MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[2591:2574]));
  assign MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_19_nl = (readslicef_28_18_10((MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_19_nl = nl_MultLoop_acc_19_nl[17:0];
  assign nl_MultLoop_acc_31_nl = (MultLoop_acc_19_nl) + (biases_rsci_idat[107:90]);
  assign MultLoop_acc_31_nl = nl_MultLoop_acc_31_nl[17:0];
  assign nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[2177:2160]));
  assign MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[2195:2178]));
  assign MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_30_nl = (readslicef_28_18_10((MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_30_nl = nl_MultLoop_acc_30_nl[17:0];
  assign nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[2213:2196]));
  assign MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[2231:2214]));
  assign MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_29_nl = (readslicef_28_18_10((MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_29_nl = nl_MultLoop_acc_29_nl[17:0];
  assign nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[2249:2232]));
  assign MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[2267:2250]));
  assign MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_28_nl = (readslicef_28_18_10((MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_28_nl = nl_MultLoop_acc_28_nl[17:0];
  assign nl_MultLoop_acc_40_nl = (MultLoop_acc_31_nl) + (MultLoop_acc_30_nl) + (MultLoop_acc_29_nl)
      + (MultLoop_acc_28_nl);
  assign MultLoop_acc_40_nl = nl_MultLoop_acc_40_nl[17:0];
  assign nl_res_rsci_d_107_90  = (MultLoop_acc_41_nl) + (MultLoop_acc_40_nl);
  assign nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[269:252]));
  assign MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[287:270]));
  assign MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_138_nl = (readslicef_28_18_10((MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_138_nl = nl_MultLoop_acc_138_nl[17:0];
  assign nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[305:288]));
  assign MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[323:306]));
  assign MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_137_nl = (readslicef_28_18_10((MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_137_nl = nl_MultLoop_acc_137_nl[17:0];
  assign nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[125:108]));
  assign MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[143:126]));
  assign MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_142_nl = (readslicef_28_18_10((MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_142_nl = nl_MultLoop_acc_142_nl[17:0];
  assign nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[161:144]));
  assign MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[179:162]));
  assign MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_141_nl = (readslicef_28_18_10((MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_141_nl = nl_MultLoop_acc_141_nl[17:0];
  assign nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[197:180]));
  assign MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[215:198]));
  assign MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_140_nl = (readslicef_28_18_10((MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_140_nl = nl_MultLoop_acc_140_nl[17:0];
  assign nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[233:216]));
  assign MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[251:234]));
  assign MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_139_nl = (readslicef_28_18_10((MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_139_nl = nl_MultLoop_acc_139_nl[17:0];
  assign nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[341:324]));
  assign MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[359:342]));
  assign MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_136_nl = (readslicef_28_18_10((MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_136_nl = nl_MultLoop_acc_136_nl[17:0];
  assign nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[377:360]));
  assign MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[395:378]));
  assign MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_135_nl = (readslicef_28_18_10((MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_135_nl = nl_MultLoop_acc_135_nl[17:0];
  assign nl_MultLoop_acc_156_nl = (MultLoop_acc_138_nl) + (MultLoop_acc_137_nl) +
      (MultLoop_acc_142_nl) + (MultLoop_acc_141_nl) + (MultLoop_acc_140_nl) + (MultLoop_acc_139_nl)
      + (MultLoop_acc_136_nl) + (MultLoop_acc_135_nl);
  assign MultLoop_acc_156_nl = nl_MultLoop_acc_156_nl[17:0];
  assign nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[413:396]));
  assign MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[431:414]));
  assign MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_134_nl = (readslicef_28_18_10((MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[17:0];
  assign nl_MultLoop_acc_146_nl = (MultLoop_acc_134_nl) + (biases_rsci_idat[17:0]);
  assign MultLoop_acc_146_nl = nl_MultLoop_acc_146_nl[17:0];
  assign nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[17:0]));
  assign MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[35:18]));
  assign MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_145_nl = (readslicef_28_18_10((MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_145_nl = nl_MultLoop_acc_145_nl[17:0];
  assign nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[53:36]));
  assign MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[71:54]));
  assign MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_144_nl = (readslicef_28_18_10((MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_144_nl = nl_MultLoop_acc_144_nl[17:0];
  assign nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[89:72]));
  assign MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[107:90]));
  assign MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_143_nl = (readslicef_28_18_10((MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[17:0];
  assign nl_MultLoop_acc_155_nl = (MultLoop_acc_146_nl) + (MultLoop_acc_145_nl) +
      (MultLoop_acc_144_nl) + (MultLoop_acc_143_nl);
  assign MultLoop_acc_155_nl = nl_MultLoop_acc_155_nl[17:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_156_nl) + (MultLoop_acc_155_nl);
  assign nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[1997:1980]));
  assign MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[2015:1998]));
  assign MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_46_nl = (readslicef_28_18_10((MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_46_nl = nl_MultLoop_acc_46_nl[17:0];
  assign nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[2033:2016]));
  assign MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[2051:2034]));
  assign MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_45_nl = (readslicef_28_18_10((MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[17:0];
  assign nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[1853:1836]));
  assign MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[1871:1854]));
  assign MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_50_nl = (readslicef_28_18_10((MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_50_nl = nl_MultLoop_acc_50_nl[17:0];
  assign nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[1889:1872]));
  assign MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[1907:1890]));
  assign MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_49_nl = (readslicef_28_18_10((MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_49_nl = nl_MultLoop_acc_49_nl[17:0];
  assign nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[1925:1908]));
  assign MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[1943:1926]));
  assign MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_48_nl = (readslicef_28_18_10((MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_48_nl = nl_MultLoop_acc_48_nl[17:0];
  assign nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[1961:1944]));
  assign MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[1979:1962]));
  assign MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_47_nl = (readslicef_28_18_10((MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_47_nl = nl_MultLoop_acc_47_nl[17:0];
  assign nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[2069:2052]));
  assign MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[2087:2070]));
  assign MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_44_nl = (readslicef_28_18_10((MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_44_nl = nl_MultLoop_acc_44_nl[17:0];
  assign nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[2105:2088]));
  assign MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[2123:2106]));
  assign MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_43_nl = (readslicef_28_18_10((MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_43_nl = nl_MultLoop_acc_43_nl[17:0];
  assign nl_MultLoop_acc_64_nl = (MultLoop_acc_46_nl) + (MultLoop_acc_45_nl) + (MultLoop_acc_50_nl)
      + (MultLoop_acc_49_nl) + (MultLoop_acc_48_nl) + (MultLoop_acc_47_nl) + (MultLoop_acc_44_nl)
      + (MultLoop_acc_43_nl);
  assign MultLoop_acc_64_nl = nl_MultLoop_acc_64_nl[17:0];
  assign nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[2141:2124]));
  assign MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[2159:2142]));
  assign MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_42_nl = (readslicef_28_18_10((MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[17:0];
  assign nl_MultLoop_acc_54_nl = (MultLoop_acc_42_nl) + (biases_rsci_idat[89:72]);
  assign MultLoop_acc_54_nl = nl_MultLoop_acc_54_nl[17:0];
  assign nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[1745:1728]));
  assign MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[1763:1746]));
  assign MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_53_nl = (readslicef_28_18_10((MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[17:0];
  assign nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[1781:1764]));
  assign MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[1799:1782]));
  assign MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_52_nl = (readslicef_28_18_10((MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_52_nl = nl_MultLoop_acc_52_nl[17:0];
  assign nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[1817:1800]));
  assign MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[1835:1818]));
  assign MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_51_nl = (readslicef_28_18_10((MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_51_nl = nl_MultLoop_acc_51_nl[17:0];
  assign nl_MultLoop_acc_63_nl = (MultLoop_acc_54_nl) + (MultLoop_acc_53_nl) + (MultLoop_acc_52_nl)
      + (MultLoop_acc_51_nl);
  assign MultLoop_acc_63_nl = nl_MultLoop_acc_63_nl[17:0];
  assign nl_res_rsci_d_89_72  = (MultLoop_acc_64_nl) + (MultLoop_acc_63_nl);
  assign nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[701:684]));
  assign MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[719:702]));
  assign MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_115_nl = (readslicef_28_18_10((MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_115_nl = nl_MultLoop_acc_115_nl[17:0];
  assign nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[737:720]));
  assign MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[755:738]));
  assign MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_114_nl = (readslicef_28_18_10((MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_114_nl = nl_MultLoop_acc_114_nl[17:0];
  assign nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[557:540]));
  assign MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[575:558]));
  assign MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_119_nl = (readslicef_28_18_10((MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_119_nl = nl_MultLoop_acc_119_nl[17:0];
  assign nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[593:576]));
  assign MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[611:594]));
  assign MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_118_nl = (readslicef_28_18_10((MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_118_nl = nl_MultLoop_acc_118_nl[17:0];
  assign nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[629:612]));
  assign MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[647:630]));
  assign MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_117_nl = (readslicef_28_18_10((MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_117_nl = nl_MultLoop_acc_117_nl[17:0];
  assign nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[665:648]));
  assign MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[683:666]));
  assign MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_116_nl = (readslicef_28_18_10((MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_116_nl = nl_MultLoop_acc_116_nl[17:0];
  assign nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[773:756]));
  assign MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[791:774]));
  assign MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_113_nl = (readslicef_28_18_10((MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_113_nl = nl_MultLoop_acc_113_nl[17:0];
  assign nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[809:792]));
  assign MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[827:810]));
  assign MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_112_nl = (readslicef_28_18_10((MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_112_nl = nl_MultLoop_acc_112_nl[17:0];
  assign nl_MultLoop_acc_133_nl = (MultLoop_acc_115_nl) + (MultLoop_acc_114_nl) +
      (MultLoop_acc_119_nl) + (MultLoop_acc_118_nl) + (MultLoop_acc_117_nl) + (MultLoop_acc_116_nl)
      + (MultLoop_acc_113_nl) + (MultLoop_acc_112_nl);
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[17:0];
  assign nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[845:828]));
  assign MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[863:846]));
  assign MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_111_nl = (readslicef_28_18_10((MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_111_nl = nl_MultLoop_acc_111_nl[17:0];
  assign nl_MultLoop_acc_123_nl = (MultLoop_acc_111_nl) + (biases_rsci_idat[35:18]);
  assign MultLoop_acc_123_nl = nl_MultLoop_acc_123_nl[17:0];
  assign nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[449:432]));
  assign MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[467:450]));
  assign MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_122_nl = (readslicef_28_18_10((MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_122_nl = nl_MultLoop_acc_122_nl[17:0];
  assign nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[485:468]));
  assign MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[503:486]));
  assign MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_121_nl = (readslicef_28_18_10((MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_121_nl = nl_MultLoop_acc_121_nl[17:0];
  assign nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[521:504]));
  assign MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[539:522]));
  assign MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_120_nl = (readslicef_28_18_10((MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_120_nl = nl_MultLoop_acc_120_nl[17:0];
  assign nl_MultLoop_acc_132_nl = (MultLoop_acc_123_nl) + (MultLoop_acc_122_nl) +
      (MultLoop_acc_121_nl) + (MultLoop_acc_120_nl);
  assign MultLoop_acc_132_nl = nl_MultLoop_acc_132_nl[17:0];
  assign nl_res_rsci_d_35_18  = (MultLoop_acc_133_nl) + (MultLoop_acc_132_nl);
  assign nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[1565:1548]));
  assign MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[1583:1566]));
  assign MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_69_nl = (readslicef_28_18_10((MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_69_nl = nl_MultLoop_acc_69_nl[17:0];
  assign nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[1601:1584]));
  assign MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[1619:1602]));
  assign MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_68_nl = (readslicef_28_18_10((MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_68_nl = nl_MultLoop_acc_68_nl[17:0];
  assign nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[1421:1404]));
  assign MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[1439:1422]));
  assign MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_73_nl = (readslicef_28_18_10((MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[17:0];
  assign nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[1457:1440]));
  assign MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[1475:1458]));
  assign MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_72_nl = (readslicef_28_18_10((MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_72_nl = nl_MultLoop_acc_72_nl[17:0];
  assign nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[1493:1476]));
  assign MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[1511:1494]));
  assign MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_71_nl = (readslicef_28_18_10((MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_71_nl = nl_MultLoop_acc_71_nl[17:0];
  assign nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[1529:1512]));
  assign MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[1547:1530]));
  assign MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_70_nl = (readslicef_28_18_10((MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_70_nl = nl_MultLoop_acc_70_nl[17:0];
  assign nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[1637:1620]));
  assign MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[1655:1638]));
  assign MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_67_nl = (readslicef_28_18_10((MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_67_nl = nl_MultLoop_acc_67_nl[17:0];
  assign nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[1673:1656]));
  assign MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[1691:1674]));
  assign MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_66_nl = (readslicef_28_18_10((MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_66_nl = nl_MultLoop_acc_66_nl[17:0];
  assign nl_MultLoop_acc_87_nl = (MultLoop_acc_69_nl) + (MultLoop_acc_68_nl) + (MultLoop_acc_73_nl)
      + (MultLoop_acc_72_nl) + (MultLoop_acc_71_nl) + (MultLoop_acc_70_nl) + (MultLoop_acc_67_nl)
      + (MultLoop_acc_66_nl);
  assign MultLoop_acc_87_nl = nl_MultLoop_acc_87_nl[17:0];
  assign nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[1709:1692]));
  assign MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[1727:1710]));
  assign MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_65_nl = (readslicef_28_18_10((MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[17:0];
  assign nl_MultLoop_acc_77_nl = (MultLoop_acc_65_nl) + (biases_rsci_idat[71:54]);
  assign MultLoop_acc_77_nl = nl_MultLoop_acc_77_nl[17:0];
  assign nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[1313:1296]));
  assign MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[1331:1314]));
  assign MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_76_nl = (readslicef_28_18_10((MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_76_nl = nl_MultLoop_acc_76_nl[17:0];
  assign nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[1349:1332]));
  assign MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[1367:1350]));
  assign MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_75_nl = (readslicef_28_18_10((MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_75_nl = nl_MultLoop_acc_75_nl[17:0];
  assign nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[1385:1368]));
  assign MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[1403:1386]));
  assign MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_74_nl = (readslicef_28_18_10((MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_74_nl = nl_MultLoop_acc_74_nl[17:0];
  assign nl_MultLoop_acc_86_nl = (MultLoop_acc_77_nl) + (MultLoop_acc_76_nl) + (MultLoop_acc_75_nl)
      + (MultLoop_acc_74_nl);
  assign MultLoop_acc_86_nl = nl_MultLoop_acc_86_nl[17:0];
  assign nl_res_rsci_d_71_54  = (MultLoop_acc_87_nl) + (MultLoop_acc_86_nl);
  assign nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[1133:1116]));
  assign MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[1151:1134]));
  assign MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_92_nl = (readslicef_28_18_10((MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_92_nl = nl_MultLoop_acc_92_nl[17:0];
  assign nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[1169:1152]));
  assign MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[1187:1170]));
  assign MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_91_nl = (readslicef_28_18_10((MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_91_nl = nl_MultLoop_acc_91_nl[17:0];
  assign nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[989:972]));
  assign MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[1007:990]));
  assign MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_96_nl = (readslicef_28_18_10((MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_96_nl = nl_MultLoop_acc_96_nl[17:0];
  assign nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[1025:1008]));
  assign MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[1043:1026]));
  assign MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_95_nl = (readslicef_28_18_10((MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_95_nl = nl_MultLoop_acc_95_nl[17:0];
  assign nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[1061:1044]));
  assign MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[1079:1062]));
  assign MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_94_nl = (readslicef_28_18_10((MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_94_nl = nl_MultLoop_acc_94_nl[17:0];
  assign nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[1097:1080]));
  assign MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[1115:1098]));
  assign MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_93_nl = (readslicef_28_18_10((MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_93_nl = nl_MultLoop_acc_93_nl[17:0];
  assign nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[1205:1188]));
  assign MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[1223:1206]));
  assign MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_90_nl = (readslicef_28_18_10((MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_90_nl = nl_MultLoop_acc_90_nl[17:0];
  assign nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[1241:1224]));
  assign MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[1259:1242]));
  assign MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_89_nl = (readslicef_28_18_10((MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_89_nl = nl_MultLoop_acc_89_nl[17:0];
  assign nl_MultLoop_acc_110_nl = (MultLoop_acc_92_nl) + (MultLoop_acc_91_nl) + (MultLoop_acc_96_nl)
      + (MultLoop_acc_95_nl) + (MultLoop_acc_94_nl) + (MultLoop_acc_93_nl) + (MultLoop_acc_90_nl)
      + (MultLoop_acc_89_nl);
  assign MultLoop_acc_110_nl = nl_MultLoop_acc_110_nl[17:0];
  assign nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[1277:1260]));
  assign MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[1295:1278]));
  assign MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_88_nl = (readslicef_28_18_10((MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_88_nl = nl_MultLoop_acc_88_nl[17:0];
  assign nl_MultLoop_acc_100_nl = (MultLoop_acc_88_nl) + (biases_rsci_idat[53:36]);
  assign MultLoop_acc_100_nl = nl_MultLoop_acc_100_nl[17:0];
  assign nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[881:864]));
  assign MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[899:882]));
  assign MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_99_nl = (readslicef_28_18_10((MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_99_nl = nl_MultLoop_acc_99_nl[17:0];
  assign nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[917:900]));
  assign MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[935:918]));
  assign MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_98_nl = (readslicef_28_18_10((MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_98_nl = nl_MultLoop_acc_98_nl[17:0];
  assign nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[953:936]));
  assign MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[971:954]));
  assign MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_97_nl = (readslicef_28_18_10((MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_97_nl = nl_MultLoop_acc_97_nl[17:0];
  assign nl_MultLoop_acc_109_nl = (MultLoop_acc_100_nl) + (MultLoop_acc_99_nl) +
      (MultLoop_acc_98_nl) + (MultLoop_acc_97_nl);
  assign MultLoop_acc_109_nl = nl_MultLoop_acc_109_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_110_nl) + (MultLoop_acc_109_nl);

  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4 (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input [2591:0] weights_rsc_dat;
  input [107:0] biases_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_layer3_t_layer4_t_config4_core nnet_dense_large_layer3_t_layer4_t_config4_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .weights_rsc_dat(weights_rsc_dat),
      .biases_rsc_dat(biases_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__relu_layer2_t_layer3_t_relu_config3__f965bc8c53f54aae1e9689bf95c0a23c1350c_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:08:24 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3_core
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [431:0] data_rsci_idat;
  reg [16:0] res_rsci_d_412_396;
  reg [16:0] res_rsci_d_394_378;
  reg [16:0] res_rsci_d_376_360;
  reg [16:0] res_rsci_d_358_342;
  reg [16:0] res_rsci_d_340_324;
  reg [16:0] res_rsci_d_322_306;
  reg [16:0] res_rsci_d_304_288;
  reg [16:0] res_rsci_d_286_270;
  reg [16:0] res_rsci_d_268_252;
  reg [16:0] res_rsci_d_250_234;
  reg [16:0] res_rsci_d_232_216;
  reg [16:0] res_rsci_d_214_198;
  reg [16:0] res_rsci_d_196_180;
  reg [16:0] res_rsci_d_178_162;
  reg [16:0] res_rsci_d_160_144;
  reg [16:0] res_rsci_d_142_126;
  reg [16:0] res_rsci_d_124_108;
  reg [16:0] res_rsci_d_106_90;
  reg [16:0] res_rsci_d_88_72;
  reg [16:0] res_rsci_d_70_54;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;
  reg [16:0] res_rsci_d_430_414;

  wire[18:0] for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [431:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_430_414 , 1'b0 , res_rsci_d_412_396 ,
      1'b0 , res_rsci_d_394_378 , 1'b0 , res_rsci_d_376_360 , 1'b0 , res_rsci_d_358_342
      , 1'b0 , res_rsci_d_340_324 , 1'b0 , res_rsci_d_322_306 , 1'b0 , res_rsci_d_304_288
      , 1'b0 , res_rsci_d_286_270 , 1'b0 , res_rsci_d_268_252 , 1'b0 , res_rsci_d_250_234
      , 1'b0 , res_rsci_d_232_216 , 1'b0 , res_rsci_d_214_198 , 1'b0 , res_rsci_d_196_180
      , 1'b0 , res_rsci_d_178_162 , 1'b0 , res_rsci_d_160_144 , 1'b0 , res_rsci_d_142_126
      , 1'b0 , res_rsci_d_124_108 , 1'b0 , res_rsci_d_106_90 , 1'b0 , res_rsci_d_88_72
      , 1'b0 , res_rsci_d_70_54 , 1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18
      , 1'b0 , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd432)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd432)) res_rsci (
      .d(nl_res_rsci_d[431:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_430_414 <= 17'b00000000000000000;
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_412_396 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
      res_rsci_d_394_378 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_376_360 <= 17'b00000000000000000;
      res_rsci_d_70_54 <= 17'b00000000000000000;
      res_rsci_d_358_342 <= 17'b00000000000000000;
      res_rsci_d_88_72 <= 17'b00000000000000000;
      res_rsci_d_340_324 <= 17'b00000000000000000;
      res_rsci_d_106_90 <= 17'b00000000000000000;
      res_rsci_d_322_306 <= 17'b00000000000000000;
      res_rsci_d_124_108 <= 17'b00000000000000000;
      res_rsci_d_304_288 <= 17'b00000000000000000;
      res_rsci_d_142_126 <= 17'b00000000000000000;
      res_rsci_d_286_270 <= 17'b00000000000000000;
      res_rsci_d_160_144 <= 17'b00000000000000000;
      res_rsci_d_268_252 <= 17'b00000000000000000;
      res_rsci_d_178_162 <= 17'b00000000000000000;
      res_rsci_d_250_234 <= 17'b00000000000000000;
      res_rsci_d_196_180 <= 17'b00000000000000000;
      res_rsci_d_232_216 <= 17'b00000000000000000;
      res_rsci_d_214_198 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_430_414 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[430:414]),
          (readslicef_19_1_18((for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_412_396 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[412:396]),
          (readslicef_19_1_18((for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_394_378 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[394:378]),
          (readslicef_19_1_18((for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_376_360 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[376:360]),
          (readslicef_19_1_18((for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_70_54 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[70:54]),
          (readslicef_19_1_18((for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_358_342 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[358:342]),
          (readslicef_19_1_18((for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_88_72 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[88:72]),
          (readslicef_19_1_18((for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_340_324 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[340:324]),
          (readslicef_19_1_18((for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_106_90 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[106:90]),
          (readslicef_19_1_18((for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_322_306 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[322:306]),
          (readslicef_19_1_18((for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_124_108 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[124:108]),
          (readslicef_19_1_18((for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_304_288 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[304:288]),
          (readslicef_19_1_18((for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_142_126 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[142:126]),
          (readslicef_19_1_18((for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_286_270 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[286:270]),
          (readslicef_19_1_18((for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_160_144 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[160:144]),
          (readslicef_19_1_18((for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_268_252 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[268:252]),
          (readslicef_19_1_18((for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_178_162 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[178:162]),
          (readslicef_19_1_18((for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_250_234 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[250:234]),
          (readslicef_19_1_18((for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_196_180 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[196:180]),
          (readslicef_19_1_18((for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_232_216 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[232:216]),
          (readslicef_19_1_18((for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_214_198 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[214:198]),
          (readslicef_19_1_18((for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[431:414]);
  assign for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[413:396]);
  assign for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[395:378]);
  assign for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[377:360]);
  assign for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[71:54]);
  assign for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[359:342]);
  assign for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[89:72]);
  assign for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[341:324]);
  assign for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[107:90]);
  assign for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[323:306]);
  assign for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[125:108]);
  assign for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[305:288]);
  assign for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[143:126]);
  assign for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[287:270]);
  assign for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[161:144]);
  assign for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[269:252]);
  assign for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[179:162]);
  assign for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[251:234]);
  assign for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[197:180]);
  assign for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[233:216]);
  assign for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[215:198]);
  assign for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer2_t_layer3_t_relu_config3_core nnet_relu_layer2_t_layer3_t_relu_config3_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_input_t_layer2_t_config2__23a9a06a28f1f911c48f835db6db103c78ba1_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sun Feb 23 21:10:07 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2_core
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2_core (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [863:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input [20735:0] weights_rsc_dat;
  input [431:0] biases_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [863:0] data_rsci_idat;
  wire [20735:0] weights_rsci_idat;
  wire [431:0] biases_rsci_idat;
  reg [17:0] res_rsci_d_431_414;
  wire [18:0] nl_res_rsci_d_431_414;
  reg [17:0] res_rsci_d_413_396;
  wire [18:0] nl_res_rsci_d_413_396;
  reg [17:0] res_rsci_d_395_378;
  wire [18:0] nl_res_rsci_d_395_378;
  reg [17:0] res_rsci_d_377_360;
  wire [18:0] nl_res_rsci_d_377_360;
  reg [17:0] res_rsci_d_359_342;
  wire [18:0] nl_res_rsci_d_359_342;
  reg [17:0] res_rsci_d_341_324;
  wire [18:0] nl_res_rsci_d_341_324;
  reg [17:0] res_rsci_d_323_306;
  wire [18:0] nl_res_rsci_d_323_306;
  reg [17:0] res_rsci_d_305_288;
  wire [18:0] nl_res_rsci_d_305_288;
  reg [17:0] res_rsci_d_287_270;
  wire [18:0] nl_res_rsci_d_287_270;
  reg [17:0] res_rsci_d_269_252;
  wire [18:0] nl_res_rsci_d_269_252;
  reg [17:0] res_rsci_d_251_234;
  wire [18:0] nl_res_rsci_d_251_234;
  reg [17:0] res_rsci_d_233_216;
  wire [18:0] nl_res_rsci_d_233_216;
  reg [17:0] res_rsci_d_215_198;
  wire [18:0] nl_res_rsci_d_215_198;
  reg [17:0] res_rsci_d_197_180;
  wire [18:0] nl_res_rsci_d_197_180;
  reg [17:0] res_rsci_d_179_162;
  wire [18:0] nl_res_rsci_d_179_162;
  reg [17:0] res_rsci_d_161_144;
  wire [18:0] nl_res_rsci_d_161_144;
  reg [17:0] res_rsci_d_143_126;
  wire [18:0] nl_res_rsci_d_143_126;
  reg [17:0] res_rsci_d_125_108;
  wire [18:0] nl_res_rsci_d_125_108;
  reg [17:0] res_rsci_d_107_90;
  wire [18:0] nl_res_rsci_d_107_90;
  reg [17:0] res_rsci_d_89_72;
  wire [18:0] nl_res_rsci_d_89_72;
  reg [17:0] res_rsci_d_71_54;
  wire [18:0] nl_res_rsci_d_71_54;
  reg [17:0] res_rsci_d_53_36;
  wire [18:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [18:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [18:0] nl_res_rsci_d_17_0;

  wire[17:0] MultLoop_acc_159_nl;
  wire[21:0] nl_MultLoop_acc_159_nl;
  wire[17:0] MultLoop_acc_129_nl;
  wire[18:0] nl_MultLoop_acc_129_nl;
  wire[27:0] MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_128_nl;
  wire[18:0] nl_MultLoop_acc_128_nl;
  wire[27:0] MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_127_nl;
  wire[18:0] nl_MultLoop_acc_127_nl;
  wire[27:0] MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_126_nl;
  wire[18:0] nl_MultLoop_acc_126_nl;
  wire[27:0] MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_125_nl;
  wire[18:0] nl_MultLoop_acc_125_nl;
  wire[27:0] MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_124_nl;
  wire[18:0] nl_MultLoop_acc_124_nl;
  wire[27:0] MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_123_nl;
  wire[18:0] nl_MultLoop_acc_123_nl;
  wire[27:0] MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_122_nl;
  wire[18:0] nl_MultLoop_acc_122_nl;
  wire[27:0] MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_117_nl;
  wire[18:0] nl_MultLoop_acc_117_nl;
  wire[27:0] MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_116_nl;
  wire[18:0] nl_MultLoop_acc_116_nl;
  wire[27:0] MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_115_nl;
  wire[18:0] nl_MultLoop_acc_115_nl;
  wire[27:0] MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_114_nl;
  wire[18:0] nl_MultLoop_acc_114_nl;
  wire[27:0] MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_121_nl;
  wire[18:0] nl_MultLoop_acc_121_nl;
  wire[27:0] MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_120_nl;
  wire[18:0] nl_MultLoop_acc_120_nl;
  wire[27:0] MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_119_nl;
  wire[18:0] nl_MultLoop_acc_119_nl;
  wire[27:0] MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_118_nl;
  wire[18:0] nl_MultLoop_acc_118_nl;
  wire[27:0] MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_158_nl;
  wire[20:0] nl_MultLoop_acc_158_nl;
  wire[17:0] MultLoop_acc_133_nl;
  wire[18:0] nl_MultLoop_acc_133_nl;
  wire[27:0] MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_132_nl;
  wire[18:0] nl_MultLoop_acc_132_nl;
  wire[27:0] MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_137_nl;
  wire[18:0] nl_MultLoop_acc_137_nl;
  wire[17:0] MultLoop_acc_113_nl;
  wire[18:0] nl_MultLoop_acc_113_nl;
  wire[27:0] MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_136_nl;
  wire[18:0] nl_MultLoop_acc_136_nl;
  wire[27:0] MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_135_nl;
  wire[18:0] nl_MultLoop_acc_135_nl;
  wire[27:0] MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_134_nl;
  wire[18:0] nl_MultLoop_acc_134_nl;
  wire[27:0] MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_131_nl;
  wire[18:0] nl_MultLoop_acc_131_nl;
  wire[27:0] MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_130_nl;
  wire[18:0] nl_MultLoop_acc_130_nl;
  wire[27:0] MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1240_nl;
  wire[21:0] nl_MultLoop_acc_1240_nl;
  wire[17:0] MultLoop_acc_1210_nl;
  wire[18:0] nl_MultLoop_acc_1210_nl;
  wire[27:0] MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1209_nl;
  wire[18:0] nl_MultLoop_acc_1209_nl;
  wire[27:0] MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1208_nl;
  wire[18:0] nl_MultLoop_acc_1208_nl;
  wire[27:0] MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1207_nl;
  wire[18:0] nl_MultLoop_acc_1207_nl;
  wire[27:0] MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1206_nl;
  wire[18:0] nl_MultLoop_acc_1206_nl;
  wire[27:0] MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1205_nl;
  wire[18:0] nl_MultLoop_acc_1205_nl;
  wire[27:0] MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1204_nl;
  wire[18:0] nl_MultLoop_acc_1204_nl;
  wire[27:0] MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1203_nl;
  wire[18:0] nl_MultLoop_acc_1203_nl;
  wire[27:0] MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1198_nl;
  wire[18:0] nl_MultLoop_acc_1198_nl;
  wire[27:0] MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1197_nl;
  wire[18:0] nl_MultLoop_acc_1197_nl;
  wire[27:0] MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1196_nl;
  wire[18:0] nl_MultLoop_acc_1196_nl;
  wire[27:0] MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1195_nl;
  wire[18:0] nl_MultLoop_acc_1195_nl;
  wire[27:0] MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1202_nl;
  wire[18:0] nl_MultLoop_acc_1202_nl;
  wire[27:0] MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1201_nl;
  wire[18:0] nl_MultLoop_acc_1201_nl;
  wire[27:0] MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1200_nl;
  wire[18:0] nl_MultLoop_acc_1200_nl;
  wire[27:0] MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1199_nl;
  wire[18:0] nl_MultLoop_acc_1199_nl;
  wire[27:0] MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1239_nl;
  wire[20:0] nl_MultLoop_acc_1239_nl;
  wire[17:0] MultLoop_acc_1214_nl;
  wire[18:0] nl_MultLoop_acc_1214_nl;
  wire[27:0] MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1213_nl;
  wire[18:0] nl_MultLoop_acc_1213_nl;
  wire[27:0] MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1218_nl;
  wire[18:0] nl_MultLoop_acc_1218_nl;
  wire[17:0] MultLoop_acc_1194_nl;
  wire[18:0] nl_MultLoop_acc_1194_nl;
  wire[27:0] MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1217_nl;
  wire[18:0] nl_MultLoop_acc_1217_nl;
  wire[27:0] MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1216_nl;
  wire[18:0] nl_MultLoop_acc_1216_nl;
  wire[27:0] MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1215_nl;
  wire[18:0] nl_MultLoop_acc_1215_nl;
  wire[27:0] MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1212_nl;
  wire[18:0] nl_MultLoop_acc_1212_nl;
  wire[27:0] MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1211_nl;
  wire[18:0] nl_MultLoop_acc_1211_nl;
  wire[27:0] MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_206_nl;
  wire[21:0] nl_MultLoop_acc_206_nl;
  wire[17:0] MultLoop_acc_176_nl;
  wire[18:0] nl_MultLoop_acc_176_nl;
  wire[27:0] MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_175_nl;
  wire[18:0] nl_MultLoop_acc_175_nl;
  wire[27:0] MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_174_nl;
  wire[18:0] nl_MultLoop_acc_174_nl;
  wire[27:0] MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_173_nl;
  wire[18:0] nl_MultLoop_acc_173_nl;
  wire[27:0] MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_172_nl;
  wire[18:0] nl_MultLoop_acc_172_nl;
  wire[27:0] MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_171_nl;
  wire[18:0] nl_MultLoop_acc_171_nl;
  wire[27:0] MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_170_nl;
  wire[18:0] nl_MultLoop_acc_170_nl;
  wire[27:0] MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_169_nl;
  wire[18:0] nl_MultLoop_acc_169_nl;
  wire[27:0] MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_164_nl;
  wire[18:0] nl_MultLoop_acc_164_nl;
  wire[27:0] MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_163_nl;
  wire[18:0] nl_MultLoop_acc_163_nl;
  wire[27:0] MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_162_nl;
  wire[18:0] nl_MultLoop_acc_162_nl;
  wire[27:0] MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_161_nl;
  wire[18:0] nl_MultLoop_acc_161_nl;
  wire[27:0] MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_168_nl;
  wire[18:0] nl_MultLoop_acc_168_nl;
  wire[27:0] MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_167_nl;
  wire[18:0] nl_MultLoop_acc_167_nl;
  wire[27:0] MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_166_nl;
  wire[18:0] nl_MultLoop_acc_166_nl;
  wire[27:0] MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_165_nl;
  wire[18:0] nl_MultLoop_acc_165_nl;
  wire[27:0] MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_205_nl;
  wire[20:0] nl_MultLoop_acc_205_nl;
  wire[17:0] MultLoop_acc_180_nl;
  wire[18:0] nl_MultLoop_acc_180_nl;
  wire[27:0] MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_179_nl;
  wire[18:0] nl_MultLoop_acc_179_nl;
  wire[27:0] MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_184_nl;
  wire[18:0] nl_MultLoop_acc_184_nl;
  wire[17:0] MultLoop_acc_160_nl;
  wire[18:0] nl_MultLoop_acc_160_nl;
  wire[27:0] MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_183_nl;
  wire[18:0] nl_MultLoop_acc_183_nl;
  wire[27:0] MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_182_nl;
  wire[18:0] nl_MultLoop_acc_182_nl;
  wire[27:0] MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_181_nl;
  wire[18:0] nl_MultLoop_acc_181_nl;
  wire[27:0] MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_178_nl;
  wire[18:0] nl_MultLoop_acc_178_nl;
  wire[27:0] MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_177_nl;
  wire[18:0] nl_MultLoop_acc_177_nl;
  wire[27:0] MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1193_nl;
  wire[21:0] nl_MultLoop_acc_1193_nl;
  wire[17:0] MultLoop_acc_1163_nl;
  wire[18:0] nl_MultLoop_acc_1163_nl;
  wire[27:0] MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1162_nl;
  wire[18:0] nl_MultLoop_acc_1162_nl;
  wire[27:0] MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1161_nl;
  wire[18:0] nl_MultLoop_acc_1161_nl;
  wire[27:0] MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1160_nl;
  wire[18:0] nl_MultLoop_acc_1160_nl;
  wire[27:0] MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1159_nl;
  wire[18:0] nl_MultLoop_acc_1159_nl;
  wire[27:0] MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1158_nl;
  wire[18:0] nl_MultLoop_acc_1158_nl;
  wire[27:0] MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1157_nl;
  wire[18:0] nl_MultLoop_acc_1157_nl;
  wire[27:0] MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1156_nl;
  wire[18:0] nl_MultLoop_acc_1156_nl;
  wire[27:0] MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1151_nl;
  wire[18:0] nl_MultLoop_acc_1151_nl;
  wire[27:0] MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1150_nl;
  wire[18:0] nl_MultLoop_acc_1150_nl;
  wire[27:0] MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1149_nl;
  wire[18:0] nl_MultLoop_acc_1149_nl;
  wire[27:0] MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1148_nl;
  wire[18:0] nl_MultLoop_acc_1148_nl;
  wire[27:0] MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1155_nl;
  wire[18:0] nl_MultLoop_acc_1155_nl;
  wire[27:0] MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1154_nl;
  wire[18:0] nl_MultLoop_acc_1154_nl;
  wire[27:0] MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1153_nl;
  wire[18:0] nl_MultLoop_acc_1153_nl;
  wire[27:0] MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1152_nl;
  wire[18:0] nl_MultLoop_acc_1152_nl;
  wire[27:0] MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1192_nl;
  wire[20:0] nl_MultLoop_acc_1192_nl;
  wire[17:0] MultLoop_acc_1167_nl;
  wire[18:0] nl_MultLoop_acc_1167_nl;
  wire[27:0] MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1166_nl;
  wire[18:0] nl_MultLoop_acc_1166_nl;
  wire[27:0] MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1171_nl;
  wire[18:0] nl_MultLoop_acc_1171_nl;
  wire[17:0] MultLoop_acc_1147_nl;
  wire[18:0] nl_MultLoop_acc_1147_nl;
  wire[27:0] MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1170_nl;
  wire[18:0] nl_MultLoop_acc_1170_nl;
  wire[27:0] MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1169_nl;
  wire[18:0] nl_MultLoop_acc_1169_nl;
  wire[27:0] MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1168_nl;
  wire[18:0] nl_MultLoop_acc_1168_nl;
  wire[27:0] MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1165_nl;
  wire[18:0] nl_MultLoop_acc_1165_nl;
  wire[27:0] MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1164_nl;
  wire[18:0] nl_MultLoop_acc_1164_nl;
  wire[27:0] MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_253_nl;
  wire[21:0] nl_MultLoop_acc_253_nl;
  wire[17:0] MultLoop_acc_223_nl;
  wire[18:0] nl_MultLoop_acc_223_nl;
  wire[27:0] MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_222_nl;
  wire[18:0] nl_MultLoop_acc_222_nl;
  wire[27:0] MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_221_nl;
  wire[18:0] nl_MultLoop_acc_221_nl;
  wire[27:0] MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_220_nl;
  wire[18:0] nl_MultLoop_acc_220_nl;
  wire[27:0] MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_219_nl;
  wire[18:0] nl_MultLoop_acc_219_nl;
  wire[27:0] MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_218_nl;
  wire[18:0] nl_MultLoop_acc_218_nl;
  wire[27:0] MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_217_nl;
  wire[18:0] nl_MultLoop_acc_217_nl;
  wire[27:0] MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_216_nl;
  wire[18:0] nl_MultLoop_acc_216_nl;
  wire[27:0] MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_211_nl;
  wire[18:0] nl_MultLoop_acc_211_nl;
  wire[27:0] MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_210_nl;
  wire[18:0] nl_MultLoop_acc_210_nl;
  wire[27:0] MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_209_nl;
  wire[18:0] nl_MultLoop_acc_209_nl;
  wire[27:0] MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_208_nl;
  wire[18:0] nl_MultLoop_acc_208_nl;
  wire[27:0] MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_215_nl;
  wire[18:0] nl_MultLoop_acc_215_nl;
  wire[27:0] MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_214_nl;
  wire[18:0] nl_MultLoop_acc_214_nl;
  wire[27:0] MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_213_nl;
  wire[18:0] nl_MultLoop_acc_213_nl;
  wire[27:0] MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_212_nl;
  wire[18:0] nl_MultLoop_acc_212_nl;
  wire[27:0] MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_252_nl;
  wire[20:0] nl_MultLoop_acc_252_nl;
  wire[17:0] MultLoop_acc_227_nl;
  wire[18:0] nl_MultLoop_acc_227_nl;
  wire[27:0] MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_226_nl;
  wire[18:0] nl_MultLoop_acc_226_nl;
  wire[27:0] MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_231_nl;
  wire[18:0] nl_MultLoop_acc_231_nl;
  wire[17:0] MultLoop_acc_207_nl;
  wire[18:0] nl_MultLoop_acc_207_nl;
  wire[27:0] MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_230_nl;
  wire[18:0] nl_MultLoop_acc_230_nl;
  wire[27:0] MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_229_nl;
  wire[18:0] nl_MultLoop_acc_229_nl;
  wire[27:0] MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_228_nl;
  wire[18:0] nl_MultLoop_acc_228_nl;
  wire[27:0] MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_225_nl;
  wire[18:0] nl_MultLoop_acc_225_nl;
  wire[27:0] MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_224_nl;
  wire[18:0] nl_MultLoop_acc_224_nl;
  wire[27:0] MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1146_nl;
  wire[21:0] nl_MultLoop_acc_1146_nl;
  wire[17:0] MultLoop_acc_1116_nl;
  wire[18:0] nl_MultLoop_acc_1116_nl;
  wire[27:0] MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1115_nl;
  wire[18:0] nl_MultLoop_acc_1115_nl;
  wire[27:0] MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1114_nl;
  wire[18:0] nl_MultLoop_acc_1114_nl;
  wire[27:0] MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1113_nl;
  wire[18:0] nl_MultLoop_acc_1113_nl;
  wire[27:0] MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1112_nl;
  wire[18:0] nl_MultLoop_acc_1112_nl;
  wire[27:0] MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1111_nl;
  wire[18:0] nl_MultLoop_acc_1111_nl;
  wire[27:0] MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1110_nl;
  wire[18:0] nl_MultLoop_acc_1110_nl;
  wire[27:0] MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1109_nl;
  wire[18:0] nl_MultLoop_acc_1109_nl;
  wire[27:0] MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1104_nl;
  wire[18:0] nl_MultLoop_acc_1104_nl;
  wire[27:0] MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1103_nl;
  wire[18:0] nl_MultLoop_acc_1103_nl;
  wire[27:0] MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1102_nl;
  wire[18:0] nl_MultLoop_acc_1102_nl;
  wire[27:0] MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1101_nl;
  wire[18:0] nl_MultLoop_acc_1101_nl;
  wire[27:0] MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1108_nl;
  wire[18:0] nl_MultLoop_acc_1108_nl;
  wire[27:0] MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1107_nl;
  wire[18:0] nl_MultLoop_acc_1107_nl;
  wire[27:0] MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1106_nl;
  wire[18:0] nl_MultLoop_acc_1106_nl;
  wire[27:0] MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1105_nl;
  wire[18:0] nl_MultLoop_acc_1105_nl;
  wire[27:0] MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1145_nl;
  wire[20:0] nl_MultLoop_acc_1145_nl;
  wire[17:0] MultLoop_acc_1120_nl;
  wire[18:0] nl_MultLoop_acc_1120_nl;
  wire[27:0] MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1119_nl;
  wire[18:0] nl_MultLoop_acc_1119_nl;
  wire[27:0] MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1124_nl;
  wire[18:0] nl_MultLoop_acc_1124_nl;
  wire[17:0] MultLoop_acc_1100_nl;
  wire[18:0] nl_MultLoop_acc_1100_nl;
  wire[27:0] MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1123_nl;
  wire[18:0] nl_MultLoop_acc_1123_nl;
  wire[27:0] MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1122_nl;
  wire[18:0] nl_MultLoop_acc_1122_nl;
  wire[27:0] MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1121_nl;
  wire[18:0] nl_MultLoop_acc_1121_nl;
  wire[27:0] MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1118_nl;
  wire[18:0] nl_MultLoop_acc_1118_nl;
  wire[27:0] MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1117_nl;
  wire[18:0] nl_MultLoop_acc_1117_nl;
  wire[27:0] MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_300_nl;
  wire[21:0] nl_MultLoop_acc_300_nl;
  wire[17:0] MultLoop_acc_270_nl;
  wire[18:0] nl_MultLoop_acc_270_nl;
  wire[27:0] MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_269_nl;
  wire[18:0] nl_MultLoop_acc_269_nl;
  wire[27:0] MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_268_nl;
  wire[18:0] nl_MultLoop_acc_268_nl;
  wire[27:0] MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_267_nl;
  wire[18:0] nl_MultLoop_acc_267_nl;
  wire[27:0] MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_266_nl;
  wire[18:0] nl_MultLoop_acc_266_nl;
  wire[27:0] MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_265_nl;
  wire[18:0] nl_MultLoop_acc_265_nl;
  wire[27:0] MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_264_nl;
  wire[18:0] nl_MultLoop_acc_264_nl;
  wire[27:0] MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_263_nl;
  wire[18:0] nl_MultLoop_acc_263_nl;
  wire[27:0] MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_258_nl;
  wire[18:0] nl_MultLoop_acc_258_nl;
  wire[27:0] MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_257_nl;
  wire[18:0] nl_MultLoop_acc_257_nl;
  wire[27:0] MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_256_nl;
  wire[18:0] nl_MultLoop_acc_256_nl;
  wire[27:0] MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_255_nl;
  wire[18:0] nl_MultLoop_acc_255_nl;
  wire[27:0] MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_262_nl;
  wire[18:0] nl_MultLoop_acc_262_nl;
  wire[27:0] MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_261_nl;
  wire[18:0] nl_MultLoop_acc_261_nl;
  wire[27:0] MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_260_nl;
  wire[18:0] nl_MultLoop_acc_260_nl;
  wire[27:0] MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_259_nl;
  wire[18:0] nl_MultLoop_acc_259_nl;
  wire[27:0] MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_299_nl;
  wire[20:0] nl_MultLoop_acc_299_nl;
  wire[17:0] MultLoop_acc_274_nl;
  wire[18:0] nl_MultLoop_acc_274_nl;
  wire[27:0] MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_273_nl;
  wire[18:0] nl_MultLoop_acc_273_nl;
  wire[27:0] MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_278_nl;
  wire[18:0] nl_MultLoop_acc_278_nl;
  wire[17:0] MultLoop_acc_254_nl;
  wire[18:0] nl_MultLoop_acc_254_nl;
  wire[27:0] MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_277_nl;
  wire[18:0] nl_MultLoop_acc_277_nl;
  wire[27:0] MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_276_nl;
  wire[18:0] nl_MultLoop_acc_276_nl;
  wire[27:0] MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_275_nl;
  wire[18:0] nl_MultLoop_acc_275_nl;
  wire[27:0] MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_272_nl;
  wire[18:0] nl_MultLoop_acc_272_nl;
  wire[27:0] MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_271_nl;
  wire[18:0] nl_MultLoop_acc_271_nl;
  wire[27:0] MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1099_nl;
  wire[21:0] nl_MultLoop_acc_1099_nl;
  wire[17:0] MultLoop_acc_1069_nl;
  wire[18:0] nl_MultLoop_acc_1069_nl;
  wire[27:0] MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1068_nl;
  wire[18:0] nl_MultLoop_acc_1068_nl;
  wire[27:0] MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1067_nl;
  wire[18:0] nl_MultLoop_acc_1067_nl;
  wire[27:0] MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1066_nl;
  wire[18:0] nl_MultLoop_acc_1066_nl;
  wire[27:0] MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1065_nl;
  wire[18:0] nl_MultLoop_acc_1065_nl;
  wire[27:0] MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1064_nl;
  wire[18:0] nl_MultLoop_acc_1064_nl;
  wire[27:0] MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1063_nl;
  wire[18:0] nl_MultLoop_acc_1063_nl;
  wire[27:0] MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1062_nl;
  wire[18:0] nl_MultLoop_acc_1062_nl;
  wire[27:0] MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1057_nl;
  wire[18:0] nl_MultLoop_acc_1057_nl;
  wire[27:0] MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1056_nl;
  wire[18:0] nl_MultLoop_acc_1056_nl;
  wire[27:0] MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1055_nl;
  wire[18:0] nl_MultLoop_acc_1055_nl;
  wire[27:0] MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1054_nl;
  wire[18:0] nl_MultLoop_acc_1054_nl;
  wire[27:0] MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1061_nl;
  wire[18:0] nl_MultLoop_acc_1061_nl;
  wire[27:0] MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1060_nl;
  wire[18:0] nl_MultLoop_acc_1060_nl;
  wire[27:0] MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1059_nl;
  wire[18:0] nl_MultLoop_acc_1059_nl;
  wire[27:0] MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1058_nl;
  wire[18:0] nl_MultLoop_acc_1058_nl;
  wire[27:0] MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1098_nl;
  wire[20:0] nl_MultLoop_acc_1098_nl;
  wire[17:0] MultLoop_acc_1073_nl;
  wire[18:0] nl_MultLoop_acc_1073_nl;
  wire[27:0] MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1072_nl;
  wire[18:0] nl_MultLoop_acc_1072_nl;
  wire[27:0] MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1077_nl;
  wire[18:0] nl_MultLoop_acc_1077_nl;
  wire[17:0] MultLoop_acc_1053_nl;
  wire[18:0] nl_MultLoop_acc_1053_nl;
  wire[27:0] MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1076_nl;
  wire[18:0] nl_MultLoop_acc_1076_nl;
  wire[27:0] MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1075_nl;
  wire[18:0] nl_MultLoop_acc_1075_nl;
  wire[27:0] MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1074_nl;
  wire[18:0] nl_MultLoop_acc_1074_nl;
  wire[27:0] MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1071_nl;
  wire[18:0] nl_MultLoop_acc_1071_nl;
  wire[27:0] MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1070_nl;
  wire[18:0] nl_MultLoop_acc_1070_nl;
  wire[27:0] MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_347_nl;
  wire[21:0] nl_MultLoop_acc_347_nl;
  wire[17:0] MultLoop_acc_317_nl;
  wire[18:0] nl_MultLoop_acc_317_nl;
  wire[27:0] MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_316_nl;
  wire[18:0] nl_MultLoop_acc_316_nl;
  wire[27:0] MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_315_nl;
  wire[18:0] nl_MultLoop_acc_315_nl;
  wire[27:0] MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_314_nl;
  wire[18:0] nl_MultLoop_acc_314_nl;
  wire[27:0] MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_313_nl;
  wire[18:0] nl_MultLoop_acc_313_nl;
  wire[27:0] MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_312_nl;
  wire[18:0] nl_MultLoop_acc_312_nl;
  wire[27:0] MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_311_nl;
  wire[18:0] nl_MultLoop_acc_311_nl;
  wire[27:0] MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_310_nl;
  wire[18:0] nl_MultLoop_acc_310_nl;
  wire[27:0] MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_305_nl;
  wire[18:0] nl_MultLoop_acc_305_nl;
  wire[27:0] MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_304_nl;
  wire[18:0] nl_MultLoop_acc_304_nl;
  wire[27:0] MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_303_nl;
  wire[18:0] nl_MultLoop_acc_303_nl;
  wire[27:0] MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_302_nl;
  wire[18:0] nl_MultLoop_acc_302_nl;
  wire[27:0] MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_309_nl;
  wire[18:0] nl_MultLoop_acc_309_nl;
  wire[27:0] MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_308_nl;
  wire[18:0] nl_MultLoop_acc_308_nl;
  wire[27:0] MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_307_nl;
  wire[18:0] nl_MultLoop_acc_307_nl;
  wire[27:0] MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_306_nl;
  wire[18:0] nl_MultLoop_acc_306_nl;
  wire[27:0] MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_346_nl;
  wire[20:0] nl_MultLoop_acc_346_nl;
  wire[17:0] MultLoop_acc_321_nl;
  wire[18:0] nl_MultLoop_acc_321_nl;
  wire[27:0] MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_320_nl;
  wire[18:0] nl_MultLoop_acc_320_nl;
  wire[27:0] MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_325_nl;
  wire[18:0] nl_MultLoop_acc_325_nl;
  wire[17:0] MultLoop_acc_301_nl;
  wire[18:0] nl_MultLoop_acc_301_nl;
  wire[27:0] MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_324_nl;
  wire[18:0] nl_MultLoop_acc_324_nl;
  wire[27:0] MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_323_nl;
  wire[18:0] nl_MultLoop_acc_323_nl;
  wire[27:0] MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_322_nl;
  wire[18:0] nl_MultLoop_acc_322_nl;
  wire[27:0] MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_319_nl;
  wire[18:0] nl_MultLoop_acc_319_nl;
  wire[27:0] MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_318_nl;
  wire[18:0] nl_MultLoop_acc_318_nl;
  wire[27:0] MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1052_nl;
  wire[21:0] nl_MultLoop_acc_1052_nl;
  wire[17:0] MultLoop_acc_1022_nl;
  wire[18:0] nl_MultLoop_acc_1022_nl;
  wire[27:0] MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1021_nl;
  wire[18:0] nl_MultLoop_acc_1021_nl;
  wire[27:0] MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1020_nl;
  wire[18:0] nl_MultLoop_acc_1020_nl;
  wire[27:0] MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1019_nl;
  wire[18:0] nl_MultLoop_acc_1019_nl;
  wire[27:0] MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1018_nl;
  wire[18:0] nl_MultLoop_acc_1018_nl;
  wire[27:0] MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1017_nl;
  wire[18:0] nl_MultLoop_acc_1017_nl;
  wire[27:0] MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1016_nl;
  wire[18:0] nl_MultLoop_acc_1016_nl;
  wire[27:0] MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1015_nl;
  wire[18:0] nl_MultLoop_acc_1015_nl;
  wire[27:0] MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1010_nl;
  wire[18:0] nl_MultLoop_acc_1010_nl;
  wire[27:0] MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1009_nl;
  wire[18:0] nl_MultLoop_acc_1009_nl;
  wire[27:0] MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1008_nl;
  wire[18:0] nl_MultLoop_acc_1008_nl;
  wire[27:0] MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1007_nl;
  wire[18:0] nl_MultLoop_acc_1007_nl;
  wire[27:0] MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1014_nl;
  wire[18:0] nl_MultLoop_acc_1014_nl;
  wire[27:0] MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1013_nl;
  wire[18:0] nl_MultLoop_acc_1013_nl;
  wire[27:0] MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1012_nl;
  wire[18:0] nl_MultLoop_acc_1012_nl;
  wire[27:0] MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1011_nl;
  wire[18:0] nl_MultLoop_acc_1011_nl;
  wire[27:0] MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1051_nl;
  wire[20:0] nl_MultLoop_acc_1051_nl;
  wire[17:0] MultLoop_acc_1026_nl;
  wire[18:0] nl_MultLoop_acc_1026_nl;
  wire[27:0] MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1025_nl;
  wire[18:0] nl_MultLoop_acc_1025_nl;
  wire[27:0] MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1030_nl;
  wire[18:0] nl_MultLoop_acc_1030_nl;
  wire[17:0] MultLoop_acc_1006_nl;
  wire[18:0] nl_MultLoop_acc_1006_nl;
  wire[27:0] MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1029_nl;
  wire[18:0] nl_MultLoop_acc_1029_nl;
  wire[27:0] MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1028_nl;
  wire[18:0] nl_MultLoop_acc_1028_nl;
  wire[27:0] MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1027_nl;
  wire[18:0] nl_MultLoop_acc_1027_nl;
  wire[27:0] MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1024_nl;
  wire[18:0] nl_MultLoop_acc_1024_nl;
  wire[27:0] MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1023_nl;
  wire[18:0] nl_MultLoop_acc_1023_nl;
  wire[27:0] MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_394_nl;
  wire[21:0] nl_MultLoop_acc_394_nl;
  wire[17:0] MultLoop_acc_364_nl;
  wire[18:0] nl_MultLoop_acc_364_nl;
  wire[27:0] MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_363_nl;
  wire[18:0] nl_MultLoop_acc_363_nl;
  wire[27:0] MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_362_nl;
  wire[18:0] nl_MultLoop_acc_362_nl;
  wire[27:0] MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_361_nl;
  wire[18:0] nl_MultLoop_acc_361_nl;
  wire[27:0] MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_360_nl;
  wire[18:0] nl_MultLoop_acc_360_nl;
  wire[27:0] MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_359_nl;
  wire[18:0] nl_MultLoop_acc_359_nl;
  wire[27:0] MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_358_nl;
  wire[18:0] nl_MultLoop_acc_358_nl;
  wire[27:0] MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_357_nl;
  wire[18:0] nl_MultLoop_acc_357_nl;
  wire[27:0] MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_352_nl;
  wire[18:0] nl_MultLoop_acc_352_nl;
  wire[27:0] MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_351_nl;
  wire[18:0] nl_MultLoop_acc_351_nl;
  wire[27:0] MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_350_nl;
  wire[18:0] nl_MultLoop_acc_350_nl;
  wire[27:0] MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_349_nl;
  wire[18:0] nl_MultLoop_acc_349_nl;
  wire[27:0] MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_356_nl;
  wire[18:0] nl_MultLoop_acc_356_nl;
  wire[27:0] MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_355_nl;
  wire[18:0] nl_MultLoop_acc_355_nl;
  wire[27:0] MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_354_nl;
  wire[18:0] nl_MultLoop_acc_354_nl;
  wire[27:0] MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_353_nl;
  wire[18:0] nl_MultLoop_acc_353_nl;
  wire[27:0] MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_393_nl;
  wire[20:0] nl_MultLoop_acc_393_nl;
  wire[17:0] MultLoop_acc_368_nl;
  wire[18:0] nl_MultLoop_acc_368_nl;
  wire[27:0] MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_367_nl;
  wire[18:0] nl_MultLoop_acc_367_nl;
  wire[27:0] MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_372_nl;
  wire[18:0] nl_MultLoop_acc_372_nl;
  wire[17:0] MultLoop_acc_348_nl;
  wire[18:0] nl_MultLoop_acc_348_nl;
  wire[27:0] MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_371_nl;
  wire[18:0] nl_MultLoop_acc_371_nl;
  wire[27:0] MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_370_nl;
  wire[18:0] nl_MultLoop_acc_370_nl;
  wire[27:0] MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_369_nl;
  wire[18:0] nl_MultLoop_acc_369_nl;
  wire[27:0] MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_366_nl;
  wire[18:0] nl_MultLoop_acc_366_nl;
  wire[27:0] MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_365_nl;
  wire[18:0] nl_MultLoop_acc_365_nl;
  wire[27:0] MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1005_nl;
  wire[21:0] nl_MultLoop_acc_1005_nl;
  wire[17:0] MultLoop_acc_975_nl;
  wire[18:0] nl_MultLoop_acc_975_nl;
  wire[27:0] MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_974_nl;
  wire[18:0] nl_MultLoop_acc_974_nl;
  wire[27:0] MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_973_nl;
  wire[18:0] nl_MultLoop_acc_973_nl;
  wire[27:0] MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_972_nl;
  wire[18:0] nl_MultLoop_acc_972_nl;
  wire[27:0] MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_971_nl;
  wire[18:0] nl_MultLoop_acc_971_nl;
  wire[27:0] MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_970_nl;
  wire[18:0] nl_MultLoop_acc_970_nl;
  wire[27:0] MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_969_nl;
  wire[18:0] nl_MultLoop_acc_969_nl;
  wire[27:0] MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_968_nl;
  wire[18:0] nl_MultLoop_acc_968_nl;
  wire[27:0] MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_963_nl;
  wire[18:0] nl_MultLoop_acc_963_nl;
  wire[27:0] MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_962_nl;
  wire[18:0] nl_MultLoop_acc_962_nl;
  wire[27:0] MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_961_nl;
  wire[18:0] nl_MultLoop_acc_961_nl;
  wire[27:0] MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_960_nl;
  wire[18:0] nl_MultLoop_acc_960_nl;
  wire[27:0] MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_967_nl;
  wire[18:0] nl_MultLoop_acc_967_nl;
  wire[27:0] MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_966_nl;
  wire[18:0] nl_MultLoop_acc_966_nl;
  wire[27:0] MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_965_nl;
  wire[18:0] nl_MultLoop_acc_965_nl;
  wire[27:0] MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_964_nl;
  wire[18:0] nl_MultLoop_acc_964_nl;
  wire[27:0] MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_1004_nl;
  wire[20:0] nl_MultLoop_acc_1004_nl;
  wire[17:0] MultLoop_acc_979_nl;
  wire[18:0] nl_MultLoop_acc_979_nl;
  wire[27:0] MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_978_nl;
  wire[18:0] nl_MultLoop_acc_978_nl;
  wire[27:0] MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_983_nl;
  wire[18:0] nl_MultLoop_acc_983_nl;
  wire[17:0] MultLoop_acc_959_nl;
  wire[18:0] nl_MultLoop_acc_959_nl;
  wire[27:0] MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_982_nl;
  wire[18:0] nl_MultLoop_acc_982_nl;
  wire[27:0] MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_981_nl;
  wire[18:0] nl_MultLoop_acc_981_nl;
  wire[27:0] MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_980_nl;
  wire[18:0] nl_MultLoop_acc_980_nl;
  wire[27:0] MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_977_nl;
  wire[18:0] nl_MultLoop_acc_977_nl;
  wire[27:0] MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_976_nl;
  wire[18:0] nl_MultLoop_acc_976_nl;
  wire[27:0] MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_441_nl;
  wire[21:0] nl_MultLoop_acc_441_nl;
  wire[17:0] MultLoop_acc_411_nl;
  wire[18:0] nl_MultLoop_acc_411_nl;
  wire[27:0] MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_410_nl;
  wire[18:0] nl_MultLoop_acc_410_nl;
  wire[27:0] MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_409_nl;
  wire[18:0] nl_MultLoop_acc_409_nl;
  wire[27:0] MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_408_nl;
  wire[18:0] nl_MultLoop_acc_408_nl;
  wire[27:0] MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_407_nl;
  wire[18:0] nl_MultLoop_acc_407_nl;
  wire[27:0] MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_406_nl;
  wire[18:0] nl_MultLoop_acc_406_nl;
  wire[27:0] MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_405_nl;
  wire[18:0] nl_MultLoop_acc_405_nl;
  wire[27:0] MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_404_nl;
  wire[18:0] nl_MultLoop_acc_404_nl;
  wire[27:0] MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_399_nl;
  wire[18:0] nl_MultLoop_acc_399_nl;
  wire[27:0] MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_398_nl;
  wire[18:0] nl_MultLoop_acc_398_nl;
  wire[27:0] MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_397_nl;
  wire[18:0] nl_MultLoop_acc_397_nl;
  wire[27:0] MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_396_nl;
  wire[18:0] nl_MultLoop_acc_396_nl;
  wire[27:0] MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_403_nl;
  wire[18:0] nl_MultLoop_acc_403_nl;
  wire[27:0] MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_402_nl;
  wire[18:0] nl_MultLoop_acc_402_nl;
  wire[27:0] MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_401_nl;
  wire[18:0] nl_MultLoop_acc_401_nl;
  wire[27:0] MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_400_nl;
  wire[18:0] nl_MultLoop_acc_400_nl;
  wire[27:0] MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_440_nl;
  wire[20:0] nl_MultLoop_acc_440_nl;
  wire[17:0] MultLoop_acc_415_nl;
  wire[18:0] nl_MultLoop_acc_415_nl;
  wire[27:0] MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_414_nl;
  wire[18:0] nl_MultLoop_acc_414_nl;
  wire[27:0] MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_419_nl;
  wire[18:0] nl_MultLoop_acc_419_nl;
  wire[17:0] MultLoop_acc_395_nl;
  wire[18:0] nl_MultLoop_acc_395_nl;
  wire[27:0] MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_418_nl;
  wire[18:0] nl_MultLoop_acc_418_nl;
  wire[27:0] MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_417_nl;
  wire[18:0] nl_MultLoop_acc_417_nl;
  wire[27:0] MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_416_nl;
  wire[18:0] nl_MultLoop_acc_416_nl;
  wire[27:0] MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_413_nl;
  wire[18:0] nl_MultLoop_acc_413_nl;
  wire[27:0] MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_412_nl;
  wire[18:0] nl_MultLoop_acc_412_nl;
  wire[27:0] MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_958_nl;
  wire[21:0] nl_MultLoop_acc_958_nl;
  wire[17:0] MultLoop_acc_928_nl;
  wire[18:0] nl_MultLoop_acc_928_nl;
  wire[27:0] MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_927_nl;
  wire[18:0] nl_MultLoop_acc_927_nl;
  wire[27:0] MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_926_nl;
  wire[18:0] nl_MultLoop_acc_926_nl;
  wire[27:0] MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_925_nl;
  wire[18:0] nl_MultLoop_acc_925_nl;
  wire[27:0] MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_924_nl;
  wire[18:0] nl_MultLoop_acc_924_nl;
  wire[27:0] MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_923_nl;
  wire[18:0] nl_MultLoop_acc_923_nl;
  wire[27:0] MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_922_nl;
  wire[18:0] nl_MultLoop_acc_922_nl;
  wire[27:0] MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_921_nl;
  wire[18:0] nl_MultLoop_acc_921_nl;
  wire[27:0] MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_916_nl;
  wire[18:0] nl_MultLoop_acc_916_nl;
  wire[27:0] MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_915_nl;
  wire[18:0] nl_MultLoop_acc_915_nl;
  wire[27:0] MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_914_nl;
  wire[18:0] nl_MultLoop_acc_914_nl;
  wire[27:0] MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_913_nl;
  wire[18:0] nl_MultLoop_acc_913_nl;
  wire[27:0] MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_920_nl;
  wire[18:0] nl_MultLoop_acc_920_nl;
  wire[27:0] MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_919_nl;
  wire[18:0] nl_MultLoop_acc_919_nl;
  wire[27:0] MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_918_nl;
  wire[18:0] nl_MultLoop_acc_918_nl;
  wire[27:0] MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_917_nl;
  wire[18:0] nl_MultLoop_acc_917_nl;
  wire[27:0] MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_957_nl;
  wire[20:0] nl_MultLoop_acc_957_nl;
  wire[17:0] MultLoop_acc_932_nl;
  wire[18:0] nl_MultLoop_acc_932_nl;
  wire[27:0] MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_931_nl;
  wire[18:0] nl_MultLoop_acc_931_nl;
  wire[27:0] MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_936_nl;
  wire[18:0] nl_MultLoop_acc_936_nl;
  wire[17:0] MultLoop_acc_912_nl;
  wire[18:0] nl_MultLoop_acc_912_nl;
  wire[27:0] MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_935_nl;
  wire[18:0] nl_MultLoop_acc_935_nl;
  wire[27:0] MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_934_nl;
  wire[18:0] nl_MultLoop_acc_934_nl;
  wire[27:0] MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_933_nl;
  wire[18:0] nl_MultLoop_acc_933_nl;
  wire[27:0] MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_930_nl;
  wire[18:0] nl_MultLoop_acc_930_nl;
  wire[27:0] MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_929_nl;
  wire[18:0] nl_MultLoop_acc_929_nl;
  wire[27:0] MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_488_nl;
  wire[21:0] nl_MultLoop_acc_488_nl;
  wire[17:0] MultLoop_acc_458_nl;
  wire[18:0] nl_MultLoop_acc_458_nl;
  wire[27:0] MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_457_nl;
  wire[18:0] nl_MultLoop_acc_457_nl;
  wire[27:0] MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_456_nl;
  wire[18:0] nl_MultLoop_acc_456_nl;
  wire[27:0] MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_455_nl;
  wire[18:0] nl_MultLoop_acc_455_nl;
  wire[27:0] MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_454_nl;
  wire[18:0] nl_MultLoop_acc_454_nl;
  wire[27:0] MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_453_nl;
  wire[18:0] nl_MultLoop_acc_453_nl;
  wire[27:0] MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_452_nl;
  wire[18:0] nl_MultLoop_acc_452_nl;
  wire[27:0] MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_451_nl;
  wire[18:0] nl_MultLoop_acc_451_nl;
  wire[27:0] MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_446_nl;
  wire[18:0] nl_MultLoop_acc_446_nl;
  wire[27:0] MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_445_nl;
  wire[18:0] nl_MultLoop_acc_445_nl;
  wire[27:0] MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_444_nl;
  wire[18:0] nl_MultLoop_acc_444_nl;
  wire[27:0] MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_443_nl;
  wire[18:0] nl_MultLoop_acc_443_nl;
  wire[27:0] MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_450_nl;
  wire[18:0] nl_MultLoop_acc_450_nl;
  wire[27:0] MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_449_nl;
  wire[18:0] nl_MultLoop_acc_449_nl;
  wire[27:0] MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_448_nl;
  wire[18:0] nl_MultLoop_acc_448_nl;
  wire[27:0] MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_447_nl;
  wire[18:0] nl_MultLoop_acc_447_nl;
  wire[27:0] MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_487_nl;
  wire[20:0] nl_MultLoop_acc_487_nl;
  wire[17:0] MultLoop_acc_462_nl;
  wire[18:0] nl_MultLoop_acc_462_nl;
  wire[27:0] MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_461_nl;
  wire[18:0] nl_MultLoop_acc_461_nl;
  wire[27:0] MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_466_nl;
  wire[18:0] nl_MultLoop_acc_466_nl;
  wire[17:0] MultLoop_acc_442_nl;
  wire[18:0] nl_MultLoop_acc_442_nl;
  wire[27:0] MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_465_nl;
  wire[18:0] nl_MultLoop_acc_465_nl;
  wire[27:0] MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_464_nl;
  wire[18:0] nl_MultLoop_acc_464_nl;
  wire[27:0] MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_463_nl;
  wire[18:0] nl_MultLoop_acc_463_nl;
  wire[27:0] MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_460_nl;
  wire[18:0] nl_MultLoop_acc_460_nl;
  wire[27:0] MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_459_nl;
  wire[18:0] nl_MultLoop_acc_459_nl;
  wire[27:0] MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_911_nl;
  wire[21:0] nl_MultLoop_acc_911_nl;
  wire[17:0] MultLoop_acc_881_nl;
  wire[18:0] nl_MultLoop_acc_881_nl;
  wire[27:0] MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_880_nl;
  wire[18:0] nl_MultLoop_acc_880_nl;
  wire[27:0] MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_879_nl;
  wire[18:0] nl_MultLoop_acc_879_nl;
  wire[27:0] MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_878_nl;
  wire[18:0] nl_MultLoop_acc_878_nl;
  wire[27:0] MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_877_nl;
  wire[18:0] nl_MultLoop_acc_877_nl;
  wire[27:0] MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_876_nl;
  wire[18:0] nl_MultLoop_acc_876_nl;
  wire[27:0] MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_875_nl;
  wire[18:0] nl_MultLoop_acc_875_nl;
  wire[27:0] MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_874_nl;
  wire[18:0] nl_MultLoop_acc_874_nl;
  wire[27:0] MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_869_nl;
  wire[18:0] nl_MultLoop_acc_869_nl;
  wire[27:0] MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_868_nl;
  wire[18:0] nl_MultLoop_acc_868_nl;
  wire[27:0] MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_867_nl;
  wire[18:0] nl_MultLoop_acc_867_nl;
  wire[27:0] MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_866_nl;
  wire[18:0] nl_MultLoop_acc_866_nl;
  wire[27:0] MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_873_nl;
  wire[18:0] nl_MultLoop_acc_873_nl;
  wire[27:0] MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_872_nl;
  wire[18:0] nl_MultLoop_acc_872_nl;
  wire[27:0] MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_871_nl;
  wire[18:0] nl_MultLoop_acc_871_nl;
  wire[27:0] MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_870_nl;
  wire[18:0] nl_MultLoop_acc_870_nl;
  wire[27:0] MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_910_nl;
  wire[20:0] nl_MultLoop_acc_910_nl;
  wire[17:0] MultLoop_acc_885_nl;
  wire[18:0] nl_MultLoop_acc_885_nl;
  wire[27:0] MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_884_nl;
  wire[18:0] nl_MultLoop_acc_884_nl;
  wire[27:0] MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_889_nl;
  wire[18:0] nl_MultLoop_acc_889_nl;
  wire[17:0] MultLoop_acc_865_nl;
  wire[18:0] nl_MultLoop_acc_865_nl;
  wire[27:0] MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_888_nl;
  wire[18:0] nl_MultLoop_acc_888_nl;
  wire[27:0] MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_887_nl;
  wire[18:0] nl_MultLoop_acc_887_nl;
  wire[27:0] MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_886_nl;
  wire[18:0] nl_MultLoop_acc_886_nl;
  wire[27:0] MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_883_nl;
  wire[18:0] nl_MultLoop_acc_883_nl;
  wire[27:0] MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_882_nl;
  wire[18:0] nl_MultLoop_acc_882_nl;
  wire[27:0] MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_535_nl;
  wire[21:0] nl_MultLoop_acc_535_nl;
  wire[17:0] MultLoop_acc_505_nl;
  wire[18:0] nl_MultLoop_acc_505_nl;
  wire[27:0] MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_504_nl;
  wire[18:0] nl_MultLoop_acc_504_nl;
  wire[27:0] MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_503_nl;
  wire[18:0] nl_MultLoop_acc_503_nl;
  wire[27:0] MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_502_nl;
  wire[18:0] nl_MultLoop_acc_502_nl;
  wire[27:0] MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_501_nl;
  wire[18:0] nl_MultLoop_acc_501_nl;
  wire[27:0] MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_500_nl;
  wire[18:0] nl_MultLoop_acc_500_nl;
  wire[27:0] MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_499_nl;
  wire[18:0] nl_MultLoop_acc_499_nl;
  wire[27:0] MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_498_nl;
  wire[18:0] nl_MultLoop_acc_498_nl;
  wire[27:0] MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_493_nl;
  wire[18:0] nl_MultLoop_acc_493_nl;
  wire[27:0] MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_492_nl;
  wire[18:0] nl_MultLoop_acc_492_nl;
  wire[27:0] MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_491_nl;
  wire[18:0] nl_MultLoop_acc_491_nl;
  wire[27:0] MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_490_nl;
  wire[18:0] nl_MultLoop_acc_490_nl;
  wire[27:0] MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_497_nl;
  wire[18:0] nl_MultLoop_acc_497_nl;
  wire[27:0] MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_496_nl;
  wire[18:0] nl_MultLoop_acc_496_nl;
  wire[27:0] MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_495_nl;
  wire[18:0] nl_MultLoop_acc_495_nl;
  wire[27:0] MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_494_nl;
  wire[18:0] nl_MultLoop_acc_494_nl;
  wire[27:0] MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_534_nl;
  wire[20:0] nl_MultLoop_acc_534_nl;
  wire[17:0] MultLoop_acc_509_nl;
  wire[18:0] nl_MultLoop_acc_509_nl;
  wire[27:0] MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_508_nl;
  wire[18:0] nl_MultLoop_acc_508_nl;
  wire[27:0] MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_513_nl;
  wire[18:0] nl_MultLoop_acc_513_nl;
  wire[17:0] MultLoop_acc_489_nl;
  wire[18:0] nl_MultLoop_acc_489_nl;
  wire[27:0] MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_512_nl;
  wire[18:0] nl_MultLoop_acc_512_nl;
  wire[27:0] MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_511_nl;
  wire[18:0] nl_MultLoop_acc_511_nl;
  wire[27:0] MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_510_nl;
  wire[18:0] nl_MultLoop_acc_510_nl;
  wire[27:0] MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_507_nl;
  wire[18:0] nl_MultLoop_acc_507_nl;
  wire[27:0] MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_506_nl;
  wire[18:0] nl_MultLoop_acc_506_nl;
  wire[27:0] MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_864_nl;
  wire[21:0] nl_MultLoop_acc_864_nl;
  wire[17:0] MultLoop_acc_834_nl;
  wire[18:0] nl_MultLoop_acc_834_nl;
  wire[27:0] MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_833_nl;
  wire[18:0] nl_MultLoop_acc_833_nl;
  wire[27:0] MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_832_nl;
  wire[18:0] nl_MultLoop_acc_832_nl;
  wire[27:0] MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_831_nl;
  wire[18:0] nl_MultLoop_acc_831_nl;
  wire[27:0] MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_830_nl;
  wire[18:0] nl_MultLoop_acc_830_nl;
  wire[27:0] MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_829_nl;
  wire[18:0] nl_MultLoop_acc_829_nl;
  wire[27:0] MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_828_nl;
  wire[18:0] nl_MultLoop_acc_828_nl;
  wire[27:0] MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_827_nl;
  wire[18:0] nl_MultLoop_acc_827_nl;
  wire[27:0] MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_822_nl;
  wire[18:0] nl_MultLoop_acc_822_nl;
  wire[27:0] MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_821_nl;
  wire[18:0] nl_MultLoop_acc_821_nl;
  wire[27:0] MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_820_nl;
  wire[18:0] nl_MultLoop_acc_820_nl;
  wire[27:0] MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_819_nl;
  wire[18:0] nl_MultLoop_acc_819_nl;
  wire[27:0] MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_826_nl;
  wire[18:0] nl_MultLoop_acc_826_nl;
  wire[27:0] MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_825_nl;
  wire[18:0] nl_MultLoop_acc_825_nl;
  wire[27:0] MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_824_nl;
  wire[18:0] nl_MultLoop_acc_824_nl;
  wire[27:0] MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_823_nl;
  wire[18:0] nl_MultLoop_acc_823_nl;
  wire[27:0] MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_863_nl;
  wire[20:0] nl_MultLoop_acc_863_nl;
  wire[17:0] MultLoop_acc_838_nl;
  wire[18:0] nl_MultLoop_acc_838_nl;
  wire[27:0] MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_837_nl;
  wire[18:0] nl_MultLoop_acc_837_nl;
  wire[27:0] MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_842_nl;
  wire[18:0] nl_MultLoop_acc_842_nl;
  wire[17:0] MultLoop_acc_818_nl;
  wire[18:0] nl_MultLoop_acc_818_nl;
  wire[27:0] MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_841_nl;
  wire[18:0] nl_MultLoop_acc_841_nl;
  wire[27:0] MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_840_nl;
  wire[18:0] nl_MultLoop_acc_840_nl;
  wire[27:0] MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_839_nl;
  wire[18:0] nl_MultLoop_acc_839_nl;
  wire[27:0] MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_836_nl;
  wire[18:0] nl_MultLoop_acc_836_nl;
  wire[27:0] MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_835_nl;
  wire[18:0] nl_MultLoop_acc_835_nl;
  wire[27:0] MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_582_nl;
  wire[21:0] nl_MultLoop_acc_582_nl;
  wire[17:0] MultLoop_acc_552_nl;
  wire[18:0] nl_MultLoop_acc_552_nl;
  wire[27:0] MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_551_nl;
  wire[18:0] nl_MultLoop_acc_551_nl;
  wire[27:0] MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_550_nl;
  wire[18:0] nl_MultLoop_acc_550_nl;
  wire[27:0] MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_549_nl;
  wire[18:0] nl_MultLoop_acc_549_nl;
  wire[27:0] MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_548_nl;
  wire[18:0] nl_MultLoop_acc_548_nl;
  wire[27:0] MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_547_nl;
  wire[18:0] nl_MultLoop_acc_547_nl;
  wire[27:0] MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_546_nl;
  wire[18:0] nl_MultLoop_acc_546_nl;
  wire[27:0] MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_545_nl;
  wire[18:0] nl_MultLoop_acc_545_nl;
  wire[27:0] MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_540_nl;
  wire[18:0] nl_MultLoop_acc_540_nl;
  wire[27:0] MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_539_nl;
  wire[18:0] nl_MultLoop_acc_539_nl;
  wire[27:0] MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_538_nl;
  wire[18:0] nl_MultLoop_acc_538_nl;
  wire[27:0] MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_537_nl;
  wire[18:0] nl_MultLoop_acc_537_nl;
  wire[27:0] MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_544_nl;
  wire[18:0] nl_MultLoop_acc_544_nl;
  wire[27:0] MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_543_nl;
  wire[18:0] nl_MultLoop_acc_543_nl;
  wire[27:0] MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_542_nl;
  wire[18:0] nl_MultLoop_acc_542_nl;
  wire[27:0] MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_541_nl;
  wire[18:0] nl_MultLoop_acc_541_nl;
  wire[27:0] MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_581_nl;
  wire[20:0] nl_MultLoop_acc_581_nl;
  wire[17:0] MultLoop_acc_556_nl;
  wire[18:0] nl_MultLoop_acc_556_nl;
  wire[27:0] MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_555_nl;
  wire[18:0] nl_MultLoop_acc_555_nl;
  wire[27:0] MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_560_nl;
  wire[18:0] nl_MultLoop_acc_560_nl;
  wire[17:0] MultLoop_acc_536_nl;
  wire[18:0] nl_MultLoop_acc_536_nl;
  wire[27:0] MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_559_nl;
  wire[18:0] nl_MultLoop_acc_559_nl;
  wire[27:0] MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_558_nl;
  wire[18:0] nl_MultLoop_acc_558_nl;
  wire[27:0] MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_557_nl;
  wire[18:0] nl_MultLoop_acc_557_nl;
  wire[27:0] MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_554_nl;
  wire[18:0] nl_MultLoop_acc_554_nl;
  wire[27:0] MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_553_nl;
  wire[18:0] nl_MultLoop_acc_553_nl;
  wire[27:0] MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_817_nl;
  wire[21:0] nl_MultLoop_acc_817_nl;
  wire[17:0] MultLoop_acc_787_nl;
  wire[18:0] nl_MultLoop_acc_787_nl;
  wire[27:0] MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_786_nl;
  wire[18:0] nl_MultLoop_acc_786_nl;
  wire[27:0] MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_785_nl;
  wire[18:0] nl_MultLoop_acc_785_nl;
  wire[27:0] MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_784_nl;
  wire[18:0] nl_MultLoop_acc_784_nl;
  wire[27:0] MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_783_nl;
  wire[18:0] nl_MultLoop_acc_783_nl;
  wire[27:0] MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_782_nl;
  wire[18:0] nl_MultLoop_acc_782_nl;
  wire[27:0] MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_781_nl;
  wire[18:0] nl_MultLoop_acc_781_nl;
  wire[27:0] MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_780_nl;
  wire[18:0] nl_MultLoop_acc_780_nl;
  wire[27:0] MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_775_nl;
  wire[18:0] nl_MultLoop_acc_775_nl;
  wire[27:0] MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_774_nl;
  wire[18:0] nl_MultLoop_acc_774_nl;
  wire[27:0] MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_773_nl;
  wire[18:0] nl_MultLoop_acc_773_nl;
  wire[27:0] MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_772_nl;
  wire[18:0] nl_MultLoop_acc_772_nl;
  wire[27:0] MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_779_nl;
  wire[18:0] nl_MultLoop_acc_779_nl;
  wire[27:0] MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_778_nl;
  wire[18:0] nl_MultLoop_acc_778_nl;
  wire[27:0] MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_777_nl;
  wire[18:0] nl_MultLoop_acc_777_nl;
  wire[27:0] MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_776_nl;
  wire[18:0] nl_MultLoop_acc_776_nl;
  wire[27:0] MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_816_nl;
  wire[20:0] nl_MultLoop_acc_816_nl;
  wire[17:0] MultLoop_acc_791_nl;
  wire[18:0] nl_MultLoop_acc_791_nl;
  wire[27:0] MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_790_nl;
  wire[18:0] nl_MultLoop_acc_790_nl;
  wire[27:0] MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_795_nl;
  wire[18:0] nl_MultLoop_acc_795_nl;
  wire[17:0] MultLoop_acc_771_nl;
  wire[18:0] nl_MultLoop_acc_771_nl;
  wire[27:0] MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_794_nl;
  wire[18:0] nl_MultLoop_acc_794_nl;
  wire[27:0] MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_793_nl;
  wire[18:0] nl_MultLoop_acc_793_nl;
  wire[27:0] MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_792_nl;
  wire[18:0] nl_MultLoop_acc_792_nl;
  wire[27:0] MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_789_nl;
  wire[18:0] nl_MultLoop_acc_789_nl;
  wire[27:0] MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_788_nl;
  wire[18:0] nl_MultLoop_acc_788_nl;
  wire[27:0] MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_629_nl;
  wire[21:0] nl_MultLoop_acc_629_nl;
  wire[17:0] MultLoop_acc_599_nl;
  wire[18:0] nl_MultLoop_acc_599_nl;
  wire[27:0] MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_598_nl;
  wire[18:0] nl_MultLoop_acc_598_nl;
  wire[27:0] MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_597_nl;
  wire[18:0] nl_MultLoop_acc_597_nl;
  wire[27:0] MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_596_nl;
  wire[18:0] nl_MultLoop_acc_596_nl;
  wire[27:0] MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_595_nl;
  wire[18:0] nl_MultLoop_acc_595_nl;
  wire[27:0] MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_594_nl;
  wire[18:0] nl_MultLoop_acc_594_nl;
  wire[27:0] MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_593_nl;
  wire[18:0] nl_MultLoop_acc_593_nl;
  wire[27:0] MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_592_nl;
  wire[18:0] nl_MultLoop_acc_592_nl;
  wire[27:0] MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_587_nl;
  wire[18:0] nl_MultLoop_acc_587_nl;
  wire[27:0] MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_586_nl;
  wire[18:0] nl_MultLoop_acc_586_nl;
  wire[27:0] MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_585_nl;
  wire[18:0] nl_MultLoop_acc_585_nl;
  wire[27:0] MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_584_nl;
  wire[18:0] nl_MultLoop_acc_584_nl;
  wire[27:0] MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_591_nl;
  wire[18:0] nl_MultLoop_acc_591_nl;
  wire[27:0] MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_590_nl;
  wire[18:0] nl_MultLoop_acc_590_nl;
  wire[27:0] MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_589_nl;
  wire[18:0] nl_MultLoop_acc_589_nl;
  wire[27:0] MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_588_nl;
  wire[18:0] nl_MultLoop_acc_588_nl;
  wire[27:0] MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_628_nl;
  wire[20:0] nl_MultLoop_acc_628_nl;
  wire[17:0] MultLoop_acc_603_nl;
  wire[18:0] nl_MultLoop_acc_603_nl;
  wire[27:0] MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_602_nl;
  wire[18:0] nl_MultLoop_acc_602_nl;
  wire[27:0] MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_607_nl;
  wire[18:0] nl_MultLoop_acc_607_nl;
  wire[17:0] MultLoop_acc_583_nl;
  wire[18:0] nl_MultLoop_acc_583_nl;
  wire[27:0] MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_606_nl;
  wire[18:0] nl_MultLoop_acc_606_nl;
  wire[27:0] MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_605_nl;
  wire[18:0] nl_MultLoop_acc_605_nl;
  wire[27:0] MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_604_nl;
  wire[18:0] nl_MultLoop_acc_604_nl;
  wire[27:0] MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_601_nl;
  wire[18:0] nl_MultLoop_acc_601_nl;
  wire[27:0] MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_600_nl;
  wire[18:0] nl_MultLoop_acc_600_nl;
  wire[27:0] MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_770_nl;
  wire[21:0] nl_MultLoop_acc_770_nl;
  wire[17:0] MultLoop_acc_740_nl;
  wire[18:0] nl_MultLoop_acc_740_nl;
  wire[27:0] MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_739_nl;
  wire[18:0] nl_MultLoop_acc_739_nl;
  wire[27:0] MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_738_nl;
  wire[18:0] nl_MultLoop_acc_738_nl;
  wire[27:0] MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_737_nl;
  wire[18:0] nl_MultLoop_acc_737_nl;
  wire[27:0] MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_736_nl;
  wire[18:0] nl_MultLoop_acc_736_nl;
  wire[27:0] MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_735_nl;
  wire[18:0] nl_MultLoop_acc_735_nl;
  wire[27:0] MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_734_nl;
  wire[18:0] nl_MultLoop_acc_734_nl;
  wire[27:0] MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_733_nl;
  wire[18:0] nl_MultLoop_acc_733_nl;
  wire[27:0] MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_728_nl;
  wire[18:0] nl_MultLoop_acc_728_nl;
  wire[27:0] MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_727_nl;
  wire[18:0] nl_MultLoop_acc_727_nl;
  wire[27:0] MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_726_nl;
  wire[18:0] nl_MultLoop_acc_726_nl;
  wire[27:0] MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_725_nl;
  wire[18:0] nl_MultLoop_acc_725_nl;
  wire[27:0] MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_732_nl;
  wire[18:0] nl_MultLoop_acc_732_nl;
  wire[27:0] MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_731_nl;
  wire[18:0] nl_MultLoop_acc_731_nl;
  wire[27:0] MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_730_nl;
  wire[18:0] nl_MultLoop_acc_730_nl;
  wire[27:0] MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_729_nl;
  wire[18:0] nl_MultLoop_acc_729_nl;
  wire[27:0] MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_769_nl;
  wire[20:0] nl_MultLoop_acc_769_nl;
  wire[17:0] MultLoop_acc_744_nl;
  wire[18:0] nl_MultLoop_acc_744_nl;
  wire[27:0] MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_743_nl;
  wire[18:0] nl_MultLoop_acc_743_nl;
  wire[27:0] MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_748_nl;
  wire[18:0] nl_MultLoop_acc_748_nl;
  wire[17:0] MultLoop_acc_724_nl;
  wire[18:0] nl_MultLoop_acc_724_nl;
  wire[27:0] MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_747_nl;
  wire[18:0] nl_MultLoop_acc_747_nl;
  wire[27:0] MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_746_nl;
  wire[18:0] nl_MultLoop_acc_746_nl;
  wire[27:0] MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_745_nl;
  wire[18:0] nl_MultLoop_acc_745_nl;
  wire[27:0] MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_742_nl;
  wire[18:0] nl_MultLoop_acc_742_nl;
  wire[27:0] MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_741_nl;
  wire[18:0] nl_MultLoop_acc_741_nl;
  wire[27:0] MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_676_nl;
  wire[21:0] nl_MultLoop_acc_676_nl;
  wire[17:0] MultLoop_acc_646_nl;
  wire[18:0] nl_MultLoop_acc_646_nl;
  wire[27:0] MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_645_nl;
  wire[18:0] nl_MultLoop_acc_645_nl;
  wire[27:0] MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_644_nl;
  wire[18:0] nl_MultLoop_acc_644_nl;
  wire[27:0] MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_643_nl;
  wire[18:0] nl_MultLoop_acc_643_nl;
  wire[27:0] MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_642_nl;
  wire[18:0] nl_MultLoop_acc_642_nl;
  wire[27:0] MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_641_nl;
  wire[18:0] nl_MultLoop_acc_641_nl;
  wire[27:0] MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_640_nl;
  wire[18:0] nl_MultLoop_acc_640_nl;
  wire[27:0] MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_639_nl;
  wire[18:0] nl_MultLoop_acc_639_nl;
  wire[27:0] MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_634_nl;
  wire[18:0] nl_MultLoop_acc_634_nl;
  wire[27:0] MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_633_nl;
  wire[18:0] nl_MultLoop_acc_633_nl;
  wire[27:0] MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_632_nl;
  wire[18:0] nl_MultLoop_acc_632_nl;
  wire[27:0] MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_631_nl;
  wire[18:0] nl_MultLoop_acc_631_nl;
  wire[27:0] MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_638_nl;
  wire[18:0] nl_MultLoop_acc_638_nl;
  wire[27:0] MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_637_nl;
  wire[18:0] nl_MultLoop_acc_637_nl;
  wire[27:0] MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_636_nl;
  wire[18:0] nl_MultLoop_acc_636_nl;
  wire[27:0] MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_635_nl;
  wire[18:0] nl_MultLoop_acc_635_nl;
  wire[27:0] MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_675_nl;
  wire[20:0] nl_MultLoop_acc_675_nl;
  wire[17:0] MultLoop_acc_650_nl;
  wire[18:0] nl_MultLoop_acc_650_nl;
  wire[27:0] MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_649_nl;
  wire[18:0] nl_MultLoop_acc_649_nl;
  wire[27:0] MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_654_nl;
  wire[18:0] nl_MultLoop_acc_654_nl;
  wire[17:0] MultLoop_acc_630_nl;
  wire[18:0] nl_MultLoop_acc_630_nl;
  wire[27:0] MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_653_nl;
  wire[18:0] nl_MultLoop_acc_653_nl;
  wire[27:0] MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_652_nl;
  wire[18:0] nl_MultLoop_acc_652_nl;
  wire[27:0] MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_651_nl;
  wire[18:0] nl_MultLoop_acc_651_nl;
  wire[27:0] MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_648_nl;
  wire[18:0] nl_MultLoop_acc_648_nl;
  wire[27:0] MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_647_nl;
  wire[18:0] nl_MultLoop_acc_647_nl;
  wire[27:0] MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_723_nl;
  wire[21:0] nl_MultLoop_acc_723_nl;
  wire[17:0] MultLoop_acc_693_nl;
  wire[18:0] nl_MultLoop_acc_693_nl;
  wire[27:0] MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_692_nl;
  wire[18:0] nl_MultLoop_acc_692_nl;
  wire[27:0] MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_691_nl;
  wire[18:0] nl_MultLoop_acc_691_nl;
  wire[27:0] MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_690_nl;
  wire[18:0] nl_MultLoop_acc_690_nl;
  wire[27:0] MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_689_nl;
  wire[18:0] nl_MultLoop_acc_689_nl;
  wire[27:0] MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_688_nl;
  wire[18:0] nl_MultLoop_acc_688_nl;
  wire[27:0] MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_687_nl;
  wire[18:0] nl_MultLoop_acc_687_nl;
  wire[27:0] MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_686_nl;
  wire[18:0] nl_MultLoop_acc_686_nl;
  wire[27:0] MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_681_nl;
  wire[18:0] nl_MultLoop_acc_681_nl;
  wire[27:0] MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_680_nl;
  wire[18:0] nl_MultLoop_acc_680_nl;
  wire[27:0] MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_679_nl;
  wire[18:0] nl_MultLoop_acc_679_nl;
  wire[27:0] MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_678_nl;
  wire[18:0] nl_MultLoop_acc_678_nl;
  wire[27:0] MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_685_nl;
  wire[18:0] nl_MultLoop_acc_685_nl;
  wire[27:0] MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_684_nl;
  wire[18:0] nl_MultLoop_acc_684_nl;
  wire[27:0] MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_683_nl;
  wire[18:0] nl_MultLoop_acc_683_nl;
  wire[27:0] MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_682_nl;
  wire[18:0] nl_MultLoop_acc_682_nl;
  wire[27:0] MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_722_nl;
  wire[20:0] nl_MultLoop_acc_722_nl;
  wire[17:0] MultLoop_acc_697_nl;
  wire[18:0] nl_MultLoop_acc_697_nl;
  wire[27:0] MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_696_nl;
  wire[18:0] nl_MultLoop_acc_696_nl;
  wire[27:0] MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_701_nl;
  wire[18:0] nl_MultLoop_acc_701_nl;
  wire[17:0] MultLoop_acc_677_nl;
  wire[18:0] nl_MultLoop_acc_677_nl;
  wire[27:0] MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_700_nl;
  wire[18:0] nl_MultLoop_acc_700_nl;
  wire[27:0] MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_699_nl;
  wire[18:0] nl_MultLoop_acc_699_nl;
  wire[27:0] MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_698_nl;
  wire[18:0] nl_MultLoop_acc_698_nl;
  wire[27:0] MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_695_nl;
  wire[18:0] nl_MultLoop_acc_695_nl;
  wire[27:0] MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[17:0] MultLoop_acc_694_nl;
  wire[18:0] nl_MultLoop_acc_694_nl;
  wire[27:0] MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire[27:0] MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;
  wire signed [35:0] nl_MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [431:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_431_414 , res_rsci_d_413_396 , res_rsci_d_395_378
      , res_rsci_d_377_360 , res_rsci_d_359_342 , res_rsci_d_341_324 , res_rsci_d_323_306
      , res_rsci_d_305_288 , res_rsci_d_287_270 , res_rsci_d_269_252 , res_rsci_d_251_234
      , res_rsci_d_233_216 , res_rsci_d_215_198 , res_rsci_d_197_180 , res_rsci_d_179_162
      , res_rsci_d_161_144 , res_rsci_d_143_126 , res_rsci_d_125_108 , res_rsci_d_107_90
      , res_rsci_d_89_72 , res_rsci_d_71_54 , res_rsci_d_53_36 , res_rsci_d_35_18
      , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd864)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd2),
  .width(32'sd432)) res_rsci (
      .d(nl_res_rsci_d[431:0]),
      .z(res_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd20736)) weights_rsci (
      .dat(weights_rsc_dat),
      .idat(weights_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd432)) biases_rsci (
      .dat(biases_rsc_dat),
      .idat(biases_rsci_idat)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_431_414 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_413_396 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
      res_rsci_d_395_378 <= 18'b000000000000000000;
      res_rsci_d_53_36 <= 18'b000000000000000000;
      res_rsci_d_377_360 <= 18'b000000000000000000;
      res_rsci_d_71_54 <= 18'b000000000000000000;
      res_rsci_d_359_342 <= 18'b000000000000000000;
      res_rsci_d_89_72 <= 18'b000000000000000000;
      res_rsci_d_341_324 <= 18'b000000000000000000;
      res_rsci_d_107_90 <= 18'b000000000000000000;
      res_rsci_d_323_306 <= 18'b000000000000000000;
      res_rsci_d_125_108 <= 18'b000000000000000000;
      res_rsci_d_305_288 <= 18'b000000000000000000;
      res_rsci_d_143_126 <= 18'b000000000000000000;
      res_rsci_d_287_270 <= 18'b000000000000000000;
      res_rsci_d_161_144 <= 18'b000000000000000000;
      res_rsci_d_269_252 <= 18'b000000000000000000;
      res_rsci_d_179_162 <= 18'b000000000000000000;
      res_rsci_d_251_234 <= 18'b000000000000000000;
      res_rsci_d_197_180 <= 18'b000000000000000000;
      res_rsci_d_233_216 <= 18'b000000000000000000;
      res_rsci_d_215_198 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_431_414 <= nl_res_rsci_d_431_414[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_413_396 <= nl_res_rsci_d_413_396[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
      res_rsci_d_395_378 <= nl_res_rsci_d_395_378[17:0];
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
      res_rsci_d_377_360 <= nl_res_rsci_d_377_360[17:0];
      res_rsci_d_71_54 <= nl_res_rsci_d_71_54[17:0];
      res_rsci_d_359_342 <= nl_res_rsci_d_359_342[17:0];
      res_rsci_d_89_72 <= nl_res_rsci_d_89_72[17:0];
      res_rsci_d_341_324 <= nl_res_rsci_d_341_324[17:0];
      res_rsci_d_107_90 <= nl_res_rsci_d_107_90[17:0];
      res_rsci_d_323_306 <= nl_res_rsci_d_323_306[17:0];
      res_rsci_d_125_108 <= nl_res_rsci_d_125_108[17:0];
      res_rsci_d_305_288 <= nl_res_rsci_d_305_288[17:0];
      res_rsci_d_143_126 <= nl_res_rsci_d_143_126[17:0];
      res_rsci_d_287_270 <= nl_res_rsci_d_287_270[17:0];
      res_rsci_d_161_144 <= nl_res_rsci_d_161_144[17:0];
      res_rsci_d_269_252 <= nl_res_rsci_d_269_252[17:0];
      res_rsci_d_179_162 <= nl_res_rsci_d_179_162[17:0];
      res_rsci_d_251_234 <= nl_res_rsci_d_251_234[17:0];
      res_rsci_d_197_180 <= nl_res_rsci_d_197_180[17:0];
      res_rsci_d_233_216 <= nl_res_rsci_d_233_216[17:0];
      res_rsci_d_215_198 <= nl_res_rsci_d_215_198[17:0];
    end
  end
  assign nl_MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[20141:20124]));
  assign MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[20159:20142]));
  assign MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_129_nl = (readslicef_28_18_10((MultLoop_1119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_129_nl = nl_MultLoop_acc_129_nl[17:0];
  assign nl_MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[20177:20160]));
  assign MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[20195:20178]));
  assign MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_128_nl = (readslicef_28_18_10((MultLoop_1121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_128_nl = nl_MultLoop_acc_128_nl[17:0];
  assign nl_MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[20213:20196]));
  assign MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[20231:20214]));
  assign MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_127_nl = (readslicef_28_18_10((MultLoop_1123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_127_nl = nl_MultLoop_acc_127_nl[17:0];
  assign nl_MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[20249:20232]));
  assign MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[20267:20250]));
  assign MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_126_nl = (readslicef_28_18_10((MultLoop_1125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_126_nl = nl_MultLoop_acc_126_nl[17:0];
  assign nl_MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[20285:20268]));
  assign MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[20303:20286]));
  assign MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_125_nl = (readslicef_28_18_10((MultLoop_1127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_125_nl = nl_MultLoop_acc_125_nl[17:0];
  assign nl_MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[20321:20304]));
  assign MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[20339:20322]));
  assign MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_124_nl = (readslicef_28_18_10((MultLoop_1129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_124_nl = nl_MultLoop_acc_124_nl[17:0];
  assign nl_MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[20357:20340]));
  assign MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[20375:20358]));
  assign MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_123_nl = (readslicef_28_18_10((MultLoop_1131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_123_nl = nl_MultLoop_acc_123_nl[17:0];
  assign nl_MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[20393:20376]));
  assign MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[20411:20394]));
  assign MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_122_nl = (readslicef_28_18_10((MultLoop_1133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_122_nl = nl_MultLoop_acc_122_nl[17:0];
  assign nl_MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[20573:20556]));
  assign MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[20591:20574]));
  assign MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_117_nl = (readslicef_28_18_10((MultLoop_1143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_117_nl = nl_MultLoop_acc_117_nl[17:0];
  assign nl_MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[20609:20592]));
  assign MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[20627:20610]));
  assign MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_116_nl = (readslicef_28_18_10((MultLoop_1145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_116_nl = nl_MultLoop_acc_116_nl[17:0];
  assign nl_MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[20645:20628]));
  assign MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[20663:20646]));
  assign MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_115_nl = (readslicef_28_18_10((MultLoop_1147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_115_nl = nl_MultLoop_acc_115_nl[17:0];
  assign nl_MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[20681:20664]));
  assign MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[20699:20682]));
  assign MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_114_nl = (readslicef_28_18_10((MultLoop_1149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_114_nl = nl_MultLoop_acc_114_nl[17:0];
  assign nl_MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[20429:20412]));
  assign MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[20447:20430]));
  assign MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_121_nl = (readslicef_28_18_10((MultLoop_1135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_121_nl = nl_MultLoop_acc_121_nl[17:0];
  assign nl_MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[20465:20448]));
  assign MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[20483:20466]));
  assign MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_120_nl = (readslicef_28_18_10((MultLoop_1137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_120_nl = nl_MultLoop_acc_120_nl[17:0];
  assign nl_MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[20501:20484]));
  assign MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[20519:20502]));
  assign MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_119_nl = (readslicef_28_18_10((MultLoop_1139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_119_nl = nl_MultLoop_acc_119_nl[17:0];
  assign nl_MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[20537:20520]));
  assign MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[20555:20538]));
  assign MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_118_nl = (readslicef_28_18_10((MultLoop_1141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_118_nl = nl_MultLoop_acc_118_nl[17:0];
  assign nl_MultLoop_acc_159_nl = (MultLoop_acc_129_nl) + (MultLoop_acc_128_nl) +
      (MultLoop_acc_127_nl) + (MultLoop_acc_126_nl) + (MultLoop_acc_125_nl) + (MultLoop_acc_124_nl)
      + (MultLoop_acc_123_nl) + (MultLoop_acc_122_nl) + (MultLoop_acc_117_nl) + (MultLoop_acc_116_nl)
      + (MultLoop_acc_115_nl) + (MultLoop_acc_114_nl) + (MultLoop_acc_121_nl) + (MultLoop_acc_120_nl)
      + (MultLoop_acc_119_nl) + (MultLoop_acc_118_nl);
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[17:0];
  assign nl_MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[19997:19980]));
  assign MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[20015:19998]));
  assign MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_133_nl = (readslicef_28_18_10((MultLoop_1111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[17:0];
  assign nl_MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[20033:20016]));
  assign MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[20051:20034]));
  assign MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_132_nl = (readslicef_28_18_10((MultLoop_1113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_132_nl = nl_MultLoop_acc_132_nl[17:0];
  assign nl_MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[20717:20700]));
  assign MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[20735:20718]));
  assign MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_113_nl = (readslicef_28_18_10((MultLoop_1151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_113_nl = nl_MultLoop_acc_113_nl[17:0];
  assign nl_MultLoop_acc_137_nl = (MultLoop_acc_113_nl) + (biases_rsci_idat[431:414]);
  assign MultLoop_acc_137_nl = nl_MultLoop_acc_137_nl[17:0];
  assign nl_MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[19889:19872]));
  assign MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[19907:19890]));
  assign MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_136_nl = (readslicef_28_18_10((MultLoop_1105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_136_nl = nl_MultLoop_acc_136_nl[17:0];
  assign nl_MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[19925:19908]));
  assign MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[19943:19926]));
  assign MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_135_nl = (readslicef_28_18_10((MultLoop_1107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_135_nl = nl_MultLoop_acc_135_nl[17:0];
  assign nl_MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[19961:19944]));
  assign MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[19979:19962]));
  assign MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_134_nl = (readslicef_28_18_10((MultLoop_1109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[17:0];
  assign nl_MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[20069:20052]));
  assign MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[20087:20070]));
  assign MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_131_nl = (readslicef_28_18_10((MultLoop_1115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_131_nl = nl_MultLoop_acc_131_nl[17:0];
  assign nl_MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[20105:20088]));
  assign MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[20123:20106]));
  assign MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_130_nl = (readslicef_28_18_10((MultLoop_1117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_130_nl = nl_MultLoop_acc_130_nl[17:0];
  assign nl_MultLoop_acc_158_nl = (MultLoop_acc_133_nl) + (MultLoop_acc_132_nl) +
      (MultLoop_acc_137_nl) + (MultLoop_acc_136_nl) + (MultLoop_acc_135_nl) + (MultLoop_acc_134_nl)
      + (MultLoop_acc_131_nl) + (MultLoop_acc_130_nl);
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[17:0];
  assign nl_res_rsci_d_431_414  = (MultLoop_acc_159_nl) + (MultLoop_acc_158_nl);
  assign nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[269:252]));
  assign MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[287:270]));
  assign MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1210_nl = (readslicef_28_18_10((MultLoop_15_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_16_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1210_nl = nl_MultLoop_acc_1210_nl[17:0];
  assign nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[305:288]));
  assign MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[323:306]));
  assign MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1209_nl = (readslicef_28_18_10((MultLoop_17_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_18_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1209_nl = nl_MultLoop_acc_1209_nl[17:0];
  assign nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[341:324]));
  assign MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[359:342]));
  assign MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1208_nl = (readslicef_28_18_10((MultLoop_19_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_20_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1208_nl = nl_MultLoop_acc_1208_nl[17:0];
  assign nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[377:360]));
  assign MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[395:378]));
  assign MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1207_nl = (readslicef_28_18_10((MultLoop_21_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_22_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1207_nl = nl_MultLoop_acc_1207_nl[17:0];
  assign nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[413:396]));
  assign MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[431:414]));
  assign MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1206_nl = (readslicef_28_18_10((MultLoop_23_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_24_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1206_nl = nl_MultLoop_acc_1206_nl[17:0];
  assign nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[449:432]));
  assign MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[467:450]));
  assign MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1205_nl = (readslicef_28_18_10((MultLoop_25_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_26_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1205_nl = nl_MultLoop_acc_1205_nl[17:0];
  assign nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[485:468]));
  assign MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[503:486]));
  assign MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1204_nl = (readslicef_28_18_10((MultLoop_27_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_28_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1204_nl = nl_MultLoop_acc_1204_nl[17:0];
  assign nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[521:504]));
  assign MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[539:522]));
  assign MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1203_nl = (readslicef_28_18_10((MultLoop_29_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_30_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1203_nl = nl_MultLoop_acc_1203_nl[17:0];
  assign nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[701:684]));
  assign MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[719:702]));
  assign MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1198_nl = (readslicef_28_18_10((MultLoop_39_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_40_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1198_nl = nl_MultLoop_acc_1198_nl[17:0];
  assign nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[737:720]));
  assign MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[755:738]));
  assign MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1197_nl = (readslicef_28_18_10((MultLoop_41_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_42_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1197_nl = nl_MultLoop_acc_1197_nl[17:0];
  assign nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[773:756]));
  assign MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[791:774]));
  assign MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1196_nl = (readslicef_28_18_10((MultLoop_43_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_44_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1196_nl = nl_MultLoop_acc_1196_nl[17:0];
  assign nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[809:792]));
  assign MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[827:810]));
  assign MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1195_nl = (readslicef_28_18_10((MultLoop_45_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_46_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1195_nl = nl_MultLoop_acc_1195_nl[17:0];
  assign nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[557:540]));
  assign MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[575:558]));
  assign MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1202_nl = (readslicef_28_18_10((MultLoop_31_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_32_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1202_nl = nl_MultLoop_acc_1202_nl[17:0];
  assign nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[593:576]));
  assign MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[611:594]));
  assign MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1201_nl = (readslicef_28_18_10((MultLoop_33_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_34_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1201_nl = nl_MultLoop_acc_1201_nl[17:0];
  assign nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[629:612]));
  assign MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[647:630]));
  assign MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1200_nl = (readslicef_28_18_10((MultLoop_35_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_36_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1200_nl = nl_MultLoop_acc_1200_nl[17:0];
  assign nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[665:648]));
  assign MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[683:666]));
  assign MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1199_nl = (readslicef_28_18_10((MultLoop_37_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_38_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1199_nl = nl_MultLoop_acc_1199_nl[17:0];
  assign nl_MultLoop_acc_1240_nl = (MultLoop_acc_1210_nl) + (MultLoop_acc_1209_nl)
      + (MultLoop_acc_1208_nl) + (MultLoop_acc_1207_nl) + (MultLoop_acc_1206_nl)
      + (MultLoop_acc_1205_nl) + (MultLoop_acc_1204_nl) + (MultLoop_acc_1203_nl)
      + (MultLoop_acc_1198_nl) + (MultLoop_acc_1197_nl) + (MultLoop_acc_1196_nl)
      + (MultLoop_acc_1195_nl) + (MultLoop_acc_1202_nl) + (MultLoop_acc_1201_nl)
      + (MultLoop_acc_1200_nl) + (MultLoop_acc_1199_nl);
  assign MultLoop_acc_1240_nl = nl_MultLoop_acc_1240_nl[17:0];
  assign nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[125:108]));
  assign MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[143:126]));
  assign MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1214_nl = (readslicef_28_18_10((MultLoop_7_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_8_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1214_nl = nl_MultLoop_acc_1214_nl[17:0];
  assign nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[161:144]));
  assign MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[179:162]));
  assign MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1213_nl = (readslicef_28_18_10((MultLoop_9_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_10_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1213_nl = nl_MultLoop_acc_1213_nl[17:0];
  assign nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[845:828]));
  assign MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[863:846]));
  assign MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1194_nl = (readslicef_28_18_10((MultLoop_47_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_48_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1194_nl = nl_MultLoop_acc_1194_nl[17:0];
  assign nl_MultLoop_acc_1218_nl = (MultLoop_acc_1194_nl) + (biases_rsci_idat[17:0]);
  assign MultLoop_acc_1218_nl = nl_MultLoop_acc_1218_nl[17:0];
  assign nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[17:0]));
  assign MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[35:18]));
  assign MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1217_nl = (readslicef_28_18_10((MultLoop_1_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_2_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1217_nl = nl_MultLoop_acc_1217_nl[17:0];
  assign nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[53:36]));
  assign MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[71:54]));
  assign MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1216_nl = (readslicef_28_18_10((MultLoop_3_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_4_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1216_nl = nl_MultLoop_acc_1216_nl[17:0];
  assign nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[89:72]));
  assign MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[107:90]));
  assign MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1215_nl = (readslicef_28_18_10((MultLoop_5_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_6_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1215_nl = nl_MultLoop_acc_1215_nl[17:0];
  assign nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[197:180]));
  assign MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[215:198]));
  assign MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1212_nl = (readslicef_28_18_10((MultLoop_11_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_12_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1212_nl = nl_MultLoop_acc_1212_nl[17:0];
  assign nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[233:216]));
  assign MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[251:234]));
  assign MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1211_nl = (readslicef_28_18_10((MultLoop_13_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_14_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1211_nl = nl_MultLoop_acc_1211_nl[17:0];
  assign nl_MultLoop_acc_1239_nl = (MultLoop_acc_1214_nl) + (MultLoop_acc_1213_nl)
      + (MultLoop_acc_1218_nl) + (MultLoop_acc_1217_nl) + (MultLoop_acc_1216_nl)
      + (MultLoop_acc_1215_nl) + (MultLoop_acc_1212_nl) + (MultLoop_acc_1211_nl);
  assign MultLoop_acc_1239_nl = nl_MultLoop_acc_1239_nl[17:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_1240_nl) + (MultLoop_acc_1239_nl);
  assign nl_MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[19277:19260]));
  assign MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[19295:19278]));
  assign MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_176_nl = (readslicef_28_18_10((MultLoop_1071_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1072_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_176_nl = nl_MultLoop_acc_176_nl[17:0];
  assign nl_MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[19313:19296]));
  assign MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[19331:19314]));
  assign MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_175_nl = (readslicef_28_18_10((MultLoop_1073_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1074_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_175_nl = nl_MultLoop_acc_175_nl[17:0];
  assign nl_MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[19349:19332]));
  assign MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[19367:19350]));
  assign MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_174_nl = (readslicef_28_18_10((MultLoop_1075_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1076_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_174_nl = nl_MultLoop_acc_174_nl[17:0];
  assign nl_MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[19385:19368]));
  assign MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[19403:19386]));
  assign MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_173_nl = (readslicef_28_18_10((MultLoop_1077_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1078_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_173_nl = nl_MultLoop_acc_173_nl[17:0];
  assign nl_MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[19421:19404]));
  assign MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[19439:19422]));
  assign MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_172_nl = (readslicef_28_18_10((MultLoop_1079_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1080_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_172_nl = nl_MultLoop_acc_172_nl[17:0];
  assign nl_MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[19457:19440]));
  assign MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[19475:19458]));
  assign MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_171_nl = (readslicef_28_18_10((MultLoop_1081_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1082_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_171_nl = nl_MultLoop_acc_171_nl[17:0];
  assign nl_MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[19493:19476]));
  assign MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[19511:19494]));
  assign MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_170_nl = (readslicef_28_18_10((MultLoop_1083_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1084_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_170_nl = nl_MultLoop_acc_170_nl[17:0];
  assign nl_MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[19529:19512]));
  assign MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[19547:19530]));
  assign MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_169_nl = (readslicef_28_18_10((MultLoop_1085_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1086_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_169_nl = nl_MultLoop_acc_169_nl[17:0];
  assign nl_MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[19709:19692]));
  assign MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[19727:19710]));
  assign MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_164_nl = (readslicef_28_18_10((MultLoop_1095_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1096_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_164_nl = nl_MultLoop_acc_164_nl[17:0];
  assign nl_MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[19745:19728]));
  assign MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[19763:19746]));
  assign MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_163_nl = (readslicef_28_18_10((MultLoop_1097_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1098_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_163_nl = nl_MultLoop_acc_163_nl[17:0];
  assign nl_MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[19781:19764]));
  assign MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[19799:19782]));
  assign MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_162_nl = (readslicef_28_18_10((MultLoop_1099_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_162_nl = nl_MultLoop_acc_162_nl[17:0];
  assign nl_MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[19817:19800]));
  assign MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[19835:19818]));
  assign MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_161_nl = (readslicef_28_18_10((MultLoop_1101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_161_nl = nl_MultLoop_acc_161_nl[17:0];
  assign nl_MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[19565:19548]));
  assign MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[19583:19566]));
  assign MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_168_nl = (readslicef_28_18_10((MultLoop_1087_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1088_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_168_nl = nl_MultLoop_acc_168_nl[17:0];
  assign nl_MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[19601:19584]));
  assign MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[19619:19602]));
  assign MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_167_nl = (readslicef_28_18_10((MultLoop_1089_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1090_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_167_nl = nl_MultLoop_acc_167_nl[17:0];
  assign nl_MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[19637:19620]));
  assign MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[19655:19638]));
  assign MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_166_nl = (readslicef_28_18_10((MultLoop_1091_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1092_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_166_nl = nl_MultLoop_acc_166_nl[17:0];
  assign nl_MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[19673:19656]));
  assign MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[19691:19674]));
  assign MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_165_nl = (readslicef_28_18_10((MultLoop_1093_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1094_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[17:0];
  assign nl_MultLoop_acc_206_nl = (MultLoop_acc_176_nl) + (MultLoop_acc_175_nl) +
      (MultLoop_acc_174_nl) + (MultLoop_acc_173_nl) + (MultLoop_acc_172_nl) + (MultLoop_acc_171_nl)
      + (MultLoop_acc_170_nl) + (MultLoop_acc_169_nl) + (MultLoop_acc_164_nl) + (MultLoop_acc_163_nl)
      + (MultLoop_acc_162_nl) + (MultLoop_acc_161_nl) + (MultLoop_acc_168_nl) + (MultLoop_acc_167_nl)
      + (MultLoop_acc_166_nl) + (MultLoop_acc_165_nl);
  assign MultLoop_acc_206_nl = nl_MultLoop_acc_206_nl[17:0];
  assign nl_MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[19133:19116]));
  assign MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[19151:19134]));
  assign MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_180_nl = (readslicef_28_18_10((MultLoop_1063_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1064_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_180_nl = nl_MultLoop_acc_180_nl[17:0];
  assign nl_MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[19169:19152]));
  assign MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[19187:19170]));
  assign MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_179_nl = (readslicef_28_18_10((MultLoop_1065_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1066_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_179_nl = nl_MultLoop_acc_179_nl[17:0];
  assign nl_MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[19853:19836]));
  assign MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[19871:19854]));
  assign MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_160_nl = (readslicef_28_18_10((MultLoop_1103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_160_nl = nl_MultLoop_acc_160_nl[17:0];
  assign nl_MultLoop_acc_184_nl = (MultLoop_acc_160_nl) + (biases_rsci_idat[413:396]);
  assign MultLoop_acc_184_nl = nl_MultLoop_acc_184_nl[17:0];
  assign nl_MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[19025:19008]));
  assign MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[19043:19026]));
  assign MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_183_nl = (readslicef_28_18_10((MultLoop_1057_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1058_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_183_nl = nl_MultLoop_acc_183_nl[17:0];
  assign nl_MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[19061:19044]));
  assign MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[19079:19062]));
  assign MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_182_nl = (readslicef_28_18_10((MultLoop_1059_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1060_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_182_nl = nl_MultLoop_acc_182_nl[17:0];
  assign nl_MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[19097:19080]));
  assign MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[19115:19098]));
  assign MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_181_nl = (readslicef_28_18_10((MultLoop_1061_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1062_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_181_nl = nl_MultLoop_acc_181_nl[17:0];
  assign nl_MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[19205:19188]));
  assign MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[19223:19206]));
  assign MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_178_nl = (readslicef_28_18_10((MultLoop_1067_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1068_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_178_nl = nl_MultLoop_acc_178_nl[17:0];
  assign nl_MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[19241:19224]));
  assign MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[19259:19242]));
  assign MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_177_nl = (readslicef_28_18_10((MultLoop_1069_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1070_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_177_nl = nl_MultLoop_acc_177_nl[17:0];
  assign nl_MultLoop_acc_205_nl = (MultLoop_acc_180_nl) + (MultLoop_acc_179_nl) +
      (MultLoop_acc_184_nl) + (MultLoop_acc_183_nl) + (MultLoop_acc_182_nl) + (MultLoop_acc_181_nl)
      + (MultLoop_acc_178_nl) + (MultLoop_acc_177_nl);
  assign MultLoop_acc_205_nl = nl_MultLoop_acc_205_nl[17:0];
  assign nl_res_rsci_d_413_396  = (MultLoop_acc_206_nl) + (MultLoop_acc_205_nl);
  assign nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[1133:1116]));
  assign MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[1151:1134]));
  assign MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1163_nl = (readslicef_28_18_10((MultLoop_63_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_64_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1163_nl = nl_MultLoop_acc_1163_nl[17:0];
  assign nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[1169:1152]));
  assign MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[1187:1170]));
  assign MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1162_nl = (readslicef_28_18_10((MultLoop_65_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_66_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1162_nl = nl_MultLoop_acc_1162_nl[17:0];
  assign nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[1205:1188]));
  assign MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[1223:1206]));
  assign MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1161_nl = (readslicef_28_18_10((MultLoop_67_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_68_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1161_nl = nl_MultLoop_acc_1161_nl[17:0];
  assign nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[1241:1224]));
  assign MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[1259:1242]));
  assign MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1160_nl = (readslicef_28_18_10((MultLoop_69_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_70_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1160_nl = nl_MultLoop_acc_1160_nl[17:0];
  assign nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[1277:1260]));
  assign MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[1295:1278]));
  assign MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1159_nl = (readslicef_28_18_10((MultLoop_71_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_72_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1159_nl = nl_MultLoop_acc_1159_nl[17:0];
  assign nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[1313:1296]));
  assign MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[1331:1314]));
  assign MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1158_nl = (readslicef_28_18_10((MultLoop_73_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_74_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1158_nl = nl_MultLoop_acc_1158_nl[17:0];
  assign nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[1349:1332]));
  assign MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[1367:1350]));
  assign MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1157_nl = (readslicef_28_18_10((MultLoop_75_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_76_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1157_nl = nl_MultLoop_acc_1157_nl[17:0];
  assign nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[1385:1368]));
  assign MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[1403:1386]));
  assign MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1156_nl = (readslicef_28_18_10((MultLoop_77_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_78_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1156_nl = nl_MultLoop_acc_1156_nl[17:0];
  assign nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[1565:1548]));
  assign MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[1583:1566]));
  assign MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1151_nl = (readslicef_28_18_10((MultLoop_87_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_88_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1151_nl = nl_MultLoop_acc_1151_nl[17:0];
  assign nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[1601:1584]));
  assign MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[1619:1602]));
  assign MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1150_nl = (readslicef_28_18_10((MultLoop_89_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_90_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1150_nl = nl_MultLoop_acc_1150_nl[17:0];
  assign nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[1637:1620]));
  assign MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[1655:1638]));
  assign MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1149_nl = (readslicef_28_18_10((MultLoop_91_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_92_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1149_nl = nl_MultLoop_acc_1149_nl[17:0];
  assign nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[1673:1656]));
  assign MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[1691:1674]));
  assign MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1148_nl = (readslicef_28_18_10((MultLoop_93_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_94_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1148_nl = nl_MultLoop_acc_1148_nl[17:0];
  assign nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[1421:1404]));
  assign MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[1439:1422]));
  assign MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1155_nl = (readslicef_28_18_10((MultLoop_79_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_80_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1155_nl = nl_MultLoop_acc_1155_nl[17:0];
  assign nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[1457:1440]));
  assign MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[1475:1458]));
  assign MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1154_nl = (readslicef_28_18_10((MultLoop_81_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_82_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1154_nl = nl_MultLoop_acc_1154_nl[17:0];
  assign nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[1493:1476]));
  assign MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[1511:1494]));
  assign MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1153_nl = (readslicef_28_18_10((MultLoop_83_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_84_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1153_nl = nl_MultLoop_acc_1153_nl[17:0];
  assign nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[1529:1512]));
  assign MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[1547:1530]));
  assign MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1152_nl = (readslicef_28_18_10((MultLoop_85_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_86_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1152_nl = nl_MultLoop_acc_1152_nl[17:0];
  assign nl_MultLoop_acc_1193_nl = (MultLoop_acc_1163_nl) + (MultLoop_acc_1162_nl)
      + (MultLoop_acc_1161_nl) + (MultLoop_acc_1160_nl) + (MultLoop_acc_1159_nl)
      + (MultLoop_acc_1158_nl) + (MultLoop_acc_1157_nl) + (MultLoop_acc_1156_nl)
      + (MultLoop_acc_1151_nl) + (MultLoop_acc_1150_nl) + (MultLoop_acc_1149_nl)
      + (MultLoop_acc_1148_nl) + (MultLoop_acc_1155_nl) + (MultLoop_acc_1154_nl)
      + (MultLoop_acc_1153_nl) + (MultLoop_acc_1152_nl);
  assign MultLoop_acc_1193_nl = nl_MultLoop_acc_1193_nl[17:0];
  assign nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[989:972]));
  assign MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[1007:990]));
  assign MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1167_nl = (readslicef_28_18_10((MultLoop_55_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_56_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1167_nl = nl_MultLoop_acc_1167_nl[17:0];
  assign nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[1025:1008]));
  assign MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[1043:1026]));
  assign MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1166_nl = (readslicef_28_18_10((MultLoop_57_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_58_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1166_nl = nl_MultLoop_acc_1166_nl[17:0];
  assign nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[1709:1692]));
  assign MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[1727:1710]));
  assign MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1147_nl = (readslicef_28_18_10((MultLoop_95_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_96_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1147_nl = nl_MultLoop_acc_1147_nl[17:0];
  assign nl_MultLoop_acc_1171_nl = (MultLoop_acc_1147_nl) + (biases_rsci_idat[35:18]);
  assign MultLoop_acc_1171_nl = nl_MultLoop_acc_1171_nl[17:0];
  assign nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[881:864]));
  assign MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[899:882]));
  assign MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1170_nl = (readslicef_28_18_10((MultLoop_49_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_50_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1170_nl = nl_MultLoop_acc_1170_nl[17:0];
  assign nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[917:900]));
  assign MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[935:918]));
  assign MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1169_nl = (readslicef_28_18_10((MultLoop_51_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_52_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1169_nl = nl_MultLoop_acc_1169_nl[17:0];
  assign nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[953:936]));
  assign MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[971:954]));
  assign MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1168_nl = (readslicef_28_18_10((MultLoop_53_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_54_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1168_nl = nl_MultLoop_acc_1168_nl[17:0];
  assign nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[1061:1044]));
  assign MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[1079:1062]));
  assign MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1165_nl = (readslicef_28_18_10((MultLoop_59_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_60_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1165_nl = nl_MultLoop_acc_1165_nl[17:0];
  assign nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[1097:1080]));
  assign MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[1115:1098]));
  assign MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1164_nl = (readslicef_28_18_10((MultLoop_61_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_62_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1164_nl = nl_MultLoop_acc_1164_nl[17:0];
  assign nl_MultLoop_acc_1192_nl = (MultLoop_acc_1167_nl) + (MultLoop_acc_1166_nl)
      + (MultLoop_acc_1171_nl) + (MultLoop_acc_1170_nl) + (MultLoop_acc_1169_nl)
      + (MultLoop_acc_1168_nl) + (MultLoop_acc_1165_nl) + (MultLoop_acc_1164_nl);
  assign MultLoop_acc_1192_nl = nl_MultLoop_acc_1192_nl[17:0];
  assign nl_res_rsci_d_35_18  = (MultLoop_acc_1193_nl) + (MultLoop_acc_1192_nl);
  assign nl_MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[18413:18396]));
  assign MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[18431:18414]));
  assign MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_223_nl = (readslicef_28_18_10((MultLoop_1023_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1024_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_223_nl = nl_MultLoop_acc_223_nl[17:0];
  assign nl_MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[18449:18432]));
  assign MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[18467:18450]));
  assign MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_222_nl = (readslicef_28_18_10((MultLoop_1025_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1026_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_222_nl = nl_MultLoop_acc_222_nl[17:0];
  assign nl_MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[18485:18468]));
  assign MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[18503:18486]));
  assign MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_221_nl = (readslicef_28_18_10((MultLoop_1027_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1028_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_221_nl = nl_MultLoop_acc_221_nl[17:0];
  assign nl_MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[18521:18504]));
  assign MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[18539:18522]));
  assign MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_220_nl = (readslicef_28_18_10((MultLoop_1029_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1030_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_220_nl = nl_MultLoop_acc_220_nl[17:0];
  assign nl_MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[18557:18540]));
  assign MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[18575:18558]));
  assign MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_219_nl = (readslicef_28_18_10((MultLoop_1031_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1032_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_219_nl = nl_MultLoop_acc_219_nl[17:0];
  assign nl_MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[18593:18576]));
  assign MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[18611:18594]));
  assign MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_218_nl = (readslicef_28_18_10((MultLoop_1033_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1034_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_218_nl = nl_MultLoop_acc_218_nl[17:0];
  assign nl_MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[18629:18612]));
  assign MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[18647:18630]));
  assign MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_217_nl = (readslicef_28_18_10((MultLoop_1035_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1036_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_217_nl = nl_MultLoop_acc_217_nl[17:0];
  assign nl_MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[18665:18648]));
  assign MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[18683:18666]));
  assign MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_216_nl = (readslicef_28_18_10((MultLoop_1037_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1038_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_216_nl = nl_MultLoop_acc_216_nl[17:0];
  assign nl_MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[18845:18828]));
  assign MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[18863:18846]));
  assign MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_211_nl = (readslicef_28_18_10((MultLoop_1047_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1048_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_211_nl = nl_MultLoop_acc_211_nl[17:0];
  assign nl_MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[18881:18864]));
  assign MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[18899:18882]));
  assign MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_210_nl = (readslicef_28_18_10((MultLoop_1049_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1050_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_210_nl = nl_MultLoop_acc_210_nl[17:0];
  assign nl_MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[18917:18900]));
  assign MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[18935:18918]));
  assign MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_209_nl = (readslicef_28_18_10((MultLoop_1051_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1052_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_209_nl = nl_MultLoop_acc_209_nl[17:0];
  assign nl_MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[18953:18936]));
  assign MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[18971:18954]));
  assign MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_208_nl = (readslicef_28_18_10((MultLoop_1053_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1054_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_208_nl = nl_MultLoop_acc_208_nl[17:0];
  assign nl_MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[18701:18684]));
  assign MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[18719:18702]));
  assign MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_215_nl = (readslicef_28_18_10((MultLoop_1039_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1040_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_215_nl = nl_MultLoop_acc_215_nl[17:0];
  assign nl_MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[18737:18720]));
  assign MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[18755:18738]));
  assign MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_214_nl = (readslicef_28_18_10((MultLoop_1041_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1042_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_214_nl = nl_MultLoop_acc_214_nl[17:0];
  assign nl_MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[18773:18756]));
  assign MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[18791:18774]));
  assign MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_213_nl = (readslicef_28_18_10((MultLoop_1043_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1044_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_213_nl = nl_MultLoop_acc_213_nl[17:0];
  assign nl_MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[18809:18792]));
  assign MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[18827:18810]));
  assign MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_212_nl = (readslicef_28_18_10((MultLoop_1045_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1046_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_212_nl = nl_MultLoop_acc_212_nl[17:0];
  assign nl_MultLoop_acc_253_nl = (MultLoop_acc_223_nl) + (MultLoop_acc_222_nl) +
      (MultLoop_acc_221_nl) + (MultLoop_acc_220_nl) + (MultLoop_acc_219_nl) + (MultLoop_acc_218_nl)
      + (MultLoop_acc_217_nl) + (MultLoop_acc_216_nl) + (MultLoop_acc_211_nl) + (MultLoop_acc_210_nl)
      + (MultLoop_acc_209_nl) + (MultLoop_acc_208_nl) + (MultLoop_acc_215_nl) + (MultLoop_acc_214_nl)
      + (MultLoop_acc_213_nl) + (MultLoop_acc_212_nl);
  assign MultLoop_acc_253_nl = nl_MultLoop_acc_253_nl[17:0];
  assign nl_MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[18269:18252]));
  assign MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[18287:18270]));
  assign MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_227_nl = (readslicef_28_18_10((MultLoop_1015_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1016_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_227_nl = nl_MultLoop_acc_227_nl[17:0];
  assign nl_MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[18305:18288]));
  assign MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[18323:18306]));
  assign MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_226_nl = (readslicef_28_18_10((MultLoop_1017_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1018_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_226_nl = nl_MultLoop_acc_226_nl[17:0];
  assign nl_MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[18989:18972]));
  assign MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[19007:18990]));
  assign MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_207_nl = (readslicef_28_18_10((MultLoop_1055_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1056_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_207_nl = nl_MultLoop_acc_207_nl[17:0];
  assign nl_MultLoop_acc_231_nl = (MultLoop_acc_207_nl) + (biases_rsci_idat[395:378]);
  assign MultLoop_acc_231_nl = nl_MultLoop_acc_231_nl[17:0];
  assign nl_MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[18161:18144]));
  assign MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[18179:18162]));
  assign MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_230_nl = (readslicef_28_18_10((MultLoop_1009_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1010_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_230_nl = nl_MultLoop_acc_230_nl[17:0];
  assign nl_MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[18197:18180]));
  assign MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[18215:18198]));
  assign MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_229_nl = (readslicef_28_18_10((MultLoop_1011_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1012_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_229_nl = nl_MultLoop_acc_229_nl[17:0];
  assign nl_MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[18233:18216]));
  assign MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[18251:18234]));
  assign MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_228_nl = (readslicef_28_18_10((MultLoop_1013_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1014_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_228_nl = nl_MultLoop_acc_228_nl[17:0];
  assign nl_MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[18341:18324]));
  assign MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[18359:18342]));
  assign MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_225_nl = (readslicef_28_18_10((MultLoop_1019_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1020_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_225_nl = nl_MultLoop_acc_225_nl[17:0];
  assign nl_MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[18377:18360]));
  assign MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[18395:18378]));
  assign MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_224_nl = (readslicef_28_18_10((MultLoop_1021_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1022_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_224_nl = nl_MultLoop_acc_224_nl[17:0];
  assign nl_MultLoop_acc_252_nl = (MultLoop_acc_227_nl) + (MultLoop_acc_226_nl) +
      (MultLoop_acc_231_nl) + (MultLoop_acc_230_nl) + (MultLoop_acc_229_nl) + (MultLoop_acc_228_nl)
      + (MultLoop_acc_225_nl) + (MultLoop_acc_224_nl);
  assign MultLoop_acc_252_nl = nl_MultLoop_acc_252_nl[17:0];
  assign nl_res_rsci_d_395_378  = (MultLoop_acc_253_nl) + (MultLoop_acc_252_nl);
  assign nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[1997:1980]));
  assign MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[2015:1998]));
  assign MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1116_nl = (readslicef_28_18_10((MultLoop_111_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_112_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1116_nl = nl_MultLoop_acc_1116_nl[17:0];
  assign nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[2033:2016]));
  assign MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[2051:2034]));
  assign MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1115_nl = (readslicef_28_18_10((MultLoop_113_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_114_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1115_nl = nl_MultLoop_acc_1115_nl[17:0];
  assign nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[2069:2052]));
  assign MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[2087:2070]));
  assign MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1114_nl = (readslicef_28_18_10((MultLoop_115_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_116_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1114_nl = nl_MultLoop_acc_1114_nl[17:0];
  assign nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[2105:2088]));
  assign MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[2123:2106]));
  assign MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1113_nl = (readslicef_28_18_10((MultLoop_117_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_118_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1113_nl = nl_MultLoop_acc_1113_nl[17:0];
  assign nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[2141:2124]));
  assign MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[2159:2142]));
  assign MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1112_nl = (readslicef_28_18_10((MultLoop_119_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_120_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1112_nl = nl_MultLoop_acc_1112_nl[17:0];
  assign nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[2177:2160]));
  assign MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[2195:2178]));
  assign MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1111_nl = (readslicef_28_18_10((MultLoop_121_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_122_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1111_nl = nl_MultLoop_acc_1111_nl[17:0];
  assign nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[2213:2196]));
  assign MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[2231:2214]));
  assign MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1110_nl = (readslicef_28_18_10((MultLoop_123_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_124_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1110_nl = nl_MultLoop_acc_1110_nl[17:0];
  assign nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[2249:2232]));
  assign MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[2267:2250]));
  assign MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1109_nl = (readslicef_28_18_10((MultLoop_125_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_126_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1109_nl = nl_MultLoop_acc_1109_nl[17:0];
  assign nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[2429:2412]));
  assign MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[2447:2430]));
  assign MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1104_nl = (readslicef_28_18_10((MultLoop_135_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_136_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1104_nl = nl_MultLoop_acc_1104_nl[17:0];
  assign nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[2465:2448]));
  assign MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[2483:2466]));
  assign MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1103_nl = (readslicef_28_18_10((MultLoop_137_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_138_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1103_nl = nl_MultLoop_acc_1103_nl[17:0];
  assign nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[2501:2484]));
  assign MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[2519:2502]));
  assign MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1102_nl = (readslicef_28_18_10((MultLoop_139_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_140_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1102_nl = nl_MultLoop_acc_1102_nl[17:0];
  assign nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[2537:2520]));
  assign MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[2555:2538]));
  assign MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1101_nl = (readslicef_28_18_10((MultLoop_141_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_142_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1101_nl = nl_MultLoop_acc_1101_nl[17:0];
  assign nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[2285:2268]));
  assign MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[2303:2286]));
  assign MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1108_nl = (readslicef_28_18_10((MultLoop_127_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_128_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1108_nl = nl_MultLoop_acc_1108_nl[17:0];
  assign nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[2321:2304]));
  assign MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[2339:2322]));
  assign MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1107_nl = (readslicef_28_18_10((MultLoop_129_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_130_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1107_nl = nl_MultLoop_acc_1107_nl[17:0];
  assign nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[2357:2340]));
  assign MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[2375:2358]));
  assign MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1106_nl = (readslicef_28_18_10((MultLoop_131_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_132_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1106_nl = nl_MultLoop_acc_1106_nl[17:0];
  assign nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[2393:2376]));
  assign MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[2411:2394]));
  assign MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1105_nl = (readslicef_28_18_10((MultLoop_133_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_134_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1105_nl = nl_MultLoop_acc_1105_nl[17:0];
  assign nl_MultLoop_acc_1146_nl = (MultLoop_acc_1116_nl) + (MultLoop_acc_1115_nl)
      + (MultLoop_acc_1114_nl) + (MultLoop_acc_1113_nl) + (MultLoop_acc_1112_nl)
      + (MultLoop_acc_1111_nl) + (MultLoop_acc_1110_nl) + (MultLoop_acc_1109_nl)
      + (MultLoop_acc_1104_nl) + (MultLoop_acc_1103_nl) + (MultLoop_acc_1102_nl)
      + (MultLoop_acc_1101_nl) + (MultLoop_acc_1108_nl) + (MultLoop_acc_1107_nl)
      + (MultLoop_acc_1106_nl) + (MultLoop_acc_1105_nl);
  assign MultLoop_acc_1146_nl = nl_MultLoop_acc_1146_nl[17:0];
  assign nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[1853:1836]));
  assign MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[1871:1854]));
  assign MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1120_nl = (readslicef_28_18_10((MultLoop_103_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_104_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1120_nl = nl_MultLoop_acc_1120_nl[17:0];
  assign nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[1889:1872]));
  assign MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[1907:1890]));
  assign MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1119_nl = (readslicef_28_18_10((MultLoop_105_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_106_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1119_nl = nl_MultLoop_acc_1119_nl[17:0];
  assign nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[2573:2556]));
  assign MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[2591:2574]));
  assign MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1100_nl = (readslicef_28_18_10((MultLoop_143_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_144_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1100_nl = nl_MultLoop_acc_1100_nl[17:0];
  assign nl_MultLoop_acc_1124_nl = (MultLoop_acc_1100_nl) + (biases_rsci_idat[53:36]);
  assign MultLoop_acc_1124_nl = nl_MultLoop_acc_1124_nl[17:0];
  assign nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[1745:1728]));
  assign MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[1763:1746]));
  assign MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1123_nl = (readslicef_28_18_10((MultLoop_97_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_98_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1123_nl = nl_MultLoop_acc_1123_nl[17:0];
  assign nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[1781:1764]));
  assign MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[1799:1782]));
  assign MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1122_nl = (readslicef_28_18_10((MultLoop_99_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_100_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1122_nl = nl_MultLoop_acc_1122_nl[17:0];
  assign nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[1817:1800]));
  assign MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[1835:1818]));
  assign MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1121_nl = (readslicef_28_18_10((MultLoop_101_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_102_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1121_nl = nl_MultLoop_acc_1121_nl[17:0];
  assign nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[1925:1908]));
  assign MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[1943:1926]));
  assign MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1118_nl = (readslicef_28_18_10((MultLoop_107_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_108_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1118_nl = nl_MultLoop_acc_1118_nl[17:0];
  assign nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[1961:1944]));
  assign MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[1979:1962]));
  assign MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1117_nl = (readslicef_28_18_10((MultLoop_109_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_110_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1117_nl = nl_MultLoop_acc_1117_nl[17:0];
  assign nl_MultLoop_acc_1145_nl = (MultLoop_acc_1120_nl) + (MultLoop_acc_1119_nl)
      + (MultLoop_acc_1124_nl) + (MultLoop_acc_1123_nl) + (MultLoop_acc_1122_nl)
      + (MultLoop_acc_1121_nl) + (MultLoop_acc_1118_nl) + (MultLoop_acc_1117_nl);
  assign MultLoop_acc_1145_nl = nl_MultLoop_acc_1145_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_1146_nl) + (MultLoop_acc_1145_nl);
  assign nl_MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[17549:17532]));
  assign MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[17567:17550]));
  assign MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_270_nl = (readslicef_28_18_10((MultLoop_975_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_976_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[17:0];
  assign nl_MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[17585:17568]));
  assign MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[17603:17586]));
  assign MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_269_nl = (readslicef_28_18_10((MultLoop_977_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_978_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_269_nl = nl_MultLoop_acc_269_nl[17:0];
  assign nl_MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[17621:17604]));
  assign MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[17639:17622]));
  assign MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_268_nl = (readslicef_28_18_10((MultLoop_979_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_980_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_268_nl = nl_MultLoop_acc_268_nl[17:0];
  assign nl_MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[17657:17640]));
  assign MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[17675:17658]));
  assign MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_267_nl = (readslicef_28_18_10((MultLoop_981_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_982_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_267_nl = nl_MultLoop_acc_267_nl[17:0];
  assign nl_MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[17693:17676]));
  assign MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[17711:17694]));
  assign MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_266_nl = (readslicef_28_18_10((MultLoop_983_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_984_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_266_nl = nl_MultLoop_acc_266_nl[17:0];
  assign nl_MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[17729:17712]));
  assign MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[17747:17730]));
  assign MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_265_nl = (readslicef_28_18_10((MultLoop_985_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_986_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_265_nl = nl_MultLoop_acc_265_nl[17:0];
  assign nl_MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[17765:17748]));
  assign MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[17783:17766]));
  assign MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_264_nl = (readslicef_28_18_10((MultLoop_987_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_988_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_264_nl = nl_MultLoop_acc_264_nl[17:0];
  assign nl_MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[17801:17784]));
  assign MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[17819:17802]));
  assign MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_263_nl = (readslicef_28_18_10((MultLoop_989_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_990_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_263_nl = nl_MultLoop_acc_263_nl[17:0];
  assign nl_MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[17981:17964]));
  assign MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[17999:17982]));
  assign MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_258_nl = (readslicef_28_18_10((MultLoop_999_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1000_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_258_nl = nl_MultLoop_acc_258_nl[17:0];
  assign nl_MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[18017:18000]));
  assign MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[18035:18018]));
  assign MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_257_nl = (readslicef_28_18_10((MultLoop_1001_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1002_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_257_nl = nl_MultLoop_acc_257_nl[17:0];
  assign nl_MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[18053:18036]));
  assign MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[18071:18054]));
  assign MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_256_nl = (readslicef_28_18_10((MultLoop_1003_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1004_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_256_nl = nl_MultLoop_acc_256_nl[17:0];
  assign nl_MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[18089:18072]));
  assign MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[18107:18090]));
  assign MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_255_nl = (readslicef_28_18_10((MultLoop_1005_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1006_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_255_nl = nl_MultLoop_acc_255_nl[17:0];
  assign nl_MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[17837:17820]));
  assign MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[17855:17838]));
  assign MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_262_nl = (readslicef_28_18_10((MultLoop_991_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_992_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_262_nl = nl_MultLoop_acc_262_nl[17:0];
  assign nl_MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[17873:17856]));
  assign MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[17891:17874]));
  assign MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_261_nl = (readslicef_28_18_10((MultLoop_993_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_994_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_261_nl = nl_MultLoop_acc_261_nl[17:0];
  assign nl_MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[17909:17892]));
  assign MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[17927:17910]));
  assign MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_260_nl = (readslicef_28_18_10((MultLoop_995_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_996_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_260_nl = nl_MultLoop_acc_260_nl[17:0];
  assign nl_MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[17945:17928]));
  assign MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[17963:17946]));
  assign MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_259_nl = (readslicef_28_18_10((MultLoop_997_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_998_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_259_nl = nl_MultLoop_acc_259_nl[17:0];
  assign nl_MultLoop_acc_300_nl = (MultLoop_acc_270_nl) + (MultLoop_acc_269_nl) +
      (MultLoop_acc_268_nl) + (MultLoop_acc_267_nl) + (MultLoop_acc_266_nl) + (MultLoop_acc_265_nl)
      + (MultLoop_acc_264_nl) + (MultLoop_acc_263_nl) + (MultLoop_acc_258_nl) + (MultLoop_acc_257_nl)
      + (MultLoop_acc_256_nl) + (MultLoop_acc_255_nl) + (MultLoop_acc_262_nl) + (MultLoop_acc_261_nl)
      + (MultLoop_acc_260_nl) + (MultLoop_acc_259_nl);
  assign MultLoop_acc_300_nl = nl_MultLoop_acc_300_nl[17:0];
  assign nl_MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[17405:17388]));
  assign MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[17423:17406]));
  assign MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_274_nl = (readslicef_28_18_10((MultLoop_967_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_968_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_274_nl = nl_MultLoop_acc_274_nl[17:0];
  assign nl_MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[17441:17424]));
  assign MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[17459:17442]));
  assign MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_273_nl = (readslicef_28_18_10((MultLoop_969_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_970_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_273_nl = nl_MultLoop_acc_273_nl[17:0];
  assign nl_MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[18125:18108]));
  assign MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[18143:18126]));
  assign MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_254_nl = (readslicef_28_18_10((MultLoop_1007_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_1008_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_254_nl = nl_MultLoop_acc_254_nl[17:0];
  assign nl_MultLoop_acc_278_nl = (MultLoop_acc_254_nl) + (biases_rsci_idat[377:360]);
  assign MultLoop_acc_278_nl = nl_MultLoop_acc_278_nl[17:0];
  assign nl_MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[17297:17280]));
  assign MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[17315:17298]));
  assign MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_277_nl = (readslicef_28_18_10((MultLoop_961_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_962_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_277_nl = nl_MultLoop_acc_277_nl[17:0];
  assign nl_MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[17333:17316]));
  assign MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[17351:17334]));
  assign MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_276_nl = (readslicef_28_18_10((MultLoop_963_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_964_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_276_nl = nl_MultLoop_acc_276_nl[17:0];
  assign nl_MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[17369:17352]));
  assign MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[17387:17370]));
  assign MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_275_nl = (readslicef_28_18_10((MultLoop_965_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_966_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_275_nl = nl_MultLoop_acc_275_nl[17:0];
  assign nl_MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[17477:17460]));
  assign MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[17495:17478]));
  assign MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_272_nl = (readslicef_28_18_10((MultLoop_971_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_972_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_272_nl = nl_MultLoop_acc_272_nl[17:0];
  assign nl_MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[17513:17496]));
  assign MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[17531:17514]));
  assign MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_271_nl = (readslicef_28_18_10((MultLoop_973_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_974_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[17:0];
  assign nl_MultLoop_acc_299_nl = (MultLoop_acc_274_nl) + (MultLoop_acc_273_nl) +
      (MultLoop_acc_278_nl) + (MultLoop_acc_277_nl) + (MultLoop_acc_276_nl) + (MultLoop_acc_275_nl)
      + (MultLoop_acc_272_nl) + (MultLoop_acc_271_nl);
  assign MultLoop_acc_299_nl = nl_MultLoop_acc_299_nl[17:0];
  assign nl_res_rsci_d_377_360  = (MultLoop_acc_300_nl) + (MultLoop_acc_299_nl);
  assign nl_MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[2861:2844]));
  assign MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[2879:2862]));
  assign MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1069_nl = (readslicef_28_18_10((MultLoop_159_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_160_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1069_nl = nl_MultLoop_acc_1069_nl[17:0];
  assign nl_MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[2897:2880]));
  assign MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[2915:2898]));
  assign MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1068_nl = (readslicef_28_18_10((MultLoop_161_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_162_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1068_nl = nl_MultLoop_acc_1068_nl[17:0];
  assign nl_MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[2933:2916]));
  assign MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[2951:2934]));
  assign MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1067_nl = (readslicef_28_18_10((MultLoop_163_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_164_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1067_nl = nl_MultLoop_acc_1067_nl[17:0];
  assign nl_MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[2969:2952]));
  assign MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[2987:2970]));
  assign MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1066_nl = (readslicef_28_18_10((MultLoop_165_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_166_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1066_nl = nl_MultLoop_acc_1066_nl[17:0];
  assign nl_MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[3005:2988]));
  assign MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[3023:3006]));
  assign MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1065_nl = (readslicef_28_18_10((MultLoop_167_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_168_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1065_nl = nl_MultLoop_acc_1065_nl[17:0];
  assign nl_MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[3041:3024]));
  assign MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[3059:3042]));
  assign MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1064_nl = (readslicef_28_18_10((MultLoop_169_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_170_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1064_nl = nl_MultLoop_acc_1064_nl[17:0];
  assign nl_MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[3077:3060]));
  assign MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[3095:3078]));
  assign MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1063_nl = (readslicef_28_18_10((MultLoop_171_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_172_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1063_nl = nl_MultLoop_acc_1063_nl[17:0];
  assign nl_MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[3113:3096]));
  assign MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[3131:3114]));
  assign MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1062_nl = (readslicef_28_18_10((MultLoop_173_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_174_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1062_nl = nl_MultLoop_acc_1062_nl[17:0];
  assign nl_MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[3293:3276]));
  assign MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[3311:3294]));
  assign MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1057_nl = (readslicef_28_18_10((MultLoop_183_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_184_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1057_nl = nl_MultLoop_acc_1057_nl[17:0];
  assign nl_MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[3329:3312]));
  assign MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[3347:3330]));
  assign MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1056_nl = (readslicef_28_18_10((MultLoop_185_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_186_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1056_nl = nl_MultLoop_acc_1056_nl[17:0];
  assign nl_MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[3365:3348]));
  assign MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[3383:3366]));
  assign MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1055_nl = (readslicef_28_18_10((MultLoop_187_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_188_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1055_nl = nl_MultLoop_acc_1055_nl[17:0];
  assign nl_MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[3401:3384]));
  assign MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[3419:3402]));
  assign MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1054_nl = (readslicef_28_18_10((MultLoop_189_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_190_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1054_nl = nl_MultLoop_acc_1054_nl[17:0];
  assign nl_MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[3149:3132]));
  assign MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[3167:3150]));
  assign MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1061_nl = (readslicef_28_18_10((MultLoop_175_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_176_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1061_nl = nl_MultLoop_acc_1061_nl[17:0];
  assign nl_MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[3185:3168]));
  assign MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[3203:3186]));
  assign MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1060_nl = (readslicef_28_18_10((MultLoop_177_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_178_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1060_nl = nl_MultLoop_acc_1060_nl[17:0];
  assign nl_MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[3221:3204]));
  assign MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[3239:3222]));
  assign MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1059_nl = (readslicef_28_18_10((MultLoop_179_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_180_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1059_nl = nl_MultLoop_acc_1059_nl[17:0];
  assign nl_MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[3257:3240]));
  assign MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[3275:3258]));
  assign MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1058_nl = (readslicef_28_18_10((MultLoop_181_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_182_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1058_nl = nl_MultLoop_acc_1058_nl[17:0];
  assign nl_MultLoop_acc_1099_nl = (MultLoop_acc_1069_nl) + (MultLoop_acc_1068_nl)
      + (MultLoop_acc_1067_nl) + (MultLoop_acc_1066_nl) + (MultLoop_acc_1065_nl)
      + (MultLoop_acc_1064_nl) + (MultLoop_acc_1063_nl) + (MultLoop_acc_1062_nl)
      + (MultLoop_acc_1057_nl) + (MultLoop_acc_1056_nl) + (MultLoop_acc_1055_nl)
      + (MultLoop_acc_1054_nl) + (MultLoop_acc_1061_nl) + (MultLoop_acc_1060_nl)
      + (MultLoop_acc_1059_nl) + (MultLoop_acc_1058_nl);
  assign MultLoop_acc_1099_nl = nl_MultLoop_acc_1099_nl[17:0];
  assign nl_MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[2717:2700]));
  assign MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[2735:2718]));
  assign MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1073_nl = (readslicef_28_18_10((MultLoop_151_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_152_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1073_nl = nl_MultLoop_acc_1073_nl[17:0];
  assign nl_MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[2753:2736]));
  assign MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[2771:2754]));
  assign MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1072_nl = (readslicef_28_18_10((MultLoop_153_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_154_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1072_nl = nl_MultLoop_acc_1072_nl[17:0];
  assign nl_MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[3437:3420]));
  assign MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[3455:3438]));
  assign MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1053_nl = (readslicef_28_18_10((MultLoop_191_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_192_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1053_nl = nl_MultLoop_acc_1053_nl[17:0];
  assign nl_MultLoop_acc_1077_nl = (MultLoop_acc_1053_nl) + (biases_rsci_idat[71:54]);
  assign MultLoop_acc_1077_nl = nl_MultLoop_acc_1077_nl[17:0];
  assign nl_MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[2609:2592]));
  assign MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[2627:2610]));
  assign MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1076_nl = (readslicef_28_18_10((MultLoop_145_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_146_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1076_nl = nl_MultLoop_acc_1076_nl[17:0];
  assign nl_MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[2645:2628]));
  assign MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[2663:2646]));
  assign MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1075_nl = (readslicef_28_18_10((MultLoop_147_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_148_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1075_nl = nl_MultLoop_acc_1075_nl[17:0];
  assign nl_MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[2681:2664]));
  assign MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[2699:2682]));
  assign MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1074_nl = (readslicef_28_18_10((MultLoop_149_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_150_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1074_nl = nl_MultLoop_acc_1074_nl[17:0];
  assign nl_MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[2789:2772]));
  assign MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[2807:2790]));
  assign MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1071_nl = (readslicef_28_18_10((MultLoop_155_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_156_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1071_nl = nl_MultLoop_acc_1071_nl[17:0];
  assign nl_MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[2825:2808]));
  assign MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[2843:2826]));
  assign MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1070_nl = (readslicef_28_18_10((MultLoop_157_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_158_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1070_nl = nl_MultLoop_acc_1070_nl[17:0];
  assign nl_MultLoop_acc_1098_nl = (MultLoop_acc_1073_nl) + (MultLoop_acc_1072_nl)
      + (MultLoop_acc_1077_nl) + (MultLoop_acc_1076_nl) + (MultLoop_acc_1075_nl)
      + (MultLoop_acc_1074_nl) + (MultLoop_acc_1071_nl) + (MultLoop_acc_1070_nl);
  assign MultLoop_acc_1098_nl = nl_MultLoop_acc_1098_nl[17:0];
  assign nl_res_rsci_d_71_54  = (MultLoop_acc_1099_nl) + (MultLoop_acc_1098_nl);
  assign nl_MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[16685:16668]));
  assign MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[16703:16686]));
  assign MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_317_nl = (readslicef_28_18_10((MultLoop_927_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_928_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_317_nl = nl_MultLoop_acc_317_nl[17:0];
  assign nl_MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[16721:16704]));
  assign MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[16739:16722]));
  assign MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_316_nl = (readslicef_28_18_10((MultLoop_929_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_930_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_316_nl = nl_MultLoop_acc_316_nl[17:0];
  assign nl_MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[16757:16740]));
  assign MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[16775:16758]));
  assign MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_315_nl = (readslicef_28_18_10((MultLoop_931_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_932_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_315_nl = nl_MultLoop_acc_315_nl[17:0];
  assign nl_MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[16793:16776]));
  assign MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[16811:16794]));
  assign MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_314_nl = (readslicef_28_18_10((MultLoop_933_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_934_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_314_nl = nl_MultLoop_acc_314_nl[17:0];
  assign nl_MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[16829:16812]));
  assign MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[16847:16830]));
  assign MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_313_nl = (readslicef_28_18_10((MultLoop_935_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_936_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_313_nl = nl_MultLoop_acc_313_nl[17:0];
  assign nl_MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[16865:16848]));
  assign MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[16883:16866]));
  assign MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_312_nl = (readslicef_28_18_10((MultLoop_937_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_938_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_312_nl = nl_MultLoop_acc_312_nl[17:0];
  assign nl_MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[16901:16884]));
  assign MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[16919:16902]));
  assign MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_311_nl = (readslicef_28_18_10((MultLoop_939_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_940_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_311_nl = nl_MultLoop_acc_311_nl[17:0];
  assign nl_MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[16937:16920]));
  assign MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[16955:16938]));
  assign MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_310_nl = (readslicef_28_18_10((MultLoop_941_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_942_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[17:0];
  assign nl_MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[17117:17100]));
  assign MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[17135:17118]));
  assign MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_305_nl = (readslicef_28_18_10((MultLoop_951_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_952_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_305_nl = nl_MultLoop_acc_305_nl[17:0];
  assign nl_MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[17153:17136]));
  assign MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[17171:17154]));
  assign MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_304_nl = (readslicef_28_18_10((MultLoop_953_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_954_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[17:0];
  assign nl_MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[17189:17172]));
  assign MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[17207:17190]));
  assign MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_303_nl = (readslicef_28_18_10((MultLoop_955_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_956_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_303_nl = nl_MultLoop_acc_303_nl[17:0];
  assign nl_MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[17225:17208]));
  assign MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[17243:17226]));
  assign MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_302_nl = (readslicef_28_18_10((MultLoop_957_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_958_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_302_nl = nl_MultLoop_acc_302_nl[17:0];
  assign nl_MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[16973:16956]));
  assign MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[16991:16974]));
  assign MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_309_nl = (readslicef_28_18_10((MultLoop_943_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_944_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_309_nl = nl_MultLoop_acc_309_nl[17:0];
  assign nl_MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[17009:16992]));
  assign MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[17027:17010]));
  assign MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_308_nl = (readslicef_28_18_10((MultLoop_945_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_946_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_308_nl = nl_MultLoop_acc_308_nl[17:0];
  assign nl_MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[17045:17028]));
  assign MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[17063:17046]));
  assign MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_307_nl = (readslicef_28_18_10((MultLoop_947_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_948_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[17:0];
  assign nl_MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[17081:17064]));
  assign MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[17099:17082]));
  assign MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_306_nl = (readslicef_28_18_10((MultLoop_949_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_950_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_306_nl = nl_MultLoop_acc_306_nl[17:0];
  assign nl_MultLoop_acc_347_nl = (MultLoop_acc_317_nl) + (MultLoop_acc_316_nl) +
      (MultLoop_acc_315_nl) + (MultLoop_acc_314_nl) + (MultLoop_acc_313_nl) + (MultLoop_acc_312_nl)
      + (MultLoop_acc_311_nl) + (MultLoop_acc_310_nl) + (MultLoop_acc_305_nl) + (MultLoop_acc_304_nl)
      + (MultLoop_acc_303_nl) + (MultLoop_acc_302_nl) + (MultLoop_acc_309_nl) + (MultLoop_acc_308_nl)
      + (MultLoop_acc_307_nl) + (MultLoop_acc_306_nl);
  assign MultLoop_acc_347_nl = nl_MultLoop_acc_347_nl[17:0];
  assign nl_MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[16541:16524]));
  assign MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[16559:16542]));
  assign MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_321_nl = (readslicef_28_18_10((MultLoop_919_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_920_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_321_nl = nl_MultLoop_acc_321_nl[17:0];
  assign nl_MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[16577:16560]));
  assign MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[16595:16578]));
  assign MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_320_nl = (readslicef_28_18_10((MultLoop_921_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_922_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_320_nl = nl_MultLoop_acc_320_nl[17:0];
  assign nl_MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[17261:17244]));
  assign MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[17279:17262]));
  assign MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_301_nl = (readslicef_28_18_10((MultLoop_959_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_960_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_301_nl = nl_MultLoop_acc_301_nl[17:0];
  assign nl_MultLoop_acc_325_nl = (MultLoop_acc_301_nl) + (biases_rsci_idat[359:342]);
  assign MultLoop_acc_325_nl = nl_MultLoop_acc_325_nl[17:0];
  assign nl_MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[16433:16416]));
  assign MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[16451:16434]));
  assign MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_324_nl = (readslicef_28_18_10((MultLoop_913_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_914_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_324_nl = nl_MultLoop_acc_324_nl[17:0];
  assign nl_MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[16469:16452]));
  assign MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[16487:16470]));
  assign MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_323_nl = (readslicef_28_18_10((MultLoop_915_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_916_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_323_nl = nl_MultLoop_acc_323_nl[17:0];
  assign nl_MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[16505:16488]));
  assign MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[16523:16506]));
  assign MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_322_nl = (readslicef_28_18_10((MultLoop_917_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_918_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_322_nl = nl_MultLoop_acc_322_nl[17:0];
  assign nl_MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[16613:16596]));
  assign MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[16631:16614]));
  assign MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_319_nl = (readslicef_28_18_10((MultLoop_923_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_924_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_319_nl = nl_MultLoop_acc_319_nl[17:0];
  assign nl_MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[16649:16632]));
  assign MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[16667:16650]));
  assign MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_318_nl = (readslicef_28_18_10((MultLoop_925_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_926_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_318_nl = nl_MultLoop_acc_318_nl[17:0];
  assign nl_MultLoop_acc_346_nl = (MultLoop_acc_321_nl) + (MultLoop_acc_320_nl) +
      (MultLoop_acc_325_nl) + (MultLoop_acc_324_nl) + (MultLoop_acc_323_nl) + (MultLoop_acc_322_nl)
      + (MultLoop_acc_319_nl) + (MultLoop_acc_318_nl);
  assign MultLoop_acc_346_nl = nl_MultLoop_acc_346_nl[17:0];
  assign nl_res_rsci_d_359_342  = (MultLoop_acc_347_nl) + (MultLoop_acc_346_nl);
  assign nl_MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[3725:3708]));
  assign MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[3743:3726]));
  assign MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1022_nl = (readslicef_28_18_10((MultLoop_207_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_208_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1022_nl = nl_MultLoop_acc_1022_nl[17:0];
  assign nl_MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[3761:3744]));
  assign MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[3779:3762]));
  assign MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1021_nl = (readslicef_28_18_10((MultLoop_209_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_210_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1021_nl = nl_MultLoop_acc_1021_nl[17:0];
  assign nl_MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[3797:3780]));
  assign MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[3815:3798]));
  assign MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1020_nl = (readslicef_28_18_10((MultLoop_211_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_212_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1020_nl = nl_MultLoop_acc_1020_nl[17:0];
  assign nl_MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[3833:3816]));
  assign MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[3851:3834]));
  assign MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1019_nl = (readslicef_28_18_10((MultLoop_213_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_214_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1019_nl = nl_MultLoop_acc_1019_nl[17:0];
  assign nl_MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[3869:3852]));
  assign MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[3887:3870]));
  assign MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1018_nl = (readslicef_28_18_10((MultLoop_215_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_216_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1018_nl = nl_MultLoop_acc_1018_nl[17:0];
  assign nl_MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[3905:3888]));
  assign MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[3923:3906]));
  assign MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1017_nl = (readslicef_28_18_10((MultLoop_217_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_218_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1017_nl = nl_MultLoop_acc_1017_nl[17:0];
  assign nl_MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[3941:3924]));
  assign MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[3959:3942]));
  assign MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1016_nl = (readslicef_28_18_10((MultLoop_219_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_220_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1016_nl = nl_MultLoop_acc_1016_nl[17:0];
  assign nl_MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[3977:3960]));
  assign MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[3995:3978]));
  assign MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1015_nl = (readslicef_28_18_10((MultLoop_221_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_222_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1015_nl = nl_MultLoop_acc_1015_nl[17:0];
  assign nl_MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[4157:4140]));
  assign MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[4175:4158]));
  assign MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1010_nl = (readslicef_28_18_10((MultLoop_231_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_232_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1010_nl = nl_MultLoop_acc_1010_nl[17:0];
  assign nl_MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[4193:4176]));
  assign MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[4211:4194]));
  assign MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1009_nl = (readslicef_28_18_10((MultLoop_233_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_234_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1009_nl = nl_MultLoop_acc_1009_nl[17:0];
  assign nl_MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[4229:4212]));
  assign MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[4247:4230]));
  assign MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1008_nl = (readslicef_28_18_10((MultLoop_235_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_236_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1008_nl = nl_MultLoop_acc_1008_nl[17:0];
  assign nl_MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[4265:4248]));
  assign MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[4283:4266]));
  assign MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1007_nl = (readslicef_28_18_10((MultLoop_237_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_238_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1007_nl = nl_MultLoop_acc_1007_nl[17:0];
  assign nl_MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[4013:3996]));
  assign MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[4031:4014]));
  assign MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1014_nl = (readslicef_28_18_10((MultLoop_223_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_224_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1014_nl = nl_MultLoop_acc_1014_nl[17:0];
  assign nl_MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[4049:4032]));
  assign MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[4067:4050]));
  assign MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1013_nl = (readslicef_28_18_10((MultLoop_225_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_226_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1013_nl = nl_MultLoop_acc_1013_nl[17:0];
  assign nl_MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[4085:4068]));
  assign MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[4103:4086]));
  assign MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1012_nl = (readslicef_28_18_10((MultLoop_227_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_228_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1012_nl = nl_MultLoop_acc_1012_nl[17:0];
  assign nl_MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[4121:4104]));
  assign MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[4139:4122]));
  assign MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1011_nl = (readslicef_28_18_10((MultLoop_229_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_230_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1011_nl = nl_MultLoop_acc_1011_nl[17:0];
  assign nl_MultLoop_acc_1052_nl = (MultLoop_acc_1022_nl) + (MultLoop_acc_1021_nl)
      + (MultLoop_acc_1020_nl) + (MultLoop_acc_1019_nl) + (MultLoop_acc_1018_nl)
      + (MultLoop_acc_1017_nl) + (MultLoop_acc_1016_nl) + (MultLoop_acc_1015_nl)
      + (MultLoop_acc_1010_nl) + (MultLoop_acc_1009_nl) + (MultLoop_acc_1008_nl)
      + (MultLoop_acc_1007_nl) + (MultLoop_acc_1014_nl) + (MultLoop_acc_1013_nl)
      + (MultLoop_acc_1012_nl) + (MultLoop_acc_1011_nl);
  assign MultLoop_acc_1052_nl = nl_MultLoop_acc_1052_nl[17:0];
  assign nl_MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[3581:3564]));
  assign MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[3599:3582]));
  assign MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1026_nl = (readslicef_28_18_10((MultLoop_199_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_200_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1026_nl = nl_MultLoop_acc_1026_nl[17:0];
  assign nl_MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[3617:3600]));
  assign MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[3635:3618]));
  assign MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1025_nl = (readslicef_28_18_10((MultLoop_201_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_202_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1025_nl = nl_MultLoop_acc_1025_nl[17:0];
  assign nl_MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[4301:4284]));
  assign MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[4319:4302]));
  assign MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1006_nl = (readslicef_28_18_10((MultLoop_239_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_240_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1006_nl = nl_MultLoop_acc_1006_nl[17:0];
  assign nl_MultLoop_acc_1030_nl = (MultLoop_acc_1006_nl) + (biases_rsci_idat[89:72]);
  assign MultLoop_acc_1030_nl = nl_MultLoop_acc_1030_nl[17:0];
  assign nl_MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[3473:3456]));
  assign MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[3491:3474]));
  assign MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1029_nl = (readslicef_28_18_10((MultLoop_193_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_194_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1029_nl = nl_MultLoop_acc_1029_nl[17:0];
  assign nl_MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[3509:3492]));
  assign MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[3527:3510]));
  assign MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1028_nl = (readslicef_28_18_10((MultLoop_195_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_196_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1028_nl = nl_MultLoop_acc_1028_nl[17:0];
  assign nl_MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[3545:3528]));
  assign MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[3563:3546]));
  assign MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1027_nl = (readslicef_28_18_10((MultLoop_197_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_198_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1027_nl = nl_MultLoop_acc_1027_nl[17:0];
  assign nl_MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[3653:3636]));
  assign MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[3671:3654]));
  assign MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1024_nl = (readslicef_28_18_10((MultLoop_203_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_204_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1024_nl = nl_MultLoop_acc_1024_nl[17:0];
  assign nl_MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[3689:3672]));
  assign MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[3707:3690]));
  assign MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_1023_nl = (readslicef_28_18_10((MultLoop_205_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_206_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_1023_nl = nl_MultLoop_acc_1023_nl[17:0];
  assign nl_MultLoop_acc_1051_nl = (MultLoop_acc_1026_nl) + (MultLoop_acc_1025_nl)
      + (MultLoop_acc_1030_nl) + (MultLoop_acc_1029_nl) + (MultLoop_acc_1028_nl)
      + (MultLoop_acc_1027_nl) + (MultLoop_acc_1024_nl) + (MultLoop_acc_1023_nl);
  assign MultLoop_acc_1051_nl = nl_MultLoop_acc_1051_nl[17:0];
  assign nl_res_rsci_d_89_72  = (MultLoop_acc_1052_nl) + (MultLoop_acc_1051_nl);
  assign nl_MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[15821:15804]));
  assign MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[15839:15822]));
  assign MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_364_nl = (readslicef_28_18_10((MultLoop_879_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_880_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_364_nl = nl_MultLoop_acc_364_nl[17:0];
  assign nl_MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[15857:15840]));
  assign MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[15875:15858]));
  assign MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_363_nl = (readslicef_28_18_10((MultLoop_881_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_882_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_363_nl = nl_MultLoop_acc_363_nl[17:0];
  assign nl_MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[15893:15876]));
  assign MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[15911:15894]));
  assign MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_362_nl = (readslicef_28_18_10((MultLoop_883_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_884_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_362_nl = nl_MultLoop_acc_362_nl[17:0];
  assign nl_MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[15929:15912]));
  assign MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[15947:15930]));
  assign MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_361_nl = (readslicef_28_18_10((MultLoop_885_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_886_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_361_nl = nl_MultLoop_acc_361_nl[17:0];
  assign nl_MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[15965:15948]));
  assign MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[15983:15966]));
  assign MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_360_nl = (readslicef_28_18_10((MultLoop_887_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_888_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_360_nl = nl_MultLoop_acc_360_nl[17:0];
  assign nl_MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[16001:15984]));
  assign MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[16019:16002]));
  assign MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_359_nl = (readslicef_28_18_10((MultLoop_889_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_890_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_359_nl = nl_MultLoop_acc_359_nl[17:0];
  assign nl_MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[16037:16020]));
  assign MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[16055:16038]));
  assign MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_358_nl = (readslicef_28_18_10((MultLoop_891_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_892_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_358_nl = nl_MultLoop_acc_358_nl[17:0];
  assign nl_MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[16073:16056]));
  assign MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[16091:16074]));
  assign MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_357_nl = (readslicef_28_18_10((MultLoop_893_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_894_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_357_nl = nl_MultLoop_acc_357_nl[17:0];
  assign nl_MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[16253:16236]));
  assign MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[16271:16254]));
  assign MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_352_nl = (readslicef_28_18_10((MultLoop_903_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_904_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_352_nl = nl_MultLoop_acc_352_nl[17:0];
  assign nl_MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[16289:16272]));
  assign MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[16307:16290]));
  assign MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_351_nl = (readslicef_28_18_10((MultLoop_905_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_906_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_351_nl = nl_MultLoop_acc_351_nl[17:0];
  assign nl_MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[16325:16308]));
  assign MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[16343:16326]));
  assign MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_350_nl = (readslicef_28_18_10((MultLoop_907_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_908_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_350_nl = nl_MultLoop_acc_350_nl[17:0];
  assign nl_MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[16361:16344]));
  assign MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[16379:16362]));
  assign MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_349_nl = (readslicef_28_18_10((MultLoop_909_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_910_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_349_nl = nl_MultLoop_acc_349_nl[17:0];
  assign nl_MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[16109:16092]));
  assign MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[16127:16110]));
  assign MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_356_nl = (readslicef_28_18_10((MultLoop_895_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_896_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_356_nl = nl_MultLoop_acc_356_nl[17:0];
  assign nl_MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[16145:16128]));
  assign MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[16163:16146]));
  assign MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_355_nl = (readslicef_28_18_10((MultLoop_897_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_898_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_355_nl = nl_MultLoop_acc_355_nl[17:0];
  assign nl_MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[16181:16164]));
  assign MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[16199:16182]));
  assign MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_354_nl = (readslicef_28_18_10((MultLoop_899_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_900_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_354_nl = nl_MultLoop_acc_354_nl[17:0];
  assign nl_MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[16217:16200]));
  assign MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[16235:16218]));
  assign MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_353_nl = (readslicef_28_18_10((MultLoop_901_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_902_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_353_nl = nl_MultLoop_acc_353_nl[17:0];
  assign nl_MultLoop_acc_394_nl = (MultLoop_acc_364_nl) + (MultLoop_acc_363_nl) +
      (MultLoop_acc_362_nl) + (MultLoop_acc_361_nl) + (MultLoop_acc_360_nl) + (MultLoop_acc_359_nl)
      + (MultLoop_acc_358_nl) + (MultLoop_acc_357_nl) + (MultLoop_acc_352_nl) + (MultLoop_acc_351_nl)
      + (MultLoop_acc_350_nl) + (MultLoop_acc_349_nl) + (MultLoop_acc_356_nl) + (MultLoop_acc_355_nl)
      + (MultLoop_acc_354_nl) + (MultLoop_acc_353_nl);
  assign MultLoop_acc_394_nl = nl_MultLoop_acc_394_nl[17:0];
  assign nl_MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[15677:15660]));
  assign MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[15695:15678]));
  assign MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_368_nl = (readslicef_28_18_10((MultLoop_871_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_872_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_368_nl = nl_MultLoop_acc_368_nl[17:0];
  assign nl_MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[15713:15696]));
  assign MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[15731:15714]));
  assign MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_367_nl = (readslicef_28_18_10((MultLoop_873_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_874_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_367_nl = nl_MultLoop_acc_367_nl[17:0];
  assign nl_MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[16397:16380]));
  assign MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[16415:16398]));
  assign MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_348_nl = (readslicef_28_18_10((MultLoop_911_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_912_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_348_nl = nl_MultLoop_acc_348_nl[17:0];
  assign nl_MultLoop_acc_372_nl = (MultLoop_acc_348_nl) + (biases_rsci_idat[341:324]);
  assign MultLoop_acc_372_nl = nl_MultLoop_acc_372_nl[17:0];
  assign nl_MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[15569:15552]));
  assign MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[15587:15570]));
  assign MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_371_nl = (readslicef_28_18_10((MultLoop_865_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_866_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_371_nl = nl_MultLoop_acc_371_nl[17:0];
  assign nl_MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[15605:15588]));
  assign MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[15623:15606]));
  assign MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_370_nl = (readslicef_28_18_10((MultLoop_867_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_868_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_370_nl = nl_MultLoop_acc_370_nl[17:0];
  assign nl_MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[15641:15624]));
  assign MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[15659:15642]));
  assign MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_369_nl = (readslicef_28_18_10((MultLoop_869_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_870_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_369_nl = nl_MultLoop_acc_369_nl[17:0];
  assign nl_MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[15749:15732]));
  assign MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[15767:15750]));
  assign MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_366_nl = (readslicef_28_18_10((MultLoop_875_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_876_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_366_nl = nl_MultLoop_acc_366_nl[17:0];
  assign nl_MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[15785:15768]));
  assign MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[15803:15786]));
  assign MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_365_nl = (readslicef_28_18_10((MultLoop_877_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_878_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_365_nl = nl_MultLoop_acc_365_nl[17:0];
  assign nl_MultLoop_acc_393_nl = (MultLoop_acc_368_nl) + (MultLoop_acc_367_nl) +
      (MultLoop_acc_372_nl) + (MultLoop_acc_371_nl) + (MultLoop_acc_370_nl) + (MultLoop_acc_369_nl)
      + (MultLoop_acc_366_nl) + (MultLoop_acc_365_nl);
  assign MultLoop_acc_393_nl = nl_MultLoop_acc_393_nl[17:0];
  assign nl_res_rsci_d_341_324  = (MultLoop_acc_394_nl) + (MultLoop_acc_393_nl);
  assign nl_MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[4589:4572]));
  assign MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[4607:4590]));
  assign MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_975_nl = (readslicef_28_18_10((MultLoop_255_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_256_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_975_nl = nl_MultLoop_acc_975_nl[17:0];
  assign nl_MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[4625:4608]));
  assign MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[4643:4626]));
  assign MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_974_nl = (readslicef_28_18_10((MultLoop_257_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_258_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_974_nl = nl_MultLoop_acc_974_nl[17:0];
  assign nl_MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[4661:4644]));
  assign MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[4679:4662]));
  assign MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_973_nl = (readslicef_28_18_10((MultLoop_259_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_260_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_973_nl = nl_MultLoop_acc_973_nl[17:0];
  assign nl_MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[4697:4680]));
  assign MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[4715:4698]));
  assign MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_972_nl = (readslicef_28_18_10((MultLoop_261_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_262_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_972_nl = nl_MultLoop_acc_972_nl[17:0];
  assign nl_MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[4733:4716]));
  assign MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[4751:4734]));
  assign MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_971_nl = (readslicef_28_18_10((MultLoop_263_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_264_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_971_nl = nl_MultLoop_acc_971_nl[17:0];
  assign nl_MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[4769:4752]));
  assign MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[4787:4770]));
  assign MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_970_nl = (readslicef_28_18_10((MultLoop_265_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_266_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_970_nl = nl_MultLoop_acc_970_nl[17:0];
  assign nl_MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[4805:4788]));
  assign MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[4823:4806]));
  assign MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_969_nl = (readslicef_28_18_10((MultLoop_267_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_268_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_969_nl = nl_MultLoop_acc_969_nl[17:0];
  assign nl_MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[4841:4824]));
  assign MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[4859:4842]));
  assign MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_968_nl = (readslicef_28_18_10((MultLoop_269_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_270_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_968_nl = nl_MultLoop_acc_968_nl[17:0];
  assign nl_MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[5021:5004]));
  assign MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[5039:5022]));
  assign MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_963_nl = (readslicef_28_18_10((MultLoop_279_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_280_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_963_nl = nl_MultLoop_acc_963_nl[17:0];
  assign nl_MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[5057:5040]));
  assign MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[5075:5058]));
  assign MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_962_nl = (readslicef_28_18_10((MultLoop_281_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_282_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_962_nl = nl_MultLoop_acc_962_nl[17:0];
  assign nl_MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[5093:5076]));
  assign MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[5111:5094]));
  assign MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_961_nl = (readslicef_28_18_10((MultLoop_283_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_284_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_961_nl = nl_MultLoop_acc_961_nl[17:0];
  assign nl_MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[5129:5112]));
  assign MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[5147:5130]));
  assign MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_960_nl = (readslicef_28_18_10((MultLoop_285_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_286_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_960_nl = nl_MultLoop_acc_960_nl[17:0];
  assign nl_MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[4877:4860]));
  assign MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[4895:4878]));
  assign MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_967_nl = (readslicef_28_18_10((MultLoop_271_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_272_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_967_nl = nl_MultLoop_acc_967_nl[17:0];
  assign nl_MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[4913:4896]));
  assign MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[4931:4914]));
  assign MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_966_nl = (readslicef_28_18_10((MultLoop_273_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_274_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_966_nl = nl_MultLoop_acc_966_nl[17:0];
  assign nl_MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[4949:4932]));
  assign MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[4967:4950]));
  assign MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_965_nl = (readslicef_28_18_10((MultLoop_275_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_276_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_965_nl = nl_MultLoop_acc_965_nl[17:0];
  assign nl_MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[4985:4968]));
  assign MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[5003:4986]));
  assign MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_964_nl = (readslicef_28_18_10((MultLoop_277_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_278_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_964_nl = nl_MultLoop_acc_964_nl[17:0];
  assign nl_MultLoop_acc_1005_nl = (MultLoop_acc_975_nl) + (MultLoop_acc_974_nl)
      + (MultLoop_acc_973_nl) + (MultLoop_acc_972_nl) + (MultLoop_acc_971_nl) + (MultLoop_acc_970_nl)
      + (MultLoop_acc_969_nl) + (MultLoop_acc_968_nl) + (MultLoop_acc_963_nl) + (MultLoop_acc_962_nl)
      + (MultLoop_acc_961_nl) + (MultLoop_acc_960_nl) + (MultLoop_acc_967_nl) + (MultLoop_acc_966_nl)
      + (MultLoop_acc_965_nl) + (MultLoop_acc_964_nl);
  assign MultLoop_acc_1005_nl = nl_MultLoop_acc_1005_nl[17:0];
  assign nl_MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[4445:4428]));
  assign MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[4463:4446]));
  assign MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_979_nl = (readslicef_28_18_10((MultLoop_247_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_248_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_979_nl = nl_MultLoop_acc_979_nl[17:0];
  assign nl_MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[4481:4464]));
  assign MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[4499:4482]));
  assign MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_978_nl = (readslicef_28_18_10((MultLoop_249_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_250_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_978_nl = nl_MultLoop_acc_978_nl[17:0];
  assign nl_MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[5165:5148]));
  assign MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[5183:5166]));
  assign MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_959_nl = (readslicef_28_18_10((MultLoop_287_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_288_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_959_nl = nl_MultLoop_acc_959_nl[17:0];
  assign nl_MultLoop_acc_983_nl = (MultLoop_acc_959_nl) + (biases_rsci_idat[107:90]);
  assign MultLoop_acc_983_nl = nl_MultLoop_acc_983_nl[17:0];
  assign nl_MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[4337:4320]));
  assign MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[4355:4338]));
  assign MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_982_nl = (readslicef_28_18_10((MultLoop_241_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_242_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_982_nl = nl_MultLoop_acc_982_nl[17:0];
  assign nl_MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[4373:4356]));
  assign MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[4391:4374]));
  assign MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_981_nl = (readslicef_28_18_10((MultLoop_243_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_244_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_981_nl = nl_MultLoop_acc_981_nl[17:0];
  assign nl_MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[4409:4392]));
  assign MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[4427:4410]));
  assign MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_980_nl = (readslicef_28_18_10((MultLoop_245_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_246_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_980_nl = nl_MultLoop_acc_980_nl[17:0];
  assign nl_MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[4517:4500]));
  assign MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[4535:4518]));
  assign MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_977_nl = (readslicef_28_18_10((MultLoop_251_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_252_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_977_nl = nl_MultLoop_acc_977_nl[17:0];
  assign nl_MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[4553:4536]));
  assign MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[4571:4554]));
  assign MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_976_nl = (readslicef_28_18_10((MultLoop_253_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_254_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_976_nl = nl_MultLoop_acc_976_nl[17:0];
  assign nl_MultLoop_acc_1004_nl = (MultLoop_acc_979_nl) + (MultLoop_acc_978_nl)
      + (MultLoop_acc_983_nl) + (MultLoop_acc_982_nl) + (MultLoop_acc_981_nl) + (MultLoop_acc_980_nl)
      + (MultLoop_acc_977_nl) + (MultLoop_acc_976_nl);
  assign MultLoop_acc_1004_nl = nl_MultLoop_acc_1004_nl[17:0];
  assign nl_res_rsci_d_107_90  = (MultLoop_acc_1005_nl) + (MultLoop_acc_1004_nl);
  assign nl_MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[14957:14940]));
  assign MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[14975:14958]));
  assign MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_411_nl = (readslicef_28_18_10((MultLoop_831_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_832_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_411_nl = nl_MultLoop_acc_411_nl[17:0];
  assign nl_MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[14993:14976]));
  assign MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[15011:14994]));
  assign MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_410_nl = (readslicef_28_18_10((MultLoop_833_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_834_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_410_nl = nl_MultLoop_acc_410_nl[17:0];
  assign nl_MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[15029:15012]));
  assign MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[15047:15030]));
  assign MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_409_nl = (readslicef_28_18_10((MultLoop_835_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_836_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_409_nl = nl_MultLoop_acc_409_nl[17:0];
  assign nl_MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[15065:15048]));
  assign MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[15083:15066]));
  assign MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_408_nl = (readslicef_28_18_10((MultLoop_837_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_838_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_408_nl = nl_MultLoop_acc_408_nl[17:0];
  assign nl_MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[15101:15084]));
  assign MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[15119:15102]));
  assign MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_407_nl = (readslicef_28_18_10((MultLoop_839_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_840_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_407_nl = nl_MultLoop_acc_407_nl[17:0];
  assign nl_MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[15137:15120]));
  assign MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[15155:15138]));
  assign MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_406_nl = (readslicef_28_18_10((MultLoop_841_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_842_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_406_nl = nl_MultLoop_acc_406_nl[17:0];
  assign nl_MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[15173:15156]));
  assign MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[15191:15174]));
  assign MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_405_nl = (readslicef_28_18_10((MultLoop_843_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_844_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_405_nl = nl_MultLoop_acc_405_nl[17:0];
  assign nl_MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[15209:15192]));
  assign MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[15227:15210]));
  assign MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_404_nl = (readslicef_28_18_10((MultLoop_845_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_846_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_404_nl = nl_MultLoop_acc_404_nl[17:0];
  assign nl_MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[15389:15372]));
  assign MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[15407:15390]));
  assign MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_399_nl = (readslicef_28_18_10((MultLoop_855_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_856_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_399_nl = nl_MultLoop_acc_399_nl[17:0];
  assign nl_MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[15425:15408]));
  assign MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[15443:15426]));
  assign MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_398_nl = (readslicef_28_18_10((MultLoop_857_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_858_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_398_nl = nl_MultLoop_acc_398_nl[17:0];
  assign nl_MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[15461:15444]));
  assign MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[15479:15462]));
  assign MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_397_nl = (readslicef_28_18_10((MultLoop_859_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_860_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_397_nl = nl_MultLoop_acc_397_nl[17:0];
  assign nl_MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[15497:15480]));
  assign MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[15515:15498]));
  assign MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_396_nl = (readslicef_28_18_10((MultLoop_861_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_862_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_396_nl = nl_MultLoop_acc_396_nl[17:0];
  assign nl_MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[15245:15228]));
  assign MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[15263:15246]));
  assign MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_403_nl = (readslicef_28_18_10((MultLoop_847_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_848_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_403_nl = nl_MultLoop_acc_403_nl[17:0];
  assign nl_MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[15281:15264]));
  assign MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[15299:15282]));
  assign MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_402_nl = (readslicef_28_18_10((MultLoop_849_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_850_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_402_nl = nl_MultLoop_acc_402_nl[17:0];
  assign nl_MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[15317:15300]));
  assign MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[15335:15318]));
  assign MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_401_nl = (readslicef_28_18_10((MultLoop_851_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_852_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_401_nl = nl_MultLoop_acc_401_nl[17:0];
  assign nl_MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[15353:15336]));
  assign MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[15371:15354]));
  assign MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_400_nl = (readslicef_28_18_10((MultLoop_853_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_854_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_400_nl = nl_MultLoop_acc_400_nl[17:0];
  assign nl_MultLoop_acc_441_nl = (MultLoop_acc_411_nl) + (MultLoop_acc_410_nl) +
      (MultLoop_acc_409_nl) + (MultLoop_acc_408_nl) + (MultLoop_acc_407_nl) + (MultLoop_acc_406_nl)
      + (MultLoop_acc_405_nl) + (MultLoop_acc_404_nl) + (MultLoop_acc_399_nl) + (MultLoop_acc_398_nl)
      + (MultLoop_acc_397_nl) + (MultLoop_acc_396_nl) + (MultLoop_acc_403_nl) + (MultLoop_acc_402_nl)
      + (MultLoop_acc_401_nl) + (MultLoop_acc_400_nl);
  assign MultLoop_acc_441_nl = nl_MultLoop_acc_441_nl[17:0];
  assign nl_MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[14813:14796]));
  assign MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[14831:14814]));
  assign MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_415_nl = (readslicef_28_18_10((MultLoop_823_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_824_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_415_nl = nl_MultLoop_acc_415_nl[17:0];
  assign nl_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[14849:14832]));
  assign MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[14867:14850]));
  assign MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_414_nl = (readslicef_28_18_10((MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_826_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_414_nl = nl_MultLoop_acc_414_nl[17:0];
  assign nl_MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[15533:15516]));
  assign MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[15551:15534]));
  assign MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_395_nl = (readslicef_28_18_10((MultLoop_863_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_864_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_395_nl = nl_MultLoop_acc_395_nl[17:0];
  assign nl_MultLoop_acc_419_nl = (MultLoop_acc_395_nl) + (biases_rsci_idat[323:306]);
  assign MultLoop_acc_419_nl = nl_MultLoop_acc_419_nl[17:0];
  assign nl_MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[14705:14688]));
  assign MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[14723:14706]));
  assign MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_418_nl = (readslicef_28_18_10((MultLoop_817_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_818_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_418_nl = nl_MultLoop_acc_418_nl[17:0];
  assign nl_MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[14741:14724]));
  assign MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[14759:14742]));
  assign MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_417_nl = (readslicef_28_18_10((MultLoop_819_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_820_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_417_nl = nl_MultLoop_acc_417_nl[17:0];
  assign nl_MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[14777:14760]));
  assign MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[14795:14778]));
  assign MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_416_nl = (readslicef_28_18_10((MultLoop_821_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_822_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_416_nl = nl_MultLoop_acc_416_nl[17:0];
  assign nl_MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[14885:14868]));
  assign MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[14903:14886]));
  assign MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_413_nl = (readslicef_28_18_10((MultLoop_827_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_828_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_413_nl = nl_MultLoop_acc_413_nl[17:0];
  assign nl_MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[14921:14904]));
  assign MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[14939:14922]));
  assign MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_412_nl = (readslicef_28_18_10((MultLoop_829_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_830_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_412_nl = nl_MultLoop_acc_412_nl[17:0];
  assign nl_MultLoop_acc_440_nl = (MultLoop_acc_415_nl) + (MultLoop_acc_414_nl) +
      (MultLoop_acc_419_nl) + (MultLoop_acc_418_nl) + (MultLoop_acc_417_nl) + (MultLoop_acc_416_nl)
      + (MultLoop_acc_413_nl) + (MultLoop_acc_412_nl);
  assign MultLoop_acc_440_nl = nl_MultLoop_acc_440_nl[17:0];
  assign nl_res_rsci_d_323_306  = (MultLoop_acc_441_nl) + (MultLoop_acc_440_nl);
  assign nl_MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[5453:5436]));
  assign MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[5471:5454]));
  assign MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_928_nl = (readslicef_28_18_10((MultLoop_303_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_304_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_928_nl = nl_MultLoop_acc_928_nl[17:0];
  assign nl_MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[5489:5472]));
  assign MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[5507:5490]));
  assign MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_927_nl = (readslicef_28_18_10((MultLoop_305_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_306_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_927_nl = nl_MultLoop_acc_927_nl[17:0];
  assign nl_MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[5525:5508]));
  assign MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[5543:5526]));
  assign MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_926_nl = (readslicef_28_18_10((MultLoop_307_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_308_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_926_nl = nl_MultLoop_acc_926_nl[17:0];
  assign nl_MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[5561:5544]));
  assign MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[5579:5562]));
  assign MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_925_nl = (readslicef_28_18_10((MultLoop_309_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_310_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_925_nl = nl_MultLoop_acc_925_nl[17:0];
  assign nl_MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[5597:5580]));
  assign MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[5615:5598]));
  assign MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_924_nl = (readslicef_28_18_10((MultLoop_311_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_312_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_924_nl = nl_MultLoop_acc_924_nl[17:0];
  assign nl_MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[5633:5616]));
  assign MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[5651:5634]));
  assign MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_923_nl = (readslicef_28_18_10((MultLoop_313_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_314_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_923_nl = nl_MultLoop_acc_923_nl[17:0];
  assign nl_MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[5669:5652]));
  assign MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[5687:5670]));
  assign MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_922_nl = (readslicef_28_18_10((MultLoop_315_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_316_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_922_nl = nl_MultLoop_acc_922_nl[17:0];
  assign nl_MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[5705:5688]));
  assign MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[5723:5706]));
  assign MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_921_nl = (readslicef_28_18_10((MultLoop_317_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_318_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_921_nl = nl_MultLoop_acc_921_nl[17:0];
  assign nl_MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[5885:5868]));
  assign MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[5903:5886]));
  assign MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_916_nl = (readslicef_28_18_10((MultLoop_327_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_328_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_916_nl = nl_MultLoop_acc_916_nl[17:0];
  assign nl_MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[5921:5904]));
  assign MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[5939:5922]));
  assign MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_915_nl = (readslicef_28_18_10((MultLoop_329_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_330_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_915_nl = nl_MultLoop_acc_915_nl[17:0];
  assign nl_MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[5957:5940]));
  assign MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[5975:5958]));
  assign MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_914_nl = (readslicef_28_18_10((MultLoop_331_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_332_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_914_nl = nl_MultLoop_acc_914_nl[17:0];
  assign nl_MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[5993:5976]));
  assign MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[6011:5994]));
  assign MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_913_nl = (readslicef_28_18_10((MultLoop_333_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_334_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_913_nl = nl_MultLoop_acc_913_nl[17:0];
  assign nl_MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[5741:5724]));
  assign MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[5759:5742]));
  assign MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_920_nl = (readslicef_28_18_10((MultLoop_319_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_320_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_920_nl = nl_MultLoop_acc_920_nl[17:0];
  assign nl_MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[5777:5760]));
  assign MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[5795:5778]));
  assign MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_919_nl = (readslicef_28_18_10((MultLoop_321_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_322_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_919_nl = nl_MultLoop_acc_919_nl[17:0];
  assign nl_MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[5813:5796]));
  assign MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[5831:5814]));
  assign MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_918_nl = (readslicef_28_18_10((MultLoop_323_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_324_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_918_nl = nl_MultLoop_acc_918_nl[17:0];
  assign nl_MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[5849:5832]));
  assign MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[5867:5850]));
  assign MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_917_nl = (readslicef_28_18_10((MultLoop_325_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_326_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_917_nl = nl_MultLoop_acc_917_nl[17:0];
  assign nl_MultLoop_acc_958_nl = (MultLoop_acc_928_nl) + (MultLoop_acc_927_nl) +
      (MultLoop_acc_926_nl) + (MultLoop_acc_925_nl) + (MultLoop_acc_924_nl) + (MultLoop_acc_923_nl)
      + (MultLoop_acc_922_nl) + (MultLoop_acc_921_nl) + (MultLoop_acc_916_nl) + (MultLoop_acc_915_nl)
      + (MultLoop_acc_914_nl) + (MultLoop_acc_913_nl) + (MultLoop_acc_920_nl) + (MultLoop_acc_919_nl)
      + (MultLoop_acc_918_nl) + (MultLoop_acc_917_nl);
  assign MultLoop_acc_958_nl = nl_MultLoop_acc_958_nl[17:0];
  assign nl_MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[5309:5292]));
  assign MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[5327:5310]));
  assign MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_932_nl = (readslicef_28_18_10((MultLoop_295_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_296_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_932_nl = nl_MultLoop_acc_932_nl[17:0];
  assign nl_MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[5345:5328]));
  assign MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[5363:5346]));
  assign MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_931_nl = (readslicef_28_18_10((MultLoop_297_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_298_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_931_nl = nl_MultLoop_acc_931_nl[17:0];
  assign nl_MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[6029:6012]));
  assign MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[6047:6030]));
  assign MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_912_nl = (readslicef_28_18_10((MultLoop_335_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_336_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_912_nl = nl_MultLoop_acc_912_nl[17:0];
  assign nl_MultLoop_acc_936_nl = (MultLoop_acc_912_nl) + (biases_rsci_idat[125:108]);
  assign MultLoop_acc_936_nl = nl_MultLoop_acc_936_nl[17:0];
  assign nl_MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[5201:5184]));
  assign MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[5219:5202]));
  assign MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_935_nl = (readslicef_28_18_10((MultLoop_289_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_290_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_935_nl = nl_MultLoop_acc_935_nl[17:0];
  assign nl_MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[5237:5220]));
  assign MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[5255:5238]));
  assign MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_934_nl = (readslicef_28_18_10((MultLoop_291_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_292_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_934_nl = nl_MultLoop_acc_934_nl[17:0];
  assign nl_MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[5273:5256]));
  assign MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[5291:5274]));
  assign MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_933_nl = (readslicef_28_18_10((MultLoop_293_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_294_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_933_nl = nl_MultLoop_acc_933_nl[17:0];
  assign nl_MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[5381:5364]));
  assign MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[5399:5382]));
  assign MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_930_nl = (readslicef_28_18_10((MultLoop_299_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_300_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_930_nl = nl_MultLoop_acc_930_nl[17:0];
  assign nl_MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[5417:5400]));
  assign MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[5435:5418]));
  assign MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_929_nl = (readslicef_28_18_10((MultLoop_301_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_302_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_929_nl = nl_MultLoop_acc_929_nl[17:0];
  assign nl_MultLoop_acc_957_nl = (MultLoop_acc_932_nl) + (MultLoop_acc_931_nl) +
      (MultLoop_acc_936_nl) + (MultLoop_acc_935_nl) + (MultLoop_acc_934_nl) + (MultLoop_acc_933_nl)
      + (MultLoop_acc_930_nl) + (MultLoop_acc_929_nl);
  assign MultLoop_acc_957_nl = nl_MultLoop_acc_957_nl[17:0];
  assign nl_res_rsci_d_125_108  = (MultLoop_acc_958_nl) + (MultLoop_acc_957_nl);
  assign nl_MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[14093:14076]));
  assign MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[14111:14094]));
  assign MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_458_nl = (readslicef_28_18_10((MultLoop_783_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_784_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_458_nl = nl_MultLoop_acc_458_nl[17:0];
  assign nl_MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[14129:14112]));
  assign MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[14147:14130]));
  assign MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_457_nl = (readslicef_28_18_10((MultLoop_785_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_786_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_457_nl = nl_MultLoop_acc_457_nl[17:0];
  assign nl_MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[14165:14148]));
  assign MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[14183:14166]));
  assign MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_456_nl = (readslicef_28_18_10((MultLoop_787_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_788_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_456_nl = nl_MultLoop_acc_456_nl[17:0];
  assign nl_MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[14201:14184]));
  assign MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[14219:14202]));
  assign MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_455_nl = (readslicef_28_18_10((MultLoop_789_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_790_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_455_nl = nl_MultLoop_acc_455_nl[17:0];
  assign nl_MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[14237:14220]));
  assign MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[14255:14238]));
  assign MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_454_nl = (readslicef_28_18_10((MultLoop_791_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_792_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_454_nl = nl_MultLoop_acc_454_nl[17:0];
  assign nl_MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[14273:14256]));
  assign MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[14291:14274]));
  assign MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_453_nl = (readslicef_28_18_10((MultLoop_793_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_794_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_453_nl = nl_MultLoop_acc_453_nl[17:0];
  assign nl_MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[14309:14292]));
  assign MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[14327:14310]));
  assign MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_452_nl = (readslicef_28_18_10((MultLoop_795_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_796_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_452_nl = nl_MultLoop_acc_452_nl[17:0];
  assign nl_MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[14345:14328]));
  assign MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[14363:14346]));
  assign MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_451_nl = (readslicef_28_18_10((MultLoop_797_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_798_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_451_nl = nl_MultLoop_acc_451_nl[17:0];
  assign nl_MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[14525:14508]));
  assign MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[14543:14526]));
  assign MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_446_nl = (readslicef_28_18_10((MultLoop_807_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_808_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_446_nl = nl_MultLoop_acc_446_nl[17:0];
  assign nl_MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[14561:14544]));
  assign MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[14579:14562]));
  assign MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_445_nl = (readslicef_28_18_10((MultLoop_809_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_810_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_445_nl = nl_MultLoop_acc_445_nl[17:0];
  assign nl_MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[14597:14580]));
  assign MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[14615:14598]));
  assign MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_444_nl = (readslicef_28_18_10((MultLoop_811_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_812_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_444_nl = nl_MultLoop_acc_444_nl[17:0];
  assign nl_MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[14633:14616]));
  assign MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[14651:14634]));
  assign MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_443_nl = (readslicef_28_18_10((MultLoop_813_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_814_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_443_nl = nl_MultLoop_acc_443_nl[17:0];
  assign nl_MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[14381:14364]));
  assign MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[14399:14382]));
  assign MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_450_nl = (readslicef_28_18_10((MultLoop_799_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_800_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_450_nl = nl_MultLoop_acc_450_nl[17:0];
  assign nl_MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[14417:14400]));
  assign MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[14435:14418]));
  assign MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_449_nl = (readslicef_28_18_10((MultLoop_801_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_802_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_449_nl = nl_MultLoop_acc_449_nl[17:0];
  assign nl_MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[14453:14436]));
  assign MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[14471:14454]));
  assign MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_448_nl = (readslicef_28_18_10((MultLoop_803_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_804_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_448_nl = nl_MultLoop_acc_448_nl[17:0];
  assign nl_MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[14489:14472]));
  assign MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[14507:14490]));
  assign MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_447_nl = (readslicef_28_18_10((MultLoop_805_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_806_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_447_nl = nl_MultLoop_acc_447_nl[17:0];
  assign nl_MultLoop_acc_488_nl = (MultLoop_acc_458_nl) + (MultLoop_acc_457_nl) +
      (MultLoop_acc_456_nl) + (MultLoop_acc_455_nl) + (MultLoop_acc_454_nl) + (MultLoop_acc_453_nl)
      + (MultLoop_acc_452_nl) + (MultLoop_acc_451_nl) + (MultLoop_acc_446_nl) + (MultLoop_acc_445_nl)
      + (MultLoop_acc_444_nl) + (MultLoop_acc_443_nl) + (MultLoop_acc_450_nl) + (MultLoop_acc_449_nl)
      + (MultLoop_acc_448_nl) + (MultLoop_acc_447_nl);
  assign MultLoop_acc_488_nl = nl_MultLoop_acc_488_nl[17:0];
  assign nl_MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[13949:13932]));
  assign MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[13967:13950]));
  assign MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_462_nl = (readslicef_28_18_10((MultLoop_775_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_776_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_462_nl = nl_MultLoop_acc_462_nl[17:0];
  assign nl_MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[13985:13968]));
  assign MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[14003:13986]));
  assign MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_461_nl = (readslicef_28_18_10((MultLoop_777_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_778_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_461_nl = nl_MultLoop_acc_461_nl[17:0];
  assign nl_MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[14669:14652]));
  assign MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[14687:14670]));
  assign MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_442_nl = (readslicef_28_18_10((MultLoop_815_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_816_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_442_nl = nl_MultLoop_acc_442_nl[17:0];
  assign nl_MultLoop_acc_466_nl = (MultLoop_acc_442_nl) + (biases_rsci_idat[305:288]);
  assign MultLoop_acc_466_nl = nl_MultLoop_acc_466_nl[17:0];
  assign nl_MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[13841:13824]));
  assign MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[13859:13842]));
  assign MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_465_nl = (readslicef_28_18_10((MultLoop_769_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_770_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_465_nl = nl_MultLoop_acc_465_nl[17:0];
  assign nl_MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[13877:13860]));
  assign MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[13895:13878]));
  assign MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_464_nl = (readslicef_28_18_10((MultLoop_771_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_772_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_464_nl = nl_MultLoop_acc_464_nl[17:0];
  assign nl_MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[13913:13896]));
  assign MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[13931:13914]));
  assign MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_463_nl = (readslicef_28_18_10((MultLoop_773_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_774_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_463_nl = nl_MultLoop_acc_463_nl[17:0];
  assign nl_MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[14021:14004]));
  assign MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[14039:14022]));
  assign MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_460_nl = (readslicef_28_18_10((MultLoop_779_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_780_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_460_nl = nl_MultLoop_acc_460_nl[17:0];
  assign nl_MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[14057:14040]));
  assign MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[14075:14058]));
  assign MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_459_nl = (readslicef_28_18_10((MultLoop_781_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_782_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_459_nl = nl_MultLoop_acc_459_nl[17:0];
  assign nl_MultLoop_acc_487_nl = (MultLoop_acc_462_nl) + (MultLoop_acc_461_nl) +
      (MultLoop_acc_466_nl) + (MultLoop_acc_465_nl) + (MultLoop_acc_464_nl) + (MultLoop_acc_463_nl)
      + (MultLoop_acc_460_nl) + (MultLoop_acc_459_nl);
  assign MultLoop_acc_487_nl = nl_MultLoop_acc_487_nl[17:0];
  assign nl_res_rsci_d_305_288  = (MultLoop_acc_488_nl) + (MultLoop_acc_487_nl);
  assign nl_MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[6317:6300]));
  assign MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[6335:6318]));
  assign MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_881_nl = (readslicef_28_18_10((MultLoop_351_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_352_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_881_nl = nl_MultLoop_acc_881_nl[17:0];
  assign nl_MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[6353:6336]));
  assign MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[6371:6354]));
  assign MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_880_nl = (readslicef_28_18_10((MultLoop_353_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_354_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_880_nl = nl_MultLoop_acc_880_nl[17:0];
  assign nl_MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[6389:6372]));
  assign MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[6407:6390]));
  assign MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_879_nl = (readslicef_28_18_10((MultLoop_355_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_356_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_879_nl = nl_MultLoop_acc_879_nl[17:0];
  assign nl_MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[6425:6408]));
  assign MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[6443:6426]));
  assign MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_878_nl = (readslicef_28_18_10((MultLoop_357_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_358_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_878_nl = nl_MultLoop_acc_878_nl[17:0];
  assign nl_MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[6461:6444]));
  assign MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[6479:6462]));
  assign MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_877_nl = (readslicef_28_18_10((MultLoop_359_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_360_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_877_nl = nl_MultLoop_acc_877_nl[17:0];
  assign nl_MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[6497:6480]));
  assign MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[6515:6498]));
  assign MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_876_nl = (readslicef_28_18_10((MultLoop_361_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_362_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_876_nl = nl_MultLoop_acc_876_nl[17:0];
  assign nl_MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[6533:6516]));
  assign MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[6551:6534]));
  assign MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_875_nl = (readslicef_28_18_10((MultLoop_363_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_364_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_875_nl = nl_MultLoop_acc_875_nl[17:0];
  assign nl_MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[6569:6552]));
  assign MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[6587:6570]));
  assign MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_874_nl = (readslicef_28_18_10((MultLoop_365_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_366_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_874_nl = nl_MultLoop_acc_874_nl[17:0];
  assign nl_MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[6749:6732]));
  assign MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[6767:6750]));
  assign MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_869_nl = (readslicef_28_18_10((MultLoop_375_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_376_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_869_nl = nl_MultLoop_acc_869_nl[17:0];
  assign nl_MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[6785:6768]));
  assign MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[6803:6786]));
  assign MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_868_nl = (readslicef_28_18_10((MultLoop_377_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_378_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_868_nl = nl_MultLoop_acc_868_nl[17:0];
  assign nl_MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[6821:6804]));
  assign MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[6839:6822]));
  assign MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_867_nl = (readslicef_28_18_10((MultLoop_379_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_380_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_867_nl = nl_MultLoop_acc_867_nl[17:0];
  assign nl_MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[6857:6840]));
  assign MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[6875:6858]));
  assign MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_866_nl = (readslicef_28_18_10((MultLoop_381_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_382_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_866_nl = nl_MultLoop_acc_866_nl[17:0];
  assign nl_MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[6605:6588]));
  assign MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[6623:6606]));
  assign MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_873_nl = (readslicef_28_18_10((MultLoop_367_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_368_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_873_nl = nl_MultLoop_acc_873_nl[17:0];
  assign nl_MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[6641:6624]));
  assign MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[6659:6642]));
  assign MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_872_nl = (readslicef_28_18_10((MultLoop_369_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_370_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_872_nl = nl_MultLoop_acc_872_nl[17:0];
  assign nl_MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[6677:6660]));
  assign MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[6695:6678]));
  assign MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_871_nl = (readslicef_28_18_10((MultLoop_371_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_372_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_871_nl = nl_MultLoop_acc_871_nl[17:0];
  assign nl_MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[6713:6696]));
  assign MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[6731:6714]));
  assign MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_870_nl = (readslicef_28_18_10((MultLoop_373_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_374_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_870_nl = nl_MultLoop_acc_870_nl[17:0];
  assign nl_MultLoop_acc_911_nl = (MultLoop_acc_881_nl) + (MultLoop_acc_880_nl) +
      (MultLoop_acc_879_nl) + (MultLoop_acc_878_nl) + (MultLoop_acc_877_nl) + (MultLoop_acc_876_nl)
      + (MultLoop_acc_875_nl) + (MultLoop_acc_874_nl) + (MultLoop_acc_869_nl) + (MultLoop_acc_868_nl)
      + (MultLoop_acc_867_nl) + (MultLoop_acc_866_nl) + (MultLoop_acc_873_nl) + (MultLoop_acc_872_nl)
      + (MultLoop_acc_871_nl) + (MultLoop_acc_870_nl);
  assign MultLoop_acc_911_nl = nl_MultLoop_acc_911_nl[17:0];
  assign nl_MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[6173:6156]));
  assign MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[6191:6174]));
  assign MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_885_nl = (readslicef_28_18_10((MultLoop_343_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_344_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_885_nl = nl_MultLoop_acc_885_nl[17:0];
  assign nl_MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[6209:6192]));
  assign MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[6227:6210]));
  assign MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_884_nl = (readslicef_28_18_10((MultLoop_345_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_346_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_884_nl = nl_MultLoop_acc_884_nl[17:0];
  assign nl_MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[6893:6876]));
  assign MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[6911:6894]));
  assign MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_865_nl = (readslicef_28_18_10((MultLoop_383_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_384_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_865_nl = nl_MultLoop_acc_865_nl[17:0];
  assign nl_MultLoop_acc_889_nl = (MultLoop_acc_865_nl) + (biases_rsci_idat[143:126]);
  assign MultLoop_acc_889_nl = nl_MultLoop_acc_889_nl[17:0];
  assign nl_MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[6065:6048]));
  assign MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[6083:6066]));
  assign MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_888_nl = (readslicef_28_18_10((MultLoop_337_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_338_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_888_nl = nl_MultLoop_acc_888_nl[17:0];
  assign nl_MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[6101:6084]));
  assign MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[6119:6102]));
  assign MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_887_nl = (readslicef_28_18_10((MultLoop_339_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_340_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_887_nl = nl_MultLoop_acc_887_nl[17:0];
  assign nl_MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[6137:6120]));
  assign MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[6155:6138]));
  assign MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_886_nl = (readslicef_28_18_10((MultLoop_341_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_342_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_886_nl = nl_MultLoop_acc_886_nl[17:0];
  assign nl_MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[6245:6228]));
  assign MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[6263:6246]));
  assign MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_883_nl = (readslicef_28_18_10((MultLoop_347_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_348_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_883_nl = nl_MultLoop_acc_883_nl[17:0];
  assign nl_MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[6281:6264]));
  assign MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[6299:6282]));
  assign MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_882_nl = (readslicef_28_18_10((MultLoop_349_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_350_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_882_nl = nl_MultLoop_acc_882_nl[17:0];
  assign nl_MultLoop_acc_910_nl = (MultLoop_acc_885_nl) + (MultLoop_acc_884_nl) +
      (MultLoop_acc_889_nl) + (MultLoop_acc_888_nl) + (MultLoop_acc_887_nl) + (MultLoop_acc_886_nl)
      + (MultLoop_acc_883_nl) + (MultLoop_acc_882_nl);
  assign MultLoop_acc_910_nl = nl_MultLoop_acc_910_nl[17:0];
  assign nl_res_rsci_d_143_126  = (MultLoop_acc_911_nl) + (MultLoop_acc_910_nl);
  assign nl_MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[13229:13212]));
  assign MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[13247:13230]));
  assign MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_505_nl = (readslicef_28_18_10((MultLoop_735_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_736_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_505_nl = nl_MultLoop_acc_505_nl[17:0];
  assign nl_MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[13265:13248]));
  assign MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[13283:13266]));
  assign MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_504_nl = (readslicef_28_18_10((MultLoop_737_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_738_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_504_nl = nl_MultLoop_acc_504_nl[17:0];
  assign nl_MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[13301:13284]));
  assign MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[13319:13302]));
  assign MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_503_nl = (readslicef_28_18_10((MultLoop_739_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_740_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_503_nl = nl_MultLoop_acc_503_nl[17:0];
  assign nl_MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[13337:13320]));
  assign MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[13355:13338]));
  assign MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_502_nl = (readslicef_28_18_10((MultLoop_741_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_742_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_502_nl = nl_MultLoop_acc_502_nl[17:0];
  assign nl_MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[13373:13356]));
  assign MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[13391:13374]));
  assign MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_501_nl = (readslicef_28_18_10((MultLoop_743_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_744_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_501_nl = nl_MultLoop_acc_501_nl[17:0];
  assign nl_MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[13409:13392]));
  assign MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[13427:13410]));
  assign MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_500_nl = (readslicef_28_18_10((MultLoop_745_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_746_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_500_nl = nl_MultLoop_acc_500_nl[17:0];
  assign nl_MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[13445:13428]));
  assign MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[13463:13446]));
  assign MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_499_nl = (readslicef_28_18_10((MultLoop_747_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_748_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_499_nl = nl_MultLoop_acc_499_nl[17:0];
  assign nl_MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[13481:13464]));
  assign MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[13499:13482]));
  assign MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_498_nl = (readslicef_28_18_10((MultLoop_749_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_750_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_498_nl = nl_MultLoop_acc_498_nl[17:0];
  assign nl_MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[13661:13644]));
  assign MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[13679:13662]));
  assign MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_493_nl = (readslicef_28_18_10((MultLoop_759_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_760_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_493_nl = nl_MultLoop_acc_493_nl[17:0];
  assign nl_MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[13697:13680]));
  assign MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[13715:13698]));
  assign MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_492_nl = (readslicef_28_18_10((MultLoop_761_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_762_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_492_nl = nl_MultLoop_acc_492_nl[17:0];
  assign nl_MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[13733:13716]));
  assign MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[13751:13734]));
  assign MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_491_nl = (readslicef_28_18_10((MultLoop_763_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_764_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_491_nl = nl_MultLoop_acc_491_nl[17:0];
  assign nl_MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[13769:13752]));
  assign MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[13787:13770]));
  assign MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_490_nl = (readslicef_28_18_10((MultLoop_765_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_766_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_490_nl = nl_MultLoop_acc_490_nl[17:0];
  assign nl_MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[13517:13500]));
  assign MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[13535:13518]));
  assign MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_497_nl = (readslicef_28_18_10((MultLoop_751_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_752_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_497_nl = nl_MultLoop_acc_497_nl[17:0];
  assign nl_MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[13553:13536]));
  assign MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[13571:13554]));
  assign MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_496_nl = (readslicef_28_18_10((MultLoop_753_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_754_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_496_nl = nl_MultLoop_acc_496_nl[17:0];
  assign nl_MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[13589:13572]));
  assign MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[13607:13590]));
  assign MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_495_nl = (readslicef_28_18_10((MultLoop_755_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_756_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_495_nl = nl_MultLoop_acc_495_nl[17:0];
  assign nl_MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[13625:13608]));
  assign MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[13643:13626]));
  assign MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_494_nl = (readslicef_28_18_10((MultLoop_757_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_758_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_494_nl = nl_MultLoop_acc_494_nl[17:0];
  assign nl_MultLoop_acc_535_nl = (MultLoop_acc_505_nl) + (MultLoop_acc_504_nl) +
      (MultLoop_acc_503_nl) + (MultLoop_acc_502_nl) + (MultLoop_acc_501_nl) + (MultLoop_acc_500_nl)
      + (MultLoop_acc_499_nl) + (MultLoop_acc_498_nl) + (MultLoop_acc_493_nl) + (MultLoop_acc_492_nl)
      + (MultLoop_acc_491_nl) + (MultLoop_acc_490_nl) + (MultLoop_acc_497_nl) + (MultLoop_acc_496_nl)
      + (MultLoop_acc_495_nl) + (MultLoop_acc_494_nl);
  assign MultLoop_acc_535_nl = nl_MultLoop_acc_535_nl[17:0];
  assign nl_MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[13085:13068]));
  assign MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[13103:13086]));
  assign MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_509_nl = (readslicef_28_18_10((MultLoop_727_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_509_nl = nl_MultLoop_acc_509_nl[17:0];
  assign nl_MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[13121:13104]));
  assign MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[13139:13122]));
  assign MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_508_nl = (readslicef_28_18_10((MultLoop_729_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_730_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_508_nl = nl_MultLoop_acc_508_nl[17:0];
  assign nl_MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[13805:13788]));
  assign MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[13823:13806]));
  assign MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_489_nl = (readslicef_28_18_10((MultLoop_767_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_768_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_489_nl = nl_MultLoop_acc_489_nl[17:0];
  assign nl_MultLoop_acc_513_nl = (MultLoop_acc_489_nl) + (biases_rsci_idat[287:270]);
  assign MultLoop_acc_513_nl = nl_MultLoop_acc_513_nl[17:0];
  assign nl_MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[12977:12960]));
  assign MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[12995:12978]));
  assign MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_512_nl = (readslicef_28_18_10((MultLoop_721_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_722_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_512_nl = nl_MultLoop_acc_512_nl[17:0];
  assign nl_MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[13013:12996]));
  assign MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[13031:13014]));
  assign MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_511_nl = (readslicef_28_18_10((MultLoop_723_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_724_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_511_nl = nl_MultLoop_acc_511_nl[17:0];
  assign nl_MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[13049:13032]));
  assign MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[13067:13050]));
  assign MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_510_nl = (readslicef_28_18_10((MultLoop_725_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_726_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_510_nl = nl_MultLoop_acc_510_nl[17:0];
  assign nl_MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[13157:13140]));
  assign MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[13175:13158]));
  assign MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_507_nl = (readslicef_28_18_10((MultLoop_731_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_732_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_507_nl = nl_MultLoop_acc_507_nl[17:0];
  assign nl_MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[13193:13176]));
  assign MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[13211:13194]));
  assign MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_506_nl = (readslicef_28_18_10((MultLoop_733_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_734_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_506_nl = nl_MultLoop_acc_506_nl[17:0];
  assign nl_MultLoop_acc_534_nl = (MultLoop_acc_509_nl) + (MultLoop_acc_508_nl) +
      (MultLoop_acc_513_nl) + (MultLoop_acc_512_nl) + (MultLoop_acc_511_nl) + (MultLoop_acc_510_nl)
      + (MultLoop_acc_507_nl) + (MultLoop_acc_506_nl);
  assign MultLoop_acc_534_nl = nl_MultLoop_acc_534_nl[17:0];
  assign nl_res_rsci_d_287_270  = (MultLoop_acc_535_nl) + (MultLoop_acc_534_nl);
  assign nl_MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[7181:7164]));
  assign MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[7199:7182]));
  assign MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_834_nl = (readslicef_28_18_10((MultLoop_399_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_400_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_834_nl = nl_MultLoop_acc_834_nl[17:0];
  assign nl_MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[7217:7200]));
  assign MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[7235:7218]));
  assign MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_833_nl = (readslicef_28_18_10((MultLoop_401_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_402_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_833_nl = nl_MultLoop_acc_833_nl[17:0];
  assign nl_MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[7253:7236]));
  assign MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[7271:7254]));
  assign MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_832_nl = (readslicef_28_18_10((MultLoop_403_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_404_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_832_nl = nl_MultLoop_acc_832_nl[17:0];
  assign nl_MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[7289:7272]));
  assign MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[7307:7290]));
  assign MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_831_nl = (readslicef_28_18_10((MultLoop_405_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_406_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_831_nl = nl_MultLoop_acc_831_nl[17:0];
  assign nl_MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[7325:7308]));
  assign MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[7343:7326]));
  assign MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_830_nl = (readslicef_28_18_10((MultLoop_407_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_408_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_830_nl = nl_MultLoop_acc_830_nl[17:0];
  assign nl_MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[7361:7344]));
  assign MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[7379:7362]));
  assign MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_829_nl = (readslicef_28_18_10((MultLoop_409_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_410_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_829_nl = nl_MultLoop_acc_829_nl[17:0];
  assign nl_MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[7397:7380]));
  assign MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[7415:7398]));
  assign MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_828_nl = (readslicef_28_18_10((MultLoop_411_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_412_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_828_nl = nl_MultLoop_acc_828_nl[17:0];
  assign nl_MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[7433:7416]));
  assign MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[7451:7434]));
  assign MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_827_nl = (readslicef_28_18_10((MultLoop_413_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_414_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_827_nl = nl_MultLoop_acc_827_nl[17:0];
  assign nl_MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[7613:7596]));
  assign MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[7631:7614]));
  assign MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_822_nl = (readslicef_28_18_10((MultLoop_423_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_424_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_822_nl = nl_MultLoop_acc_822_nl[17:0];
  assign nl_MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[7649:7632]));
  assign MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[7667:7650]));
  assign MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_821_nl = (readslicef_28_18_10((MultLoop_425_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_426_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_821_nl = nl_MultLoop_acc_821_nl[17:0];
  assign nl_MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[7685:7668]));
  assign MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[7703:7686]));
  assign MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_820_nl = (readslicef_28_18_10((MultLoop_427_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_428_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_820_nl = nl_MultLoop_acc_820_nl[17:0];
  assign nl_MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[7721:7704]));
  assign MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[7739:7722]));
  assign MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_819_nl = (readslicef_28_18_10((MultLoop_429_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_430_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_819_nl = nl_MultLoop_acc_819_nl[17:0];
  assign nl_MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[7469:7452]));
  assign MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[7487:7470]));
  assign MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_826_nl = (readslicef_28_18_10((MultLoop_415_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_416_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_826_nl = nl_MultLoop_acc_826_nl[17:0];
  assign nl_MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[7505:7488]));
  assign MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[7523:7506]));
  assign MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_825_nl = (readslicef_28_18_10((MultLoop_417_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_418_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_825_nl = nl_MultLoop_acc_825_nl[17:0];
  assign nl_MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[7541:7524]));
  assign MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[7559:7542]));
  assign MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_824_nl = (readslicef_28_18_10((MultLoop_419_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_420_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_824_nl = nl_MultLoop_acc_824_nl[17:0];
  assign nl_MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[7577:7560]));
  assign MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[7595:7578]));
  assign MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_823_nl = (readslicef_28_18_10((MultLoop_421_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_422_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_823_nl = nl_MultLoop_acc_823_nl[17:0];
  assign nl_MultLoop_acc_864_nl = (MultLoop_acc_834_nl) + (MultLoop_acc_833_nl) +
      (MultLoop_acc_832_nl) + (MultLoop_acc_831_nl) + (MultLoop_acc_830_nl) + (MultLoop_acc_829_nl)
      + (MultLoop_acc_828_nl) + (MultLoop_acc_827_nl) + (MultLoop_acc_822_nl) + (MultLoop_acc_821_nl)
      + (MultLoop_acc_820_nl) + (MultLoop_acc_819_nl) + (MultLoop_acc_826_nl) + (MultLoop_acc_825_nl)
      + (MultLoop_acc_824_nl) + (MultLoop_acc_823_nl);
  assign MultLoop_acc_864_nl = nl_MultLoop_acc_864_nl[17:0];
  assign nl_MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[7037:7020]));
  assign MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[7055:7038]));
  assign MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_838_nl = (readslicef_28_18_10((MultLoop_391_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_392_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_838_nl = nl_MultLoop_acc_838_nl[17:0];
  assign nl_MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[7073:7056]));
  assign MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[7091:7074]));
  assign MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_837_nl = (readslicef_28_18_10((MultLoop_393_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_394_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_837_nl = nl_MultLoop_acc_837_nl[17:0];
  assign nl_MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[7757:7740]));
  assign MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[7775:7758]));
  assign MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_818_nl = (readslicef_28_18_10((MultLoop_431_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_432_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_818_nl = nl_MultLoop_acc_818_nl[17:0];
  assign nl_MultLoop_acc_842_nl = (MultLoop_acc_818_nl) + (biases_rsci_idat[161:144]);
  assign MultLoop_acc_842_nl = nl_MultLoop_acc_842_nl[17:0];
  assign nl_MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[6929:6912]));
  assign MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[6947:6930]));
  assign MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_841_nl = (readslicef_28_18_10((MultLoop_385_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_386_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_841_nl = nl_MultLoop_acc_841_nl[17:0];
  assign nl_MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[6965:6948]));
  assign MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[6983:6966]));
  assign MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_840_nl = (readslicef_28_18_10((MultLoop_387_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_388_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_840_nl = nl_MultLoop_acc_840_nl[17:0];
  assign nl_MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[7001:6984]));
  assign MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[7019:7002]));
  assign MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_839_nl = (readslicef_28_18_10((MultLoop_389_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_390_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_839_nl = nl_MultLoop_acc_839_nl[17:0];
  assign nl_MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[7109:7092]));
  assign MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[7127:7110]));
  assign MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_836_nl = (readslicef_28_18_10((MultLoop_395_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_396_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_836_nl = nl_MultLoop_acc_836_nl[17:0];
  assign nl_MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[7145:7128]));
  assign MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[7163:7146]));
  assign MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_835_nl = (readslicef_28_18_10((MultLoop_397_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_398_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_835_nl = nl_MultLoop_acc_835_nl[17:0];
  assign nl_MultLoop_acc_863_nl = (MultLoop_acc_838_nl) + (MultLoop_acc_837_nl) +
      (MultLoop_acc_842_nl) + (MultLoop_acc_841_nl) + (MultLoop_acc_840_nl) + (MultLoop_acc_839_nl)
      + (MultLoop_acc_836_nl) + (MultLoop_acc_835_nl);
  assign MultLoop_acc_863_nl = nl_MultLoop_acc_863_nl[17:0];
  assign nl_res_rsci_d_161_144  = (MultLoop_acc_864_nl) + (MultLoop_acc_863_nl);
  assign nl_MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[12365:12348]));
  assign MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[12383:12366]));
  assign MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_552_nl = (readslicef_28_18_10((MultLoop_687_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_688_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_552_nl = nl_MultLoop_acc_552_nl[17:0];
  assign nl_MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[12401:12384]));
  assign MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[12419:12402]));
  assign MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_551_nl = (readslicef_28_18_10((MultLoop_689_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_690_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_551_nl = nl_MultLoop_acc_551_nl[17:0];
  assign nl_MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[12437:12420]));
  assign MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[12455:12438]));
  assign MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_550_nl = (readslicef_28_18_10((MultLoop_691_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_692_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_550_nl = nl_MultLoop_acc_550_nl[17:0];
  assign nl_MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[12473:12456]));
  assign MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[12491:12474]));
  assign MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_549_nl = (readslicef_28_18_10((MultLoop_693_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_694_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_549_nl = nl_MultLoop_acc_549_nl[17:0];
  assign nl_MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[12509:12492]));
  assign MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[12527:12510]));
  assign MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_548_nl = (readslicef_28_18_10((MultLoop_695_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_696_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_548_nl = nl_MultLoop_acc_548_nl[17:0];
  assign nl_MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[12545:12528]));
  assign MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[12563:12546]));
  assign MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_547_nl = (readslicef_28_18_10((MultLoop_697_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_698_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_547_nl = nl_MultLoop_acc_547_nl[17:0];
  assign nl_MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[12581:12564]));
  assign MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[12599:12582]));
  assign MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_546_nl = (readslicef_28_18_10((MultLoop_699_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_700_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_546_nl = nl_MultLoop_acc_546_nl[17:0];
  assign nl_MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[12617:12600]));
  assign MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[12635:12618]));
  assign MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_545_nl = (readslicef_28_18_10((MultLoop_701_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_702_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_545_nl = nl_MultLoop_acc_545_nl[17:0];
  assign nl_MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[12797:12780]));
  assign MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[12815:12798]));
  assign MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_540_nl = (readslicef_28_18_10((MultLoop_711_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_712_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_540_nl = nl_MultLoop_acc_540_nl[17:0];
  assign nl_MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[12833:12816]));
  assign MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[12851:12834]));
  assign MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_539_nl = (readslicef_28_18_10((MultLoop_713_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_714_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_539_nl = nl_MultLoop_acc_539_nl[17:0];
  assign nl_MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[12869:12852]));
  assign MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[12887:12870]));
  assign MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_538_nl = (readslicef_28_18_10((MultLoop_715_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_716_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_538_nl = nl_MultLoop_acc_538_nl[17:0];
  assign nl_MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[12905:12888]));
  assign MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[12923:12906]));
  assign MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_537_nl = (readslicef_28_18_10((MultLoop_717_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_718_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_537_nl = nl_MultLoop_acc_537_nl[17:0];
  assign nl_MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[12653:12636]));
  assign MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[12671:12654]));
  assign MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_544_nl = (readslicef_28_18_10((MultLoop_703_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_704_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_544_nl = nl_MultLoop_acc_544_nl[17:0];
  assign nl_MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[12689:12672]));
  assign MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[12707:12690]));
  assign MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_543_nl = (readslicef_28_18_10((MultLoop_705_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_706_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_543_nl = nl_MultLoop_acc_543_nl[17:0];
  assign nl_MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[12725:12708]));
  assign MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[12743:12726]));
  assign MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_542_nl = (readslicef_28_18_10((MultLoop_707_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_708_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_542_nl = nl_MultLoop_acc_542_nl[17:0];
  assign nl_MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[12761:12744]));
  assign MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[12779:12762]));
  assign MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_541_nl = (readslicef_28_18_10((MultLoop_709_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_710_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_541_nl = nl_MultLoop_acc_541_nl[17:0];
  assign nl_MultLoop_acc_582_nl = (MultLoop_acc_552_nl) + (MultLoop_acc_551_nl) +
      (MultLoop_acc_550_nl) + (MultLoop_acc_549_nl) + (MultLoop_acc_548_nl) + (MultLoop_acc_547_nl)
      + (MultLoop_acc_546_nl) + (MultLoop_acc_545_nl) + (MultLoop_acc_540_nl) + (MultLoop_acc_539_nl)
      + (MultLoop_acc_538_nl) + (MultLoop_acc_537_nl) + (MultLoop_acc_544_nl) + (MultLoop_acc_543_nl)
      + (MultLoop_acc_542_nl) + (MultLoop_acc_541_nl);
  assign MultLoop_acc_582_nl = nl_MultLoop_acc_582_nl[17:0];
  assign nl_MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[12221:12204]));
  assign MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[12239:12222]));
  assign MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_556_nl = (readslicef_28_18_10((MultLoop_679_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_680_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_556_nl = nl_MultLoop_acc_556_nl[17:0];
  assign nl_MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[12257:12240]));
  assign MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[12275:12258]));
  assign MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_555_nl = (readslicef_28_18_10((MultLoop_681_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_682_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_555_nl = nl_MultLoop_acc_555_nl[17:0];
  assign nl_MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[12941:12924]));
  assign MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[12959:12942]));
  assign MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_536_nl = (readslicef_28_18_10((MultLoop_719_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_720_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_536_nl = nl_MultLoop_acc_536_nl[17:0];
  assign nl_MultLoop_acc_560_nl = (MultLoop_acc_536_nl) + (biases_rsci_idat[269:252]);
  assign MultLoop_acc_560_nl = nl_MultLoop_acc_560_nl[17:0];
  assign nl_MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[12113:12096]));
  assign MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[12131:12114]));
  assign MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_559_nl = (readslicef_28_18_10((MultLoop_673_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_674_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_559_nl = nl_MultLoop_acc_559_nl[17:0];
  assign nl_MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[12149:12132]));
  assign MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[12167:12150]));
  assign MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_558_nl = (readslicef_28_18_10((MultLoop_675_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_676_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_558_nl = nl_MultLoop_acc_558_nl[17:0];
  assign nl_MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[12185:12168]));
  assign MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[12203:12186]));
  assign MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_557_nl = (readslicef_28_18_10((MultLoop_677_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_678_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_557_nl = nl_MultLoop_acc_557_nl[17:0];
  assign nl_MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[12293:12276]));
  assign MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[12311:12294]));
  assign MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_554_nl = (readslicef_28_18_10((MultLoop_683_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_684_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_554_nl = nl_MultLoop_acc_554_nl[17:0];
  assign nl_MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[12329:12312]));
  assign MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[12347:12330]));
  assign MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_553_nl = (readslicef_28_18_10((MultLoop_685_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_686_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_553_nl = nl_MultLoop_acc_553_nl[17:0];
  assign nl_MultLoop_acc_581_nl = (MultLoop_acc_556_nl) + (MultLoop_acc_555_nl) +
      (MultLoop_acc_560_nl) + (MultLoop_acc_559_nl) + (MultLoop_acc_558_nl) + (MultLoop_acc_557_nl)
      + (MultLoop_acc_554_nl) + (MultLoop_acc_553_nl);
  assign MultLoop_acc_581_nl = nl_MultLoop_acc_581_nl[17:0];
  assign nl_res_rsci_d_269_252  = (MultLoop_acc_582_nl) + (MultLoop_acc_581_nl);
  assign nl_MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[8045:8028]));
  assign MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[8063:8046]));
  assign MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_787_nl = (readslicef_28_18_10((MultLoop_447_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_448_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_787_nl = nl_MultLoop_acc_787_nl[17:0];
  assign nl_MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[8081:8064]));
  assign MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[8099:8082]));
  assign MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_786_nl = (readslicef_28_18_10((MultLoop_449_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_450_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_786_nl = nl_MultLoop_acc_786_nl[17:0];
  assign nl_MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[8117:8100]));
  assign MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[8135:8118]));
  assign MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_785_nl = (readslicef_28_18_10((MultLoop_451_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_452_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_785_nl = nl_MultLoop_acc_785_nl[17:0];
  assign nl_MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[8153:8136]));
  assign MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[8171:8154]));
  assign MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_784_nl = (readslicef_28_18_10((MultLoop_453_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_454_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_784_nl = nl_MultLoop_acc_784_nl[17:0];
  assign nl_MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[8189:8172]));
  assign MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[8207:8190]));
  assign MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_783_nl = (readslicef_28_18_10((MultLoop_455_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_456_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_783_nl = nl_MultLoop_acc_783_nl[17:0];
  assign nl_MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[8225:8208]));
  assign MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[8243:8226]));
  assign MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_782_nl = (readslicef_28_18_10((MultLoop_457_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_458_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_782_nl = nl_MultLoop_acc_782_nl[17:0];
  assign nl_MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[8261:8244]));
  assign MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[8279:8262]));
  assign MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_781_nl = (readslicef_28_18_10((MultLoop_459_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_460_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_781_nl = nl_MultLoop_acc_781_nl[17:0];
  assign nl_MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[8297:8280]));
  assign MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[8315:8298]));
  assign MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_780_nl = (readslicef_28_18_10((MultLoop_461_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_462_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_780_nl = nl_MultLoop_acc_780_nl[17:0];
  assign nl_MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[8477:8460]));
  assign MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[8495:8478]));
  assign MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_775_nl = (readslicef_28_18_10((MultLoop_471_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_472_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_775_nl = nl_MultLoop_acc_775_nl[17:0];
  assign nl_MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[8513:8496]));
  assign MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[8531:8514]));
  assign MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_774_nl = (readslicef_28_18_10((MultLoop_473_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_474_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_774_nl = nl_MultLoop_acc_774_nl[17:0];
  assign nl_MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[8549:8532]));
  assign MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[8567:8550]));
  assign MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_773_nl = (readslicef_28_18_10((MultLoop_475_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_476_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_773_nl = nl_MultLoop_acc_773_nl[17:0];
  assign nl_MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[8585:8568]));
  assign MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[8603:8586]));
  assign MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_772_nl = (readslicef_28_18_10((MultLoop_477_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_478_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_772_nl = nl_MultLoop_acc_772_nl[17:0];
  assign nl_MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[8333:8316]));
  assign MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[8351:8334]));
  assign MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_779_nl = (readslicef_28_18_10((MultLoop_463_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_464_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_779_nl = nl_MultLoop_acc_779_nl[17:0];
  assign nl_MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[8369:8352]));
  assign MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[8387:8370]));
  assign MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_778_nl = (readslicef_28_18_10((MultLoop_465_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_466_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_778_nl = nl_MultLoop_acc_778_nl[17:0];
  assign nl_MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[8405:8388]));
  assign MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[8423:8406]));
  assign MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_777_nl = (readslicef_28_18_10((MultLoop_467_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_468_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_777_nl = nl_MultLoop_acc_777_nl[17:0];
  assign nl_MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[8441:8424]));
  assign MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[8459:8442]));
  assign MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_776_nl = (readslicef_28_18_10((MultLoop_469_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_470_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_776_nl = nl_MultLoop_acc_776_nl[17:0];
  assign nl_MultLoop_acc_817_nl = (MultLoop_acc_787_nl) + (MultLoop_acc_786_nl) +
      (MultLoop_acc_785_nl) + (MultLoop_acc_784_nl) + (MultLoop_acc_783_nl) + (MultLoop_acc_782_nl)
      + (MultLoop_acc_781_nl) + (MultLoop_acc_780_nl) + (MultLoop_acc_775_nl) + (MultLoop_acc_774_nl)
      + (MultLoop_acc_773_nl) + (MultLoop_acc_772_nl) + (MultLoop_acc_779_nl) + (MultLoop_acc_778_nl)
      + (MultLoop_acc_777_nl) + (MultLoop_acc_776_nl);
  assign MultLoop_acc_817_nl = nl_MultLoop_acc_817_nl[17:0];
  assign nl_MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[7901:7884]));
  assign MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[7919:7902]));
  assign MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_791_nl = (readslicef_28_18_10((MultLoop_439_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_440_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_791_nl = nl_MultLoop_acc_791_nl[17:0];
  assign nl_MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[7937:7920]));
  assign MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[7955:7938]));
  assign MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_790_nl = (readslicef_28_18_10((MultLoop_441_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_442_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_790_nl = nl_MultLoop_acc_790_nl[17:0];
  assign nl_MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[8621:8604]));
  assign MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[8639:8622]));
  assign MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_771_nl = (readslicef_28_18_10((MultLoop_479_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_480_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_771_nl = nl_MultLoop_acc_771_nl[17:0];
  assign nl_MultLoop_acc_795_nl = (MultLoop_acc_771_nl) + (biases_rsci_idat[179:162]);
  assign MultLoop_acc_795_nl = nl_MultLoop_acc_795_nl[17:0];
  assign nl_MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[7793:7776]));
  assign MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[7811:7794]));
  assign MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_794_nl = (readslicef_28_18_10((MultLoop_433_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_434_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_794_nl = nl_MultLoop_acc_794_nl[17:0];
  assign nl_MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[7829:7812]));
  assign MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[7847:7830]));
  assign MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_793_nl = (readslicef_28_18_10((MultLoop_435_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_436_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_793_nl = nl_MultLoop_acc_793_nl[17:0];
  assign nl_MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[7865:7848]));
  assign MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[7883:7866]));
  assign MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_792_nl = (readslicef_28_18_10((MultLoop_437_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_438_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_792_nl = nl_MultLoop_acc_792_nl[17:0];
  assign nl_MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[7973:7956]));
  assign MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[7991:7974]));
  assign MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_789_nl = (readslicef_28_18_10((MultLoop_443_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_444_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_789_nl = nl_MultLoop_acc_789_nl[17:0];
  assign nl_MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[8009:7992]));
  assign MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[8027:8010]));
  assign MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_788_nl = (readslicef_28_18_10((MultLoop_445_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_446_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_788_nl = nl_MultLoop_acc_788_nl[17:0];
  assign nl_MultLoop_acc_816_nl = (MultLoop_acc_791_nl) + (MultLoop_acc_790_nl) +
      (MultLoop_acc_795_nl) + (MultLoop_acc_794_nl) + (MultLoop_acc_793_nl) + (MultLoop_acc_792_nl)
      + (MultLoop_acc_789_nl) + (MultLoop_acc_788_nl);
  assign MultLoop_acc_816_nl = nl_MultLoop_acc_816_nl[17:0];
  assign nl_res_rsci_d_179_162  = (MultLoop_acc_817_nl) + (MultLoop_acc_816_nl);
  assign nl_MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[11501:11484]));
  assign MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[11519:11502]));
  assign MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_599_nl = (readslicef_28_18_10((MultLoop_639_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_640_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_599_nl = nl_MultLoop_acc_599_nl[17:0];
  assign nl_MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[11537:11520]));
  assign MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[11555:11538]));
  assign MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_598_nl = (readslicef_28_18_10((MultLoop_641_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_642_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_598_nl = nl_MultLoop_acc_598_nl[17:0];
  assign nl_MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[11573:11556]));
  assign MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[11591:11574]));
  assign MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_597_nl = (readslicef_28_18_10((MultLoop_643_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_644_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_597_nl = nl_MultLoop_acc_597_nl[17:0];
  assign nl_MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[11609:11592]));
  assign MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[11627:11610]));
  assign MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_596_nl = (readslicef_28_18_10((MultLoop_645_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_646_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_596_nl = nl_MultLoop_acc_596_nl[17:0];
  assign nl_MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[11645:11628]));
  assign MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[11663:11646]));
  assign MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_595_nl = (readslicef_28_18_10((MultLoop_647_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_648_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_595_nl = nl_MultLoop_acc_595_nl[17:0];
  assign nl_MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[11681:11664]));
  assign MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[11699:11682]));
  assign MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_594_nl = (readslicef_28_18_10((MultLoop_649_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_650_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_594_nl = nl_MultLoop_acc_594_nl[17:0];
  assign nl_MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[11717:11700]));
  assign MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[11735:11718]));
  assign MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_593_nl = (readslicef_28_18_10((MultLoop_651_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_652_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_593_nl = nl_MultLoop_acc_593_nl[17:0];
  assign nl_MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[11753:11736]));
  assign MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[11771:11754]));
  assign MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_592_nl = (readslicef_28_18_10((MultLoop_653_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_654_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_592_nl = nl_MultLoop_acc_592_nl[17:0];
  assign nl_MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[11933:11916]));
  assign MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[11951:11934]));
  assign MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_587_nl = (readslicef_28_18_10((MultLoop_663_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_664_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_587_nl = nl_MultLoop_acc_587_nl[17:0];
  assign nl_MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[11969:11952]));
  assign MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[11987:11970]));
  assign MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_586_nl = (readslicef_28_18_10((MultLoop_665_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_666_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_586_nl = nl_MultLoop_acc_586_nl[17:0];
  assign nl_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[12005:11988]));
  assign MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[12023:12006]));
  assign MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_585_nl = (readslicef_28_18_10((MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_668_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_585_nl = nl_MultLoop_acc_585_nl[17:0];
  assign nl_MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[12041:12024]));
  assign MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[12059:12042]));
  assign MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_584_nl = (readslicef_28_18_10((MultLoop_669_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_670_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_584_nl = nl_MultLoop_acc_584_nl[17:0];
  assign nl_MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[11789:11772]));
  assign MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[11807:11790]));
  assign MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_591_nl = (readslicef_28_18_10((MultLoop_655_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_656_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_591_nl = nl_MultLoop_acc_591_nl[17:0];
  assign nl_MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[11825:11808]));
  assign MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[11843:11826]));
  assign MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_590_nl = (readslicef_28_18_10((MultLoop_657_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_658_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_590_nl = nl_MultLoop_acc_590_nl[17:0];
  assign nl_MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[11861:11844]));
  assign MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[11879:11862]));
  assign MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_589_nl = (readslicef_28_18_10((MultLoop_659_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_660_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_589_nl = nl_MultLoop_acc_589_nl[17:0];
  assign nl_MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[11897:11880]));
  assign MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[11915:11898]));
  assign MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_588_nl = (readslicef_28_18_10((MultLoop_661_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_662_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_588_nl = nl_MultLoop_acc_588_nl[17:0];
  assign nl_MultLoop_acc_629_nl = (MultLoop_acc_599_nl) + (MultLoop_acc_598_nl) +
      (MultLoop_acc_597_nl) + (MultLoop_acc_596_nl) + (MultLoop_acc_595_nl) + (MultLoop_acc_594_nl)
      + (MultLoop_acc_593_nl) + (MultLoop_acc_592_nl) + (MultLoop_acc_587_nl) + (MultLoop_acc_586_nl)
      + (MultLoop_acc_585_nl) + (MultLoop_acc_584_nl) + (MultLoop_acc_591_nl) + (MultLoop_acc_590_nl)
      + (MultLoop_acc_589_nl) + (MultLoop_acc_588_nl);
  assign MultLoop_acc_629_nl = nl_MultLoop_acc_629_nl[17:0];
  assign nl_MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[11357:11340]));
  assign MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[11375:11358]));
  assign MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_603_nl = (readslicef_28_18_10((MultLoop_631_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_632_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_603_nl = nl_MultLoop_acc_603_nl[17:0];
  assign nl_MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[11393:11376]));
  assign MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[11411:11394]));
  assign MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_602_nl = (readslicef_28_18_10((MultLoop_633_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_634_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_602_nl = nl_MultLoop_acc_602_nl[17:0];
  assign nl_MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[12077:12060]));
  assign MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[12095:12078]));
  assign MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_583_nl = (readslicef_28_18_10((MultLoop_671_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_672_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_583_nl = nl_MultLoop_acc_583_nl[17:0];
  assign nl_MultLoop_acc_607_nl = (MultLoop_acc_583_nl) + (biases_rsci_idat[251:234]);
  assign MultLoop_acc_607_nl = nl_MultLoop_acc_607_nl[17:0];
  assign nl_MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[11249:11232]));
  assign MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[11267:11250]));
  assign MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_606_nl = (readslicef_28_18_10((MultLoop_625_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_626_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_606_nl = nl_MultLoop_acc_606_nl[17:0];
  assign nl_MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[11285:11268]));
  assign MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[11303:11286]));
  assign MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_605_nl = (readslicef_28_18_10((MultLoop_627_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_628_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_605_nl = nl_MultLoop_acc_605_nl[17:0];
  assign nl_MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[11321:11304]));
  assign MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[11339:11322]));
  assign MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_604_nl = (readslicef_28_18_10((MultLoop_629_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_630_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_604_nl = nl_MultLoop_acc_604_nl[17:0];
  assign nl_MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[11429:11412]));
  assign MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[11447:11430]));
  assign MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_601_nl = (readslicef_28_18_10((MultLoop_635_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_636_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_601_nl = nl_MultLoop_acc_601_nl[17:0];
  assign nl_MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[11465:11448]));
  assign MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[11483:11466]));
  assign MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_600_nl = (readslicef_28_18_10((MultLoop_637_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_638_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_600_nl = nl_MultLoop_acc_600_nl[17:0];
  assign nl_MultLoop_acc_628_nl = (MultLoop_acc_603_nl) + (MultLoop_acc_602_nl) +
      (MultLoop_acc_607_nl) + (MultLoop_acc_606_nl) + (MultLoop_acc_605_nl) + (MultLoop_acc_604_nl)
      + (MultLoop_acc_601_nl) + (MultLoop_acc_600_nl);
  assign MultLoop_acc_628_nl = nl_MultLoop_acc_628_nl[17:0];
  assign nl_res_rsci_d_251_234  = (MultLoop_acc_629_nl) + (MultLoop_acc_628_nl);
  assign nl_MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[8909:8892]));
  assign MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[8927:8910]));
  assign MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_740_nl = (readslicef_28_18_10((MultLoop_495_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_496_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_740_nl = nl_MultLoop_acc_740_nl[17:0];
  assign nl_MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[8945:8928]));
  assign MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[8963:8946]));
  assign MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_739_nl = (readslicef_28_18_10((MultLoop_497_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_498_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_739_nl = nl_MultLoop_acc_739_nl[17:0];
  assign nl_MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[8981:8964]));
  assign MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[8999:8982]));
  assign MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_738_nl = (readslicef_28_18_10((MultLoop_499_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_500_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_738_nl = nl_MultLoop_acc_738_nl[17:0];
  assign nl_MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[9017:9000]));
  assign MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[9035:9018]));
  assign MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_737_nl = (readslicef_28_18_10((MultLoop_501_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_502_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_737_nl = nl_MultLoop_acc_737_nl[17:0];
  assign nl_MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[9053:9036]));
  assign MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[9071:9054]));
  assign MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_736_nl = (readslicef_28_18_10((MultLoop_503_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_504_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_736_nl = nl_MultLoop_acc_736_nl[17:0];
  assign nl_MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[9089:9072]));
  assign MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[9107:9090]));
  assign MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_735_nl = (readslicef_28_18_10((MultLoop_505_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_506_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_735_nl = nl_MultLoop_acc_735_nl[17:0];
  assign nl_MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[9125:9108]));
  assign MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[9143:9126]));
  assign MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_734_nl = (readslicef_28_18_10((MultLoop_507_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_508_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_734_nl = nl_MultLoop_acc_734_nl[17:0];
  assign nl_MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[9161:9144]));
  assign MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[9179:9162]));
  assign MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_733_nl = (readslicef_28_18_10((MultLoop_509_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_510_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_733_nl = nl_MultLoop_acc_733_nl[17:0];
  assign nl_MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[9341:9324]));
  assign MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[9359:9342]));
  assign MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_728_nl = (readslicef_28_18_10((MultLoop_519_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_520_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_728_nl = nl_MultLoop_acc_728_nl[17:0];
  assign nl_MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[9377:9360]));
  assign MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[9395:9378]));
  assign MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_727_nl = (readslicef_28_18_10((MultLoop_521_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_522_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_727_nl = nl_MultLoop_acc_727_nl[17:0];
  assign nl_MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[9413:9396]));
  assign MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[9431:9414]));
  assign MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_726_nl = (readslicef_28_18_10((MultLoop_523_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_524_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_726_nl = nl_MultLoop_acc_726_nl[17:0];
  assign nl_MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[9449:9432]));
  assign MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[9467:9450]));
  assign MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_725_nl = (readslicef_28_18_10((MultLoop_525_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_526_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_725_nl = nl_MultLoop_acc_725_nl[17:0];
  assign nl_MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[9197:9180]));
  assign MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[9215:9198]));
  assign MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_732_nl = (readslicef_28_18_10((MultLoop_511_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_512_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_732_nl = nl_MultLoop_acc_732_nl[17:0];
  assign nl_MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[9233:9216]));
  assign MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[9251:9234]));
  assign MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_731_nl = (readslicef_28_18_10((MultLoop_513_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_514_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_731_nl = nl_MultLoop_acc_731_nl[17:0];
  assign nl_MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[9269:9252]));
  assign MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[9287:9270]));
  assign MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_730_nl = (readslicef_28_18_10((MultLoop_515_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_516_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_730_nl = nl_MultLoop_acc_730_nl[17:0];
  assign nl_MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[9305:9288]));
  assign MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[9323:9306]));
  assign MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_729_nl = (readslicef_28_18_10((MultLoop_517_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_518_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_729_nl = nl_MultLoop_acc_729_nl[17:0];
  assign nl_MultLoop_acc_770_nl = (MultLoop_acc_740_nl) + (MultLoop_acc_739_nl) +
      (MultLoop_acc_738_nl) + (MultLoop_acc_737_nl) + (MultLoop_acc_736_nl) + (MultLoop_acc_735_nl)
      + (MultLoop_acc_734_nl) + (MultLoop_acc_733_nl) + (MultLoop_acc_728_nl) + (MultLoop_acc_727_nl)
      + (MultLoop_acc_726_nl) + (MultLoop_acc_725_nl) + (MultLoop_acc_732_nl) + (MultLoop_acc_731_nl)
      + (MultLoop_acc_730_nl) + (MultLoop_acc_729_nl);
  assign MultLoop_acc_770_nl = nl_MultLoop_acc_770_nl[17:0];
  assign nl_MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[8765:8748]));
  assign MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[8783:8766]));
  assign MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_744_nl = (readslicef_28_18_10((MultLoop_487_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_488_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_744_nl = nl_MultLoop_acc_744_nl[17:0];
  assign nl_MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[8801:8784]));
  assign MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[8819:8802]));
  assign MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_743_nl = (readslicef_28_18_10((MultLoop_489_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_490_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_743_nl = nl_MultLoop_acc_743_nl[17:0];
  assign nl_MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[9485:9468]));
  assign MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[9503:9486]));
  assign MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_724_nl = (readslicef_28_18_10((MultLoop_527_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_528_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_724_nl = nl_MultLoop_acc_724_nl[17:0];
  assign nl_MultLoop_acc_748_nl = (MultLoop_acc_724_nl) + (biases_rsci_idat[197:180]);
  assign MultLoop_acc_748_nl = nl_MultLoop_acc_748_nl[17:0];
  assign nl_MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[8657:8640]));
  assign MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[8675:8658]));
  assign MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_747_nl = (readslicef_28_18_10((MultLoop_481_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_482_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_747_nl = nl_MultLoop_acc_747_nl[17:0];
  assign nl_MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[8693:8676]));
  assign MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[8711:8694]));
  assign MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_746_nl = (readslicef_28_18_10((MultLoop_483_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_484_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_746_nl = nl_MultLoop_acc_746_nl[17:0];
  assign nl_MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[8729:8712]));
  assign MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[8747:8730]));
  assign MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_745_nl = (readslicef_28_18_10((MultLoop_485_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_486_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_745_nl = nl_MultLoop_acc_745_nl[17:0];
  assign nl_MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[8837:8820]));
  assign MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[8855:8838]));
  assign MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_742_nl = (readslicef_28_18_10((MultLoop_491_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_492_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_742_nl = nl_MultLoop_acc_742_nl[17:0];
  assign nl_MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[8873:8856]));
  assign MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[8891:8874]));
  assign MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_741_nl = (readslicef_28_18_10((MultLoop_493_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_494_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_741_nl = nl_MultLoop_acc_741_nl[17:0];
  assign nl_MultLoop_acc_769_nl = (MultLoop_acc_744_nl) + (MultLoop_acc_743_nl) +
      (MultLoop_acc_748_nl) + (MultLoop_acc_747_nl) + (MultLoop_acc_746_nl) + (MultLoop_acc_745_nl)
      + (MultLoop_acc_742_nl) + (MultLoop_acc_741_nl);
  assign MultLoop_acc_769_nl = nl_MultLoop_acc_769_nl[17:0];
  assign nl_res_rsci_d_197_180  = (MultLoop_acc_770_nl) + (MultLoop_acc_769_nl);
  assign nl_MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[10637:10620]));
  assign MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[10655:10638]));
  assign MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_646_nl = (readslicef_28_18_10((MultLoop_591_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_592_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_646_nl = nl_MultLoop_acc_646_nl[17:0];
  assign nl_MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[10673:10656]));
  assign MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[10691:10674]));
  assign MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_645_nl = (readslicef_28_18_10((MultLoop_593_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_594_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_645_nl = nl_MultLoop_acc_645_nl[17:0];
  assign nl_MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[10709:10692]));
  assign MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[10727:10710]));
  assign MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_644_nl = (readslicef_28_18_10((MultLoop_595_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_596_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_644_nl = nl_MultLoop_acc_644_nl[17:0];
  assign nl_MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[10745:10728]));
  assign MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[10763:10746]));
  assign MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_643_nl = (readslicef_28_18_10((MultLoop_597_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_598_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_643_nl = nl_MultLoop_acc_643_nl[17:0];
  assign nl_MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[10781:10764]));
  assign MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[10799:10782]));
  assign MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_642_nl = (readslicef_28_18_10((MultLoop_599_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_600_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_642_nl = nl_MultLoop_acc_642_nl[17:0];
  assign nl_MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[10817:10800]));
  assign MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[10835:10818]));
  assign MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_641_nl = (readslicef_28_18_10((MultLoop_601_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_602_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_641_nl = nl_MultLoop_acc_641_nl[17:0];
  assign nl_MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[10853:10836]));
  assign MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[10871:10854]));
  assign MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_640_nl = (readslicef_28_18_10((MultLoop_603_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_604_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_640_nl = nl_MultLoop_acc_640_nl[17:0];
  assign nl_MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[10889:10872]));
  assign MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[10907:10890]));
  assign MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_639_nl = (readslicef_28_18_10((MultLoop_605_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_606_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_639_nl = nl_MultLoop_acc_639_nl[17:0];
  assign nl_MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[11069:11052]));
  assign MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[11087:11070]));
  assign MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_634_nl = (readslicef_28_18_10((MultLoop_615_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_616_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_634_nl = nl_MultLoop_acc_634_nl[17:0];
  assign nl_MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[11105:11088]));
  assign MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[11123:11106]));
  assign MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_633_nl = (readslicef_28_18_10((MultLoop_617_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_618_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_633_nl = nl_MultLoop_acc_633_nl[17:0];
  assign nl_MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[11141:11124]));
  assign MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[11159:11142]));
  assign MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_632_nl = (readslicef_28_18_10((MultLoop_619_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_620_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_632_nl = nl_MultLoop_acc_632_nl[17:0];
  assign nl_MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[11177:11160]));
  assign MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[11195:11178]));
  assign MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_631_nl = (readslicef_28_18_10((MultLoop_621_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_622_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_631_nl = nl_MultLoop_acc_631_nl[17:0];
  assign nl_MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[10925:10908]));
  assign MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[10943:10926]));
  assign MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_638_nl = (readslicef_28_18_10((MultLoop_607_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_608_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_638_nl = nl_MultLoop_acc_638_nl[17:0];
  assign nl_MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[10961:10944]));
  assign MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[10979:10962]));
  assign MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_637_nl = (readslicef_28_18_10((MultLoop_609_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_610_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_637_nl = nl_MultLoop_acc_637_nl[17:0];
  assign nl_MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[10997:10980]));
  assign MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[11015:10998]));
  assign MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_636_nl = (readslicef_28_18_10((MultLoop_611_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_612_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_636_nl = nl_MultLoop_acc_636_nl[17:0];
  assign nl_MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[11033:11016]));
  assign MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[11051:11034]));
  assign MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_635_nl = (readslicef_28_18_10((MultLoop_613_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_614_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_635_nl = nl_MultLoop_acc_635_nl[17:0];
  assign nl_MultLoop_acc_676_nl = (MultLoop_acc_646_nl) + (MultLoop_acc_645_nl) +
      (MultLoop_acc_644_nl) + (MultLoop_acc_643_nl) + (MultLoop_acc_642_nl) + (MultLoop_acc_641_nl)
      + (MultLoop_acc_640_nl) + (MultLoop_acc_639_nl) + (MultLoop_acc_634_nl) + (MultLoop_acc_633_nl)
      + (MultLoop_acc_632_nl) + (MultLoop_acc_631_nl) + (MultLoop_acc_638_nl) + (MultLoop_acc_637_nl)
      + (MultLoop_acc_636_nl) + (MultLoop_acc_635_nl);
  assign MultLoop_acc_676_nl = nl_MultLoop_acc_676_nl[17:0];
  assign nl_MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[10493:10476]));
  assign MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[10511:10494]));
  assign MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_650_nl = (readslicef_28_18_10((MultLoop_583_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_584_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_650_nl = nl_MultLoop_acc_650_nl[17:0];
  assign nl_MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[10529:10512]));
  assign MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[10547:10530]));
  assign MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_649_nl = (readslicef_28_18_10((MultLoop_585_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_586_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_649_nl = nl_MultLoop_acc_649_nl[17:0];
  assign nl_MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[11213:11196]));
  assign MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[11231:11214]));
  assign MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_630_nl = (readslicef_28_18_10((MultLoop_623_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_624_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_630_nl = nl_MultLoop_acc_630_nl[17:0];
  assign nl_MultLoop_acc_654_nl = (MultLoop_acc_630_nl) + (biases_rsci_idat[233:216]);
  assign MultLoop_acc_654_nl = nl_MultLoop_acc_654_nl[17:0];
  assign nl_MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[10385:10368]));
  assign MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[10403:10386]));
  assign MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_653_nl = (readslicef_28_18_10((MultLoop_577_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_578_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_653_nl = nl_MultLoop_acc_653_nl[17:0];
  assign nl_MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[10421:10404]));
  assign MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[10439:10422]));
  assign MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_652_nl = (readslicef_28_18_10((MultLoop_579_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_580_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_652_nl = nl_MultLoop_acc_652_nl[17:0];
  assign nl_MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[10457:10440]));
  assign MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[10475:10458]));
  assign MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_651_nl = (readslicef_28_18_10((MultLoop_581_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_582_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_651_nl = nl_MultLoop_acc_651_nl[17:0];
  assign nl_MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[10565:10548]));
  assign MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[10583:10566]));
  assign MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_648_nl = (readslicef_28_18_10((MultLoop_587_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_588_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_648_nl = nl_MultLoop_acc_648_nl[17:0];
  assign nl_MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[10601:10584]));
  assign MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[10619:10602]));
  assign MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_647_nl = (readslicef_28_18_10((MultLoop_589_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_590_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_647_nl = nl_MultLoop_acc_647_nl[17:0];
  assign nl_MultLoop_acc_675_nl = (MultLoop_acc_650_nl) + (MultLoop_acc_649_nl) +
      (MultLoop_acc_654_nl) + (MultLoop_acc_653_nl) + (MultLoop_acc_652_nl) + (MultLoop_acc_651_nl)
      + (MultLoop_acc_648_nl) + (MultLoop_acc_647_nl);
  assign MultLoop_acc_675_nl = nl_MultLoop_acc_675_nl[17:0];
  assign nl_res_rsci_d_233_216  = (MultLoop_acc_676_nl) + (MultLoop_acc_675_nl);
  assign nl_MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[269:252])) * $signed((weights_rsci_idat[9773:9756]));
  assign MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[287:270])) * $signed((weights_rsci_idat[9791:9774]));
  assign MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_693_nl = (readslicef_28_18_10((MultLoop_543_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_544_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_693_nl = nl_MultLoop_acc_693_nl[17:0];
  assign nl_MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[305:288])) * $signed((weights_rsci_idat[9809:9792]));
  assign MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[323:306])) * $signed((weights_rsci_idat[9827:9810]));
  assign MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_692_nl = (readslicef_28_18_10((MultLoop_545_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_546_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_692_nl = nl_MultLoop_acc_692_nl[17:0];
  assign nl_MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[341:324])) * $signed((weights_rsci_idat[9845:9828]));
  assign MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[359:342])) * $signed((weights_rsci_idat[9863:9846]));
  assign MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_691_nl = (readslicef_28_18_10((MultLoop_547_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_548_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_691_nl = nl_MultLoop_acc_691_nl[17:0];
  assign nl_MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[377:360])) * $signed((weights_rsci_idat[9881:9864]));
  assign MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[395:378])) * $signed((weights_rsci_idat[9899:9882]));
  assign MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_690_nl = (readslicef_28_18_10((MultLoop_549_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_550_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_690_nl = nl_MultLoop_acc_690_nl[17:0];
  assign nl_MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[413:396])) * $signed((weights_rsci_idat[9917:9900]));
  assign MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[431:414])) * $signed((weights_rsci_idat[9935:9918]));
  assign MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_689_nl = (readslicef_28_18_10((MultLoop_551_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_552_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_689_nl = nl_MultLoop_acc_689_nl[17:0];
  assign nl_MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[449:432])) * $signed((weights_rsci_idat[9953:9936]));
  assign MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[467:450])) * $signed((weights_rsci_idat[9971:9954]));
  assign MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_688_nl = (readslicef_28_18_10((MultLoop_553_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_554_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_688_nl = nl_MultLoop_acc_688_nl[17:0];
  assign nl_MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[485:468])) * $signed((weights_rsci_idat[9989:9972]));
  assign MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[503:486])) * $signed((weights_rsci_idat[10007:9990]));
  assign MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_687_nl = (readslicef_28_18_10((MultLoop_555_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_556_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_687_nl = nl_MultLoop_acc_687_nl[17:0];
  assign nl_MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[521:504])) * $signed((weights_rsci_idat[10025:10008]));
  assign MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[539:522])) * $signed((weights_rsci_idat[10043:10026]));
  assign MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_686_nl = (readslicef_28_18_10((MultLoop_557_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_558_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_686_nl = nl_MultLoop_acc_686_nl[17:0];
  assign nl_MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[701:684])) * $signed((weights_rsci_idat[10205:10188]));
  assign MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[719:702])) * $signed((weights_rsci_idat[10223:10206]));
  assign MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_681_nl = (readslicef_28_18_10((MultLoop_567_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_568_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_681_nl = nl_MultLoop_acc_681_nl[17:0];
  assign nl_MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[737:720])) * $signed((weights_rsci_idat[10241:10224]));
  assign MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[755:738])) * $signed((weights_rsci_idat[10259:10242]));
  assign MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_680_nl = (readslicef_28_18_10((MultLoop_569_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_570_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_680_nl = nl_MultLoop_acc_680_nl[17:0];
  assign nl_MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[773:756])) * $signed((weights_rsci_idat[10277:10260]));
  assign MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[791:774])) * $signed((weights_rsci_idat[10295:10278]));
  assign MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_679_nl = (readslicef_28_18_10((MultLoop_571_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_572_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_679_nl = nl_MultLoop_acc_679_nl[17:0];
  assign nl_MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[809:792])) * $signed((weights_rsci_idat[10313:10296]));
  assign MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[827:810])) * $signed((weights_rsci_idat[10331:10314]));
  assign MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_678_nl = (readslicef_28_18_10((MultLoop_573_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_574_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_678_nl = nl_MultLoop_acc_678_nl[17:0];
  assign nl_MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[557:540])) * $signed((weights_rsci_idat[10061:10044]));
  assign MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[575:558])) * $signed((weights_rsci_idat[10079:10062]));
  assign MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_685_nl = (readslicef_28_18_10((MultLoop_559_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_560_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_685_nl = nl_MultLoop_acc_685_nl[17:0];
  assign nl_MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[593:576])) * $signed((weights_rsci_idat[10097:10080]));
  assign MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[611:594])) * $signed((weights_rsci_idat[10115:10098]));
  assign MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_684_nl = (readslicef_28_18_10((MultLoop_561_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_562_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_684_nl = nl_MultLoop_acc_684_nl[17:0];
  assign nl_MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[629:612])) * $signed((weights_rsci_idat[10133:10116]));
  assign MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[647:630])) * $signed((weights_rsci_idat[10151:10134]));
  assign MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_683_nl = (readslicef_28_18_10((MultLoop_563_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_564_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_683_nl = nl_MultLoop_acc_683_nl[17:0];
  assign nl_MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[665:648])) * $signed((weights_rsci_idat[10169:10152]));
  assign MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[683:666])) * $signed((weights_rsci_idat[10187:10170]));
  assign MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_682_nl = (readslicef_28_18_10((MultLoop_565_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_566_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_682_nl = nl_MultLoop_acc_682_nl[17:0];
  assign nl_MultLoop_acc_723_nl = (MultLoop_acc_693_nl) + (MultLoop_acc_692_nl) +
      (MultLoop_acc_691_nl) + (MultLoop_acc_690_nl) + (MultLoop_acc_689_nl) + (MultLoop_acc_688_nl)
      + (MultLoop_acc_687_nl) + (MultLoop_acc_686_nl) + (MultLoop_acc_681_nl) + (MultLoop_acc_680_nl)
      + (MultLoop_acc_679_nl) + (MultLoop_acc_678_nl) + (MultLoop_acc_685_nl) + (MultLoop_acc_684_nl)
      + (MultLoop_acc_683_nl) + (MultLoop_acc_682_nl);
  assign MultLoop_acc_723_nl = nl_MultLoop_acc_723_nl[17:0];
  assign nl_MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[125:108])) * $signed((weights_rsci_idat[9629:9612]));
  assign MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[143:126])) * $signed((weights_rsci_idat[9647:9630]));
  assign MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_697_nl = (readslicef_28_18_10((MultLoop_535_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_536_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_697_nl = nl_MultLoop_acc_697_nl[17:0];
  assign nl_MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[161:144])) * $signed((weights_rsci_idat[9665:9648]));
  assign MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[179:162])) * $signed((weights_rsci_idat[9683:9666]));
  assign MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_696_nl = (readslicef_28_18_10((MultLoop_537_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_538_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_696_nl = nl_MultLoop_acc_696_nl[17:0];
  assign nl_MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[845:828])) * $signed((weights_rsci_idat[10349:10332]));
  assign MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[863:846])) * $signed((weights_rsci_idat[10367:10350]));
  assign MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_677_nl = (readslicef_28_18_10((MultLoop_575_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_576_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_677_nl = nl_MultLoop_acc_677_nl[17:0];
  assign nl_MultLoop_acc_701_nl = (MultLoop_acc_677_nl) + (biases_rsci_idat[215:198]);
  assign MultLoop_acc_701_nl = nl_MultLoop_acc_701_nl[17:0];
  assign nl_MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[17:0])) * $signed((weights_rsci_idat[9521:9504]));
  assign MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[35:18])) * $signed((weights_rsci_idat[9539:9522]));
  assign MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_700_nl = (readslicef_28_18_10((MultLoop_529_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_530_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_700_nl = nl_MultLoop_acc_700_nl[17:0];
  assign nl_MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[53:36])) * $signed((weights_rsci_idat[9557:9540]));
  assign MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[71:54])) * $signed((weights_rsci_idat[9575:9558]));
  assign MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_699_nl = (readslicef_28_18_10((MultLoop_531_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_532_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_699_nl = nl_MultLoop_acc_699_nl[17:0];
  assign nl_MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[89:72])) * $signed((weights_rsci_idat[9593:9576]));
  assign MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[107:90])) * $signed((weights_rsci_idat[9611:9594]));
  assign MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_698_nl = (readslicef_28_18_10((MultLoop_533_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_534_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_698_nl = nl_MultLoop_acc_698_nl[17:0];
  assign nl_MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[197:180])) * $signed((weights_rsci_idat[9701:9684]));
  assign MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[215:198])) * $signed((weights_rsci_idat[9719:9702]));
  assign MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_695_nl = (readslicef_28_18_10((MultLoop_539_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_540_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_695_nl = nl_MultLoop_acc_695_nl[17:0];
  assign nl_MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[233:216])) * $signed((weights_rsci_idat[9737:9720]));
  assign MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = $signed((data_rsci_idat[251:234])) * $signed((weights_rsci_idat[9755:9738]));
  assign MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl
      = nl_MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl[27:0];
  assign nl_MultLoop_acc_694_nl = (readslicef_28_18_10((MultLoop_541_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)))
      + (readslicef_28_18_10((MultLoop_542_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_nl)));
  assign MultLoop_acc_694_nl = nl_MultLoop_acc_694_nl[17:0];
  assign nl_MultLoop_acc_722_nl = (MultLoop_acc_697_nl) + (MultLoop_acc_696_nl) +
      (MultLoop_acc_701_nl) + (MultLoop_acc_700_nl) + (MultLoop_acc_699_nl) + (MultLoop_acc_698_nl)
      + (MultLoop_acc_695_nl) + (MultLoop_acc_694_nl);
  assign MultLoop_acc_722_nl = nl_MultLoop_acc_722_nl[17:0];
  assign nl_res_rsci_d_215_198  = (MultLoop_acc_723_nl) + (MultLoop_acc_722_nl);

  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2 (
  data_rsc_dat, res_rsc_z, weights_rsc_dat, biases_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [863:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input [20735:0] weights_rsc_dat;
  input [431:0] biases_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_input_t_layer2_t_config2_core nnet_dense_large_input_t_layer2_t_config2_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .weights_rsc_dat(weights_rsc_dat),
      .biases_rsc_dat(biases_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Mon Feb 24 18:01:58 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    econV0_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module econV0_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;


  // FSM State Type Declaration for econV0_core_core_fsm_1
  parameter
    core_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : econV0_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 9'b000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 9'b000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 9'b000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 9'b000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 9'b001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 9'b010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 9'b100000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_staller
// ------------------------------------------------------------------


module econV0_core_staller (
  clk, rst, core_wen, core_wten, input_48_rsci_wen_comp, layer7_out_rsci_wen_comp,
      w2_rsci_wen_comp, b2_rsci_wen_comp, w4_rsci_wen_comp, b4_rsci_wen_comp, w6_rsci_wen_comp,
      b6_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_48_rsci_wen_comp;
  input layer7_out_rsci_wen_comp;
  input w2_rsci_wen_comp;
  input b2_rsci_wen_comp;
  input w4_rsci_wen_comp;
  input b4_rsci_wen_comp;
  input w6_rsci_wen_comp;
  input b6_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_48_rsci_wen_comp & layer7_out_rsci_wen_comp & w2_rsci_wen_comp
      & b2_rsci_wen_comp & w4_rsci_wen_comp & b4_rsci_wen_comp & w6_rsci_wen_comp
      & b6_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b6_rsc_triosy_obj_b6_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b6_rsc_triosy_obj_b6_rsc_triosy_wait_ctrl (
  core_wten, b6_rsc_triosy_obj_iswt0, b6_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b6_rsc_triosy_obj_iswt0;
  output b6_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b6_rsc_triosy_obj_ld_core_sct = b6_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w6_rsc_triosy_obj_w6_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w6_rsc_triosy_obj_w6_rsc_triosy_wait_ctrl (
  core_wten, w6_rsc_triosy_obj_iswt0, w6_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w6_rsc_triosy_obj_iswt0;
  output w6_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w6_rsc_triosy_obj_ld_core_sct = w6_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl (
  core_wten, b4_rsc_triosy_obj_iswt0, b4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;
  output b4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b4_rsc_triosy_obj_ld_core_sct = b4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl (
  core_wten, w4_rsc_triosy_obj_iswt0, w4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;
  output w4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w4_rsc_triosy_obj_ld_core_sct = w4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl (
  core_wten, b2_rsc_triosy_obj_iswt0, b2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;
  output b2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b2_rsc_triosy_obj_ld_core_sct = b2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl (
  core_wten, w2_rsc_triosy_obj_iswt0, w2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;
  output w2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w2_rsc_triosy_obj_ld_core_sct = w2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_out_1_rsc_triosy_obj_iswt0, const_size_out_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;
  output const_size_out_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsc_triosy_obj_ld_core_sct = const_size_out_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_in_1_rsc_triosy_obj_iswt0, const_size_in_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;
  output const_size_in_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsc_triosy_obj_ld_core_sct = const_size_in_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl (
  core_wten, layer7_out_rsc_triosy_obj_iswt0, layer7_out_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input layer7_out_rsc_triosy_obj_iswt0;
  output layer7_out_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsc_triosy_obj_ld_core_sct = layer7_out_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl (
  core_wten, input_48_rsc_triosy_obj_iswt0, input_48_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input input_48_rsc_triosy_obj_iswt0;
  output input_48_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsc_triosy_obj_ld_core_sct = input_48_rsc_triosy_obj_iswt0 & (~
      core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b6_rsci_b6_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_b6_rsci_b6_rsc_wait_dp (
  clk, rst, b6_rsci_oswt, b6_rsci_wen_comp, b6_rsci_idat_mxwt, b6_rsci_biwt, b6_rsci_bdwt,
      b6_rsci_bcwt, b6_rsci_idat
);
  input clk;
  input rst;
  input b6_rsci_oswt;
  output b6_rsci_wen_comp;
  output [53:0] b6_rsci_idat_mxwt;
  input b6_rsci_biwt;
  input b6_rsci_bdwt;
  output b6_rsci_bcwt;
  reg b6_rsci_bcwt;
  input [53:0] b6_rsci_idat;


  // Interconnect Declarations
  reg [53:0] b6_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign b6_rsci_wen_comp = (~ b6_rsci_oswt) | b6_rsci_biwt | b6_rsci_bcwt;
  assign b6_rsci_idat_mxwt = MUX_v_54_2_2(b6_rsci_idat, b6_rsci_idat_bfwt, b6_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      b6_rsci_bcwt <= 1'b0;
    end
    else begin
      b6_rsci_bcwt <= ~((~(b6_rsci_bcwt | b6_rsci_biwt)) | b6_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      b6_rsci_idat_bfwt <= 54'b000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ b6_rsci_bcwt ) begin
      b6_rsci_idat_bfwt <= b6_rsci_idat_mxwt;
    end
  end

  function automatic [53:0] MUX_v_54_2_2;
    input [53:0] input_0;
    input [53:0] input_1;
    input [0:0] sel;
    reg [53:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_54_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b6_rsci_b6_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b6_rsci_b6_rsc_wait_ctrl (
  core_wen, b6_rsci_oswt, b6_rsci_biwt, b6_rsci_bdwt, b6_rsci_bcwt, b6_rsci_irdy_core_sct,
      b6_rsci_ivld
);
  input core_wen;
  input b6_rsci_oswt;
  output b6_rsci_biwt;
  output b6_rsci_bdwt;
  input b6_rsci_bcwt;
  output b6_rsci_irdy_core_sct;
  input b6_rsci_ivld;


  // Interconnect Declarations
  wire b6_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b6_rsci_bdwt = b6_rsci_oswt & core_wen;
  assign b6_rsci_biwt = b6_rsci_ogwt & b6_rsci_ivld;
  assign b6_rsci_ogwt = b6_rsci_oswt & (~ b6_rsci_bcwt);
  assign b6_rsci_irdy_core_sct = b6_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w6_rsci_w6_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_w6_rsci_w6_rsc_wait_dp (
  clk, rst, w6_rsci_oswt, w6_rsci_wen_comp, w6_rsci_idat_mxwt, w6_rsci_biwt, w6_rsci_bdwt,
      w6_rsci_bcwt, w6_rsci_idat
);
  input clk;
  input rst;
  input w6_rsci_oswt;
  output w6_rsci_wen_comp;
  output [323:0] w6_rsci_idat_mxwt;
  input w6_rsci_biwt;
  input w6_rsci_bdwt;
  output w6_rsci_bcwt;
  reg w6_rsci_bcwt;
  input [323:0] w6_rsci_idat;


  // Interconnect Declarations
  reg [323:0] w6_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w6_rsci_wen_comp = (~ w6_rsci_oswt) | w6_rsci_biwt | w6_rsci_bcwt;
  assign w6_rsci_idat_mxwt = MUX_v_324_2_2(w6_rsci_idat, w6_rsci_idat_bfwt, w6_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      w6_rsci_bcwt <= 1'b0;
    end
    else begin
      w6_rsci_bcwt <= ~((~(w6_rsci_bcwt | w6_rsci_biwt)) | w6_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w6_rsci_idat_bfwt <= 324'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ w6_rsci_bcwt ) begin
      w6_rsci_idat_bfwt <= w6_rsci_idat_mxwt;
    end
  end

  function automatic [323:0] MUX_v_324_2_2;
    input [323:0] input_0;
    input [323:0] input_1;
    input [0:0] sel;
    reg [323:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_324_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w6_rsci_w6_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w6_rsci_w6_rsc_wait_ctrl (
  core_wen, w6_rsci_oswt, w6_rsci_biwt, w6_rsci_bdwt, w6_rsci_bcwt, w6_rsci_irdy_core_sct,
      w6_rsci_ivld
);
  input core_wen;
  input w6_rsci_oswt;
  output w6_rsci_biwt;
  output w6_rsci_bdwt;
  input w6_rsci_bcwt;
  output w6_rsci_irdy_core_sct;
  input w6_rsci_ivld;


  // Interconnect Declarations
  wire w6_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w6_rsci_bdwt = w6_rsci_oswt & core_wen;
  assign w6_rsci_biwt = w6_rsci_ogwt & w6_rsci_ivld;
  assign w6_rsci_ogwt = w6_rsci_oswt & (~ w6_rsci_bcwt);
  assign w6_rsci_irdy_core_sct = w6_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b4_rsci_b4_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_b4_rsci_b4_rsc_wait_dp (
  clk, rst, b4_rsci_oswt, b4_rsci_wen_comp, b4_rsci_idat_mxwt, b4_rsci_biwt, b4_rsci_bdwt,
      b4_rsci_bcwt, b4_rsci_idat
);
  input clk;
  input rst;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [107:0] b4_rsci_idat_mxwt;
  input b4_rsci_biwt;
  input b4_rsci_bdwt;
  output b4_rsci_bcwt;
  reg b4_rsci_bcwt;
  input [107:0] b4_rsci_idat;


  // Interconnect Declarations
  reg [107:0] b4_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign b4_rsci_wen_comp = (~ b4_rsci_oswt) | b4_rsci_biwt | b4_rsci_bcwt;
  assign b4_rsci_idat_mxwt = MUX_v_108_2_2(b4_rsci_idat, b4_rsci_idat_bfwt, b4_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      b4_rsci_bcwt <= 1'b0;
    end
    else begin
      b4_rsci_bcwt <= ~((~(b4_rsci_bcwt | b4_rsci_biwt)) | b4_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      b4_rsci_idat_bfwt <= 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ b4_rsci_bcwt ) begin
      b4_rsci_idat_bfwt <= b4_rsci_idat_mxwt;
    end
  end

  function automatic [107:0] MUX_v_108_2_2;
    input [107:0] input_0;
    input [107:0] input_1;
    input [0:0] sel;
    reg [107:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_108_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b4_rsci_b4_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b4_rsci_b4_rsc_wait_ctrl (
  core_wen, b4_rsci_oswt, b4_rsci_biwt, b4_rsci_bdwt, b4_rsci_bcwt, b4_rsci_irdy_core_sct,
      b4_rsci_ivld
);
  input core_wen;
  input b4_rsci_oswt;
  output b4_rsci_biwt;
  output b4_rsci_bdwt;
  input b4_rsci_bcwt;
  output b4_rsci_irdy_core_sct;
  input b4_rsci_ivld;


  // Interconnect Declarations
  wire b4_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b4_rsci_bdwt = b4_rsci_oswt & core_wen;
  assign b4_rsci_biwt = b4_rsci_ogwt & b4_rsci_ivld;
  assign b4_rsci_ogwt = b4_rsci_oswt & (~ b4_rsci_bcwt);
  assign b4_rsci_irdy_core_sct = b4_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w4_rsci_w4_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_w4_rsci_w4_rsc_wait_dp (
  clk, rst, w4_rsci_oswt, w4_rsci_wen_comp, w4_rsci_idat_mxwt, w4_rsci_biwt, w4_rsci_bdwt,
      w4_rsci_bcwt, w4_rsci_idat
);
  input clk;
  input rst;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [2591:0] w4_rsci_idat_mxwt;
  input w4_rsci_biwt;
  input w4_rsci_bdwt;
  output w4_rsci_bcwt;
  reg w4_rsci_bcwt;
  input [2591:0] w4_rsci_idat;


  // Interconnect Declarations
  reg [2591:0] w4_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w4_rsci_wen_comp = (~ w4_rsci_oswt) | w4_rsci_biwt | w4_rsci_bcwt;
  assign w4_rsci_idat_mxwt = MUX_v_2592_2_2(w4_rsci_idat, w4_rsci_idat_bfwt, w4_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_bcwt <= 1'b0;
    end
    else begin
      w4_rsci_bcwt <= ~((~(w4_rsci_bcwt | w4_rsci_biwt)) | w4_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_idat_bfwt <= {648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( ~ w4_rsci_bcwt ) begin
      w4_rsci_idat_bfwt <= w4_rsci_idat_mxwt;
    end
  end

  function automatic [2591:0] MUX_v_2592_2_2;
    input [2591:0] input_0;
    input [2591:0] input_1;
    input [0:0] sel;
    reg [2591:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2592_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w4_rsci_w4_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w4_rsci_w4_rsc_wait_ctrl (
  core_wen, w4_rsci_oswt, w4_rsci_biwt, w4_rsci_bdwt, w4_rsci_bcwt, w4_rsci_irdy_core_sct,
      w4_rsci_ivld
);
  input core_wen;
  input w4_rsci_oswt;
  output w4_rsci_biwt;
  output w4_rsci_bdwt;
  input w4_rsci_bcwt;
  output w4_rsci_irdy_core_sct;
  input w4_rsci_ivld;


  // Interconnect Declarations
  wire w4_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w4_rsci_bdwt = w4_rsci_oswt & core_wen;
  assign w4_rsci_biwt = w4_rsci_ogwt & w4_rsci_ivld;
  assign w4_rsci_ogwt = w4_rsci_oswt & (~ w4_rsci_bcwt);
  assign w4_rsci_irdy_core_sct = w4_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b2_rsci_b2_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_b2_rsci_b2_rsc_wait_dp (
  clk, rst, b2_rsci_oswt, b2_rsci_wen_comp, b2_rsci_idat_mxwt, b2_rsci_biwt, b2_rsci_bdwt,
      b2_rsci_bcwt, b2_rsci_idat
);
  input clk;
  input rst;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [431:0] b2_rsci_idat_mxwt;
  input b2_rsci_biwt;
  input b2_rsci_bdwt;
  output b2_rsci_bcwt;
  reg b2_rsci_bcwt;
  input [431:0] b2_rsci_idat;


  // Interconnect Declarations
  reg [431:0] b2_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign b2_rsci_wen_comp = (~ b2_rsci_oswt) | b2_rsci_biwt | b2_rsci_bcwt;
  assign b2_rsci_idat_mxwt = MUX_v_432_2_2(b2_rsci_idat, b2_rsci_idat_bfwt, b2_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      b2_rsci_bcwt <= 1'b0;
      b2_rsci_idat_bfwt <= 432'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      b2_rsci_bcwt <= ~((~(b2_rsci_bcwt | b2_rsci_biwt)) | b2_rsci_bdwt);
      b2_rsci_idat_bfwt <= b2_rsci_idat_mxwt;
    end
  end

  function automatic [431:0] MUX_v_432_2_2;
    input [431:0] input_0;
    input [431:0] input_1;
    input [0:0] sel;
    reg [431:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_432_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b2_rsci_b2_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_b2_rsci_b2_rsc_wait_ctrl (
  core_wen, b2_rsci_oswt, b2_rsci_biwt, b2_rsci_bdwt, b2_rsci_bcwt, b2_rsci_irdy_core_sct,
      b2_rsci_ivld
);
  input core_wen;
  input b2_rsci_oswt;
  output b2_rsci_biwt;
  output b2_rsci_bdwt;
  input b2_rsci_bcwt;
  output b2_rsci_irdy_core_sct;
  input b2_rsci_ivld;


  // Interconnect Declarations
  wire b2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b2_rsci_bdwt = b2_rsci_oswt & core_wen;
  assign b2_rsci_biwt = b2_rsci_ogwt & b2_rsci_ivld;
  assign b2_rsci_ogwt = b2_rsci_oswt & (~ b2_rsci_bcwt);
  assign b2_rsci_irdy_core_sct = b2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w2_rsci_w2_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_w2_rsci_w2_rsc_wait_dp (
  clk, rst, w2_rsci_oswt, w2_rsci_wen_comp, w2_rsci_idat_mxwt, w2_rsci_biwt, w2_rsci_bdwt,
      w2_rsci_bcwt, w2_rsci_idat
);
  input clk;
  input rst;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [20735:0] w2_rsci_idat_mxwt;
  input w2_rsci_biwt;
  input w2_rsci_bdwt;
  output w2_rsci_bcwt;
  reg w2_rsci_bcwt;
  input [20735:0] w2_rsci_idat;


  // Interconnect Declarations
  reg [20735:0] w2_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w2_rsci_wen_comp = (~ w2_rsci_oswt) | w2_rsci_biwt | w2_rsci_bcwt;
  assign w2_rsci_idat_mxwt = MUX_v_20736_2_2(w2_rsci_idat, w2_rsci_idat_bfwt, w2_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_bcwt <= 1'b0;
      w2_rsci_idat_bfwt <= {648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else begin
      w2_rsci_bcwt <= ~((~(w2_rsci_bcwt | w2_rsci_biwt)) | w2_rsci_bdwt);
      w2_rsci_idat_bfwt <= w2_rsci_idat_mxwt;
    end
  end

  function automatic [20735:0] MUX_v_20736_2_2;
    input [20735:0] input_0;
    input [20735:0] input_1;
    input [0:0] sel;
    reg [20735:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20736_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w2_rsci_w2_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_w2_rsci_w2_rsc_wait_ctrl (
  core_wen, w2_rsci_oswt, w2_rsci_biwt, w2_rsci_bdwt, w2_rsci_bcwt, w2_rsci_irdy_core_sct,
      w2_rsci_ivld
);
  input core_wen;
  input w2_rsci_oswt;
  output w2_rsci_biwt;
  output w2_rsci_bdwt;
  input w2_rsci_bcwt;
  output w2_rsci_irdy_core_sct;
  input w2_rsci_ivld;


  // Interconnect Declarations
  wire w2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w2_rsci_bdwt = w2_rsci_oswt & core_wen;
  assign w2_rsci_biwt = w2_rsci_ogwt & w2_rsci_ivld;
  assign w2_rsci_ogwt = w2_rsci_oswt & (~ w2_rsci_bcwt);
  assign w2_rsci_irdy_core_sct = w2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wten, const_size_out_1_rsci_iswt0, const_size_out_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_out_1_rsci_iswt0;
  output const_size_out_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wten, const_size_in_1_rsci_iswt0, const_size_in_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_in_1_rsci_iswt0;
  output const_size_in_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp (
  clk, rst, layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_biwt,
      layer7_out_rsci_bdwt, layer7_out_rsci_bcwt
);
  input clk;
  input rst;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input layer7_out_rsci_biwt;
  input layer7_out_rsci_bdwt;
  output layer7_out_rsci_bcwt;
  reg layer7_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_wen_comp = (~ layer7_out_rsci_oswt) | layer7_out_rsci_biwt
      | layer7_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_bcwt <= 1'b0;
    end
    else begin
      layer7_out_rsci_bcwt <= ~((~(layer7_out_rsci_bcwt | layer7_out_rsci_biwt))
          | layer7_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl (
  core_wen, layer7_out_rsci_oswt, layer7_out_rsci_irdy, layer7_out_rsci_biwt, layer7_out_rsci_bdwt,
      layer7_out_rsci_bcwt, layer7_out_rsci_ivld_core_sct
);
  input core_wen;
  input layer7_out_rsci_oswt;
  input layer7_out_rsci_irdy;
  output layer7_out_rsci_biwt;
  output layer7_out_rsci_bdwt;
  input layer7_out_rsci_bcwt;
  output layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire layer7_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_bdwt = layer7_out_rsci_oswt & core_wen;
  assign layer7_out_rsci_biwt = layer7_out_rsci_ogwt & layer7_out_rsci_irdy;
  assign layer7_out_rsci_ogwt = layer7_out_rsci_oswt & (~ layer7_out_rsci_bcwt);
  assign layer7_out_rsci_ivld_core_sct = layer7_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci_input_48_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_input_48_rsci_input_48_rsc_wait_dp (
  clk, rst, input_48_rsci_oswt, input_48_rsci_wen_comp, input_48_rsci_idat_mxwt,
      input_48_rsci_biwt, input_48_rsci_bdwt, input_48_rsci_bcwt, input_48_rsci_idat
);
  input clk;
  input rst;
  input input_48_rsci_oswt;
  output input_48_rsci_wen_comp;
  output [863:0] input_48_rsci_idat_mxwt;
  input input_48_rsci_biwt;
  input input_48_rsci_bdwt;
  output input_48_rsci_bcwt;
  reg input_48_rsci_bcwt;
  input [863:0] input_48_rsci_idat;


  // Interconnect Declarations
  reg [863:0] input_48_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsci_wen_comp = (~ input_48_rsci_oswt) | input_48_rsci_biwt | input_48_rsci_bcwt;
  assign input_48_rsci_idat_mxwt = MUX_v_864_2_2(input_48_rsci_idat, input_48_rsci_idat_bfwt,
      input_48_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input_48_rsci_bcwt <= 1'b0;
      input_48_rsci_idat_bfwt <= 864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      input_48_rsci_bcwt <= ~((~(input_48_rsci_bcwt | input_48_rsci_biwt)) | input_48_rsci_bdwt);
      input_48_rsci_idat_bfwt <= input_48_rsci_idat_mxwt;
    end
  end

  function automatic [863:0] MUX_v_864_2_2;
    input [863:0] input_0;
    input [863:0] input_1;
    input [0:0] sel;
    reg [863:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_864_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci_input_48_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_input_48_rsci_input_48_rsc_wait_ctrl (
  core_wen, input_48_rsci_oswt, input_48_rsci_biwt, input_48_rsci_bdwt, input_48_rsci_bcwt,
      input_48_rsci_irdy_core_sct, input_48_rsci_ivld
);
  input core_wen;
  input input_48_rsci_oswt;
  output input_48_rsci_biwt;
  output input_48_rsci_bdwt;
  input input_48_rsci_bcwt;
  output input_48_rsci_irdy_core_sct;
  input input_48_rsci_ivld;


  // Interconnect Declarations
  wire input_48_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsci_bdwt = input_48_rsci_oswt & core_wen;
  assign input_48_rsci_biwt = input_48_rsci_ogwt & input_48_rsci_ivld;
  assign input_48_rsci_ogwt = input_48_rsci_oswt & (~ input_48_rsci_bcwt);
  assign input_48_rsci_irdy_core_sct = input_48_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b6_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_b6_rsc_triosy_obj (
  b6_rsc_triosy_lz, core_wten, b6_rsc_triosy_obj_iswt0
);
  output b6_rsc_triosy_lz;
  input core_wten;
  input b6_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b6_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b6_rsc_triosy_obj (
      .ld(b6_rsc_triosy_obj_ld_core_sct),
      .lz(b6_rsc_triosy_lz)
    );
  econV0_core_b6_rsc_triosy_obj_b6_rsc_triosy_wait_ctrl econV0_core_b6_rsc_triosy_obj_b6_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b6_rsc_triosy_obj_iswt0(b6_rsc_triosy_obj_iswt0),
      .b6_rsc_triosy_obj_ld_core_sct(b6_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w6_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_w6_rsc_triosy_obj (
  w6_rsc_triosy_lz, core_wten, w6_rsc_triosy_obj_iswt0
);
  output w6_rsc_triosy_lz;
  input core_wten;
  input w6_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w6_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w6_rsc_triosy_obj (
      .ld(w6_rsc_triosy_obj_ld_core_sct),
      .lz(w6_rsc_triosy_lz)
    );
  econV0_core_w6_rsc_triosy_obj_w6_rsc_triosy_wait_ctrl econV0_core_w6_rsc_triosy_obj_w6_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w6_rsc_triosy_obj_iswt0(w6_rsc_triosy_obj_iswt0),
      .w6_rsc_triosy_obj_ld_core_sct(w6_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b4_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_b4_rsc_triosy_obj (
  b4_rsc_triosy_lz, core_wten, b4_rsc_triosy_obj_iswt0
);
  output b4_rsc_triosy_lz;
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b4_rsc_triosy_obj (
      .ld(b4_rsc_triosy_obj_ld_core_sct),
      .lz(b4_rsc_triosy_lz)
    );
  econV0_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl econV0_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(b4_rsc_triosy_obj_iswt0),
      .b4_rsc_triosy_obj_ld_core_sct(b4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w4_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_w4_rsc_triosy_obj (
  w4_rsc_triosy_lz, core_wten, w4_rsc_triosy_obj_iswt0
);
  output w4_rsc_triosy_lz;
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w4_rsc_triosy_obj (
      .ld(w4_rsc_triosy_obj_ld_core_sct),
      .lz(w4_rsc_triosy_lz)
    );
  econV0_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl econV0_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(w4_rsc_triosy_obj_iswt0),
      .w4_rsc_triosy_obj_ld_core_sct(w4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b2_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_b2_rsc_triosy_obj (
  b2_rsc_triosy_lz, core_wten, b2_rsc_triosy_obj_iswt0
);
  output b2_rsc_triosy_lz;
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b2_rsc_triosy_obj (
      .ld(b2_rsc_triosy_obj_ld_core_sct),
      .lz(b2_rsc_triosy_lz)
    );
  econV0_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl econV0_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(b2_rsc_triosy_obj_iswt0),
      .b2_rsc_triosy_obj_ld_core_sct(b2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w2_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_w2_rsc_triosy_obj (
  w2_rsc_triosy_lz, core_wten, w2_rsc_triosy_obj_iswt0
);
  output w2_rsc_triosy_lz;
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w2_rsc_triosy_obj (
      .ld(w2_rsc_triosy_obj_ld_core_sct),
      .lz(w2_rsc_triosy_lz)
    );
  econV0_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl econV0_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(w2_rsc_triosy_obj_iswt0),
      .w2_rsc_triosy_obj_ld_core_sct(w2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsc_triosy_obj (
  const_size_out_1_rsc_triosy_lz, core_wten, const_size_out_1_rsc_triosy_obj_iswt0
);
  output const_size_out_1_rsc_triosy_lz;
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_out_1_rsc_triosy_obj (
      .ld(const_size_out_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_out_1_rsc_triosy_lz)
    );
  econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
      econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(const_size_out_1_rsc_triosy_obj_iswt0),
      .const_size_out_1_rsc_triosy_obj_ld_core_sct(const_size_out_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsc_triosy_obj (
  const_size_in_1_rsc_triosy_lz, core_wten, const_size_in_1_rsc_triosy_obj_iswt0
);
  output const_size_in_1_rsc_triosy_lz;
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_in_1_rsc_triosy_obj (
      .ld(const_size_in_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_in_1_rsc_triosy_lz)
    );
  econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
      econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(const_size_in_1_rsc_triosy_obj_iswt0),
      .const_size_in_1_rsc_triosy_obj_ld_core_sct(const_size_in_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsc_triosy_obj (
  layer7_out_rsc_triosy_lz, core_wten, layer7_out_rsc_triosy_obj_iswt0
);
  output layer7_out_rsc_triosy_lz;
  input core_wten;
  input layer7_out_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire layer7_out_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) layer7_out_rsc_triosy_obj (
      .ld(layer7_out_rsc_triosy_obj_ld_core_sct),
      .lz(layer7_out_rsc_triosy_lz)
    );
  econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer7_out_rsc_triosy_obj_iswt0(layer7_out_rsc_triosy_obj_iswt0),
      .layer7_out_rsc_triosy_obj_ld_core_sct(layer7_out_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_input_48_rsc_triosy_obj (
  input_48_rsc_triosy_lz, core_wten, input_48_rsc_triosy_obj_iswt0
);
  output input_48_rsc_triosy_lz;
  input core_wten;
  input input_48_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire input_48_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) input_48_rsc_triosy_obj (
      .ld(input_48_rsc_triosy_obj_ld_core_sct),
      .lz(input_48_rsc_triosy_lz)
    );
  econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .input_48_rsc_triosy_obj_iswt0(input_48_rsc_triosy_obj_iswt0),
      .input_48_rsc_triosy_obj_ld_core_sct(input_48_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b6_rsci
// ------------------------------------------------------------------


module econV0_core_b6_rsci (
  clk, rst, b6_rsc_dat, b6_rsc_vld, b6_rsc_rdy, core_wen, b6_rsci_oswt, b6_rsci_wen_comp,
      b6_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [53:0] b6_rsc_dat;
  input b6_rsc_vld;
  output b6_rsc_rdy;
  input core_wen;
  input b6_rsci_oswt;
  output b6_rsci_wen_comp;
  output [53:0] b6_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b6_rsci_biwt;
  wire b6_rsci_bdwt;
  wire b6_rsci_bcwt;
  wire b6_rsci_irdy_core_sct;
  wire b6_rsci_ivld;
  wire [53:0] b6_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd31),
  .width(32'sd54)) b6_rsci (
      .rdy(b6_rsc_rdy),
      .vld(b6_rsc_vld),
      .dat(b6_rsc_dat),
      .irdy(b6_rsci_irdy_core_sct),
      .ivld(b6_rsci_ivld),
      .idat(b6_rsci_idat)
    );
  econV0_core_b6_rsci_b6_rsc_wait_ctrl econV0_core_b6_rsci_b6_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .b6_rsci_oswt(b6_rsci_oswt),
      .b6_rsci_biwt(b6_rsci_biwt),
      .b6_rsci_bdwt(b6_rsci_bdwt),
      .b6_rsci_bcwt(b6_rsci_bcwt),
      .b6_rsci_irdy_core_sct(b6_rsci_irdy_core_sct),
      .b6_rsci_ivld(b6_rsci_ivld)
    );
  econV0_core_b6_rsci_b6_rsc_wait_dp econV0_core_b6_rsci_b6_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .b6_rsci_oswt(b6_rsci_oswt),
      .b6_rsci_wen_comp(b6_rsci_wen_comp),
      .b6_rsci_idat_mxwt(b6_rsci_idat_mxwt),
      .b6_rsci_biwt(b6_rsci_biwt),
      .b6_rsci_bdwt(b6_rsci_bdwt),
      .b6_rsci_bcwt(b6_rsci_bcwt),
      .b6_rsci_idat(b6_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w6_rsci
// ------------------------------------------------------------------


module econV0_core_w6_rsci (
  clk, rst, w6_rsc_dat, w6_rsc_vld, w6_rsc_rdy, core_wen, w6_rsci_oswt, w6_rsci_wen_comp,
      w6_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [323:0] w6_rsc_dat;
  input w6_rsc_vld;
  output w6_rsc_rdy;
  input core_wen;
  input w6_rsci_oswt;
  output w6_rsci_wen_comp;
  output [323:0] w6_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w6_rsci_biwt;
  wire w6_rsci_bdwt;
  wire w6_rsci_bcwt;
  wire w6_rsci_irdy_core_sct;
  wire w6_rsci_ivld;
  wire [323:0] w6_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd30),
  .width(32'sd324)) w6_rsci (
      .rdy(w6_rsc_rdy),
      .vld(w6_rsc_vld),
      .dat(w6_rsc_dat),
      .irdy(w6_rsci_irdy_core_sct),
      .ivld(w6_rsci_ivld),
      .idat(w6_rsci_idat)
    );
  econV0_core_w6_rsci_w6_rsc_wait_ctrl econV0_core_w6_rsci_w6_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .w6_rsci_oswt(w6_rsci_oswt),
      .w6_rsci_biwt(w6_rsci_biwt),
      .w6_rsci_bdwt(w6_rsci_bdwt),
      .w6_rsci_bcwt(w6_rsci_bcwt),
      .w6_rsci_irdy_core_sct(w6_rsci_irdy_core_sct),
      .w6_rsci_ivld(w6_rsci_ivld)
    );
  econV0_core_w6_rsci_w6_rsc_wait_dp econV0_core_w6_rsci_w6_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .w6_rsci_oswt(w6_rsci_oswt),
      .w6_rsci_wen_comp(w6_rsci_wen_comp),
      .w6_rsci_idat_mxwt(w6_rsci_idat_mxwt),
      .w6_rsci_biwt(w6_rsci_biwt),
      .w6_rsci_bdwt(w6_rsci_bdwt),
      .w6_rsci_bcwt(w6_rsci_bcwt),
      .w6_rsci_idat(w6_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b4_rsci
// ------------------------------------------------------------------


module econV0_core_b4_rsci (
  clk, rst, b4_rsc_dat, b4_rsc_vld, b4_rsc_rdy, core_wen, b4_rsci_oswt, b4_rsci_wen_comp,
      b4_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [107:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  input core_wen;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [107:0] b4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b4_rsci_biwt;
  wire b4_rsci_bdwt;
  wire b4_rsci_bcwt;
  wire b4_rsci_irdy_core_sct;
  wire b4_rsci_ivld;
  wire [107:0] b4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd29),
  .width(32'sd108)) b4_rsci (
      .rdy(b4_rsc_rdy),
      .vld(b4_rsc_vld),
      .dat(b4_rsc_dat),
      .irdy(b4_rsci_irdy_core_sct),
      .ivld(b4_rsci_ivld),
      .idat(b4_rsci_idat)
    );
  econV0_core_b4_rsci_b4_rsc_wait_ctrl econV0_core_b4_rsci_b4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .b4_rsci_oswt(b4_rsci_oswt),
      .b4_rsci_biwt(b4_rsci_biwt),
      .b4_rsci_bdwt(b4_rsci_bdwt),
      .b4_rsci_bcwt(b4_rsci_bcwt),
      .b4_rsci_irdy_core_sct(b4_rsci_irdy_core_sct),
      .b4_rsci_ivld(b4_rsci_ivld)
    );
  econV0_core_b4_rsci_b4_rsc_wait_dp econV0_core_b4_rsci_b4_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .b4_rsci_oswt(b4_rsci_oswt),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt),
      .b4_rsci_biwt(b4_rsci_biwt),
      .b4_rsci_bdwt(b4_rsci_bdwt),
      .b4_rsci_bcwt(b4_rsci_bcwt),
      .b4_rsci_idat(b4_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w4_rsci
// ------------------------------------------------------------------


module econV0_core_w4_rsci (
  clk, rst, w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, core_wen, w4_rsci_oswt, w4_rsci_wen_comp,
      w4_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [2591:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  input core_wen;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [2591:0] w4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w4_rsci_biwt;
  wire w4_rsci_bdwt;
  wire w4_rsci_bcwt;
  wire w4_rsci_irdy_core_sct;
  wire w4_rsci_ivld;
  wire [2591:0] w4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd28),
  .width(32'sd2592)) w4_rsci (
      .rdy(w4_rsc_rdy),
      .vld(w4_rsc_vld),
      .dat(w4_rsc_dat),
      .irdy(w4_rsci_irdy_core_sct),
      .ivld(w4_rsci_ivld),
      .idat(w4_rsci_idat)
    );
  econV0_core_w4_rsci_w4_rsc_wait_ctrl econV0_core_w4_rsci_w4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .w4_rsci_oswt(w4_rsci_oswt),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_bcwt(w4_rsci_bcwt),
      .w4_rsci_irdy_core_sct(w4_rsci_irdy_core_sct),
      .w4_rsci_ivld(w4_rsci_ivld)
    );
  econV0_core_w4_rsci_w4_rsc_wait_dp econV0_core_w4_rsci_w4_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .w4_rsci_oswt(w4_rsci_oswt),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_bcwt(w4_rsci_bcwt),
      .w4_rsci_idat(w4_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_b2_rsci
// ------------------------------------------------------------------


module econV0_core_b2_rsci (
  clk, rst, b2_rsc_dat, b2_rsc_vld, b2_rsc_rdy, core_wen, b2_rsci_oswt, b2_rsci_wen_comp,
      b2_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [431:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  input core_wen;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [431:0] b2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b2_rsci_biwt;
  wire b2_rsci_bdwt;
  wire b2_rsci_bcwt;
  wire b2_rsci_irdy_core_sct;
  wire b2_rsci_ivld;
  wire [431:0] b2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd27),
  .width(32'sd432)) b2_rsci (
      .rdy(b2_rsc_rdy),
      .vld(b2_rsc_vld),
      .dat(b2_rsc_dat),
      .irdy(b2_rsci_irdy_core_sct),
      .ivld(b2_rsci_ivld),
      .idat(b2_rsci_idat)
    );
  econV0_core_b2_rsci_b2_rsc_wait_ctrl econV0_core_b2_rsci_b2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .b2_rsci_oswt(b2_rsci_oswt),
      .b2_rsci_biwt(b2_rsci_biwt),
      .b2_rsci_bdwt(b2_rsci_bdwt),
      .b2_rsci_bcwt(b2_rsci_bcwt),
      .b2_rsci_irdy_core_sct(b2_rsci_irdy_core_sct),
      .b2_rsci_ivld(b2_rsci_ivld)
    );
  econV0_core_b2_rsci_b2_rsc_wait_dp econV0_core_b2_rsci_b2_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .b2_rsci_oswt(b2_rsci_oswt),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt),
      .b2_rsci_biwt(b2_rsci_biwt),
      .b2_rsci_bdwt(b2_rsci_bdwt),
      .b2_rsci_bcwt(b2_rsci_bcwt),
      .b2_rsci_idat(b2_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_w2_rsci
// ------------------------------------------------------------------


module econV0_core_w2_rsci (
  clk, rst, w2_rsc_dat, w2_rsc_vld, w2_rsc_rdy, core_wen, w2_rsci_oswt, w2_rsci_wen_comp,
      w2_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [20735:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  input core_wen;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [20735:0] w2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w2_rsci_biwt;
  wire w2_rsci_bdwt;
  wire w2_rsci_bcwt;
  wire w2_rsci_irdy_core_sct;
  wire w2_rsci_ivld;
  wire [20735:0] w2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd26),
  .width(32'sd20736)) w2_rsci (
      .rdy(w2_rsc_rdy),
      .vld(w2_rsc_vld),
      .dat(w2_rsc_dat),
      .irdy(w2_rsci_irdy_core_sct),
      .ivld(w2_rsci_ivld),
      .idat(w2_rsci_idat)
    );
  econV0_core_w2_rsci_w2_rsc_wait_ctrl econV0_core_w2_rsci_w2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .w2_rsci_oswt(w2_rsci_oswt),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_bcwt(w2_rsci_bcwt),
      .w2_rsci_irdy_core_sct(w2_rsci_irdy_core_sct),
      .w2_rsci_ivld(w2_rsci_ivld)
    );
  econV0_core_w2_rsci_w2_rsc_wait_dp econV0_core_w2_rsci_w2_rsc_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .w2_rsci_oswt(w2_rsci_oswt),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_bcwt(w2_rsci_bcwt),
      .w2_rsci_idat(w2_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsci (
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, core_wten, const_size_out_1_rsci_iswt0
);
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input core_wten;
  input const_size_out_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd25),
  .width(32'sd16)) const_size_out_1_rsci (
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000000011),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(const_size_out_1_rsci_iswt0),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsci (
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, core_wten, const_size_in_1_rsci_iswt0
);
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input core_wten;
  input const_size_in_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd24),
  .width(32'sd16)) const_size_in_1_rsci (
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000110000),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(const_size_in_1_rsci_iswt0),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci (
  clk, rst, layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, core_wen,
      layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_idat
);
  input clk;
  input rst;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  input core_wen;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input [53:0] layer7_out_rsci_idat;


  // Interconnect Declarations
  wire layer7_out_rsci_irdy;
  wire layer7_out_rsci_biwt;
  wire layer7_out_rsci_bdwt;
  wire layer7_out_rsci_bcwt;
  wire layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd23),
  .width(32'sd54)) layer7_out_rsci (
      .irdy(layer7_out_rsci_irdy),
      .ivld(layer7_out_rsci_ivld_core_sct),
      .idat(layer7_out_rsci_idat),
      .rdy(layer7_out_rsc_rdy),
      .vld(layer7_out_rsc_vld),
      .dat(layer7_out_rsc_dat)
    );
  econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_irdy(layer7_out_rsci_irdy),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt),
      .layer7_out_rsci_ivld_core_sct(layer7_out_rsci_ivld_core_sct)
    );
  econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci
// ------------------------------------------------------------------


module econV0_core_input_48_rsci (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, core_wen, input_48_rsci_oswt,
      input_48_rsci_wen_comp, input_48_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  input core_wen;
  input input_48_rsci_oswt;
  output input_48_rsci_wen_comp;
  output [863:0] input_48_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_48_rsci_biwt;
  wire input_48_rsci_bdwt;
  wire input_48_rsci_bcwt;
  wire input_48_rsci_irdy_core_sct;
  wire input_48_rsci_ivld;
  wire [863:0] input_48_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd22),
  .width(32'sd864)) input_48_rsci (
      .rdy(input_48_rsc_rdy),
      .vld(input_48_rsc_vld),
      .dat(input_48_rsc_dat),
      .irdy(input_48_rsci_irdy_core_sct),
      .ivld(input_48_rsci_ivld),
      .idat(input_48_rsci_idat)
    );
  econV0_core_input_48_rsci_input_48_rsc_wait_ctrl econV0_core_input_48_rsci_input_48_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .input_48_rsci_oswt(input_48_rsci_oswt),
      .input_48_rsci_biwt(input_48_rsci_biwt),
      .input_48_rsci_bdwt(input_48_rsci_bdwt),
      .input_48_rsci_bcwt(input_48_rsci_bcwt),
      .input_48_rsci_irdy_core_sct(input_48_rsci_irdy_core_sct),
      .input_48_rsci_ivld(input_48_rsci_ivld)
    );
  econV0_core_input_48_rsci_input_48_rsc_wait_dp econV0_core_input_48_rsci_input_48_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_48_rsci_oswt(input_48_rsci_oswt),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .input_48_rsci_idat_mxwt(input_48_rsci_idat_mxwt),
      .input_48_rsci_biwt(input_48_rsci_biwt),
      .input_48_rsci_bdwt(input_48_rsci_bdwt),
      .input_48_rsci_bcwt(input_48_rsci_bcwt),
      .input_48_rsci_idat(input_48_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core
// ------------------------------------------------------------------


module econV0_core (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, input_48_rsc_triosy_lz,
      layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, layer7_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_triosy_lz,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_triosy_lz,
      w2_rsc_dat, w2_rsc_vld, w2_rsc_rdy, w2_rsc_triosy_lz, b2_rsc_dat, b2_rsc_vld,
      b2_rsc_rdy, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, w4_rsc_triosy_lz,
      b4_rsc_dat, b4_rsc_vld, b4_rsc_rdy, b4_rsc_triosy_lz, w6_rsc_dat, w6_rsc_vld,
      w6_rsc_rdy, w6_rsc_triosy_lz, b6_rsc_dat, b6_rsc_vld, b6_rsc_rdy, b6_rsc_triosy_lz
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  output input_48_rsc_triosy_lz;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output layer7_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [20735:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  output w2_rsc_triosy_lz;
  input [431:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  output b2_rsc_triosy_lz;
  input [2591:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  output w4_rsc_triosy_lz;
  input [107:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  output b4_rsc_triosy_lz;
  input [323:0] w6_rsc_dat;
  input w6_rsc_vld;
  output w6_rsc_rdy;
  output w6_rsc_triosy_lz;
  input [53:0] b6_rsc_dat;
  input b6_rsc_vld;
  output b6_rsc_rdy;
  output b6_rsc_triosy_lz;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_48_rsci_wen_comp;
  wire [863:0] input_48_rsci_idat_mxwt;
  wire layer7_out_rsci_wen_comp;
  reg [53:0] layer7_out_rsci_idat;
  wire w2_rsci_wen_comp;
  wire [20735:0] w2_rsci_idat_mxwt;
  wire b2_rsci_wen_comp;
  wire [431:0] b2_rsci_idat_mxwt;
  wire w4_rsci_wen_comp;
  wire [2591:0] w4_rsci_idat_mxwt;
  wire b4_rsci_wen_comp;
  wire [107:0] b4_rsci_idat_mxwt;
  wire w6_rsci_wen_comp;
  wire [323:0] w6_rsci_idat_mxwt;
  wire b6_rsci_wen_comp;
  wire [53:0] b6_rsci_idat_mxwt;
  wire [53:0] nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z;
  wire [53:0] nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z;
  wire [107:0] nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z;
  wire [107:0] nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z;
  wire [431:0] nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z;
  wire [431:0] nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z;
  wire [8:0] fsm_output;
  reg reg_b6_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse;
  wire and_cse;
  reg [323:0] nnet_dense_large_layer5_t_layer6_t_config6_w6_sva;
  reg [53:0] nnet_dense_large_layer5_t_layer6_t_config6_b6_sva;
  reg [2591:0] nnet_dense_large_layer3_t_layer4_t_config4_w4_sva;
  reg [107:0] nnet_dense_large_layer3_t_layer4_t_config4_b4_sva;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[6];
  wire [323:0] nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_weights_rsc_dat;
  assign nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_weights_rsc_dat = nnet_dense_large_layer5_t_layer6_t_config6_w6_sva;
  wire [53:0] nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_biases_rsc_dat;
  assign nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_biases_rsc_dat = nnet_dense_large_layer5_t_layer6_t_config6_b6_sva;
  wire [0:0] nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[5];
  wire [0:0] nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[4];
  wire [2591:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_weights_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_weights_rsc_dat = nnet_dense_large_layer3_t_layer4_t_config4_w4_sva;
  wire [107:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_biases_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_biases_rsc_dat = nnet_dense_large_layer3_t_layer4_t_config4_b4_sva;
  wire [0:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[3];
  wire [0:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[2];
  wire [0:0] nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[1];
  nnet_relu_layer6_t_result_t_relu_config7  nnet_relu_layer6_t_result_t_relu_config7_cmp
      (
      .data_rsc_dat(nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_layer5_t_layer6_t_config6  nnet_dense_large_layer5_t_layer6_t_config6_cmp
      (
      .data_rsc_dat(nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z),
      .res_rsc_z(nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z),
      .weights_rsc_dat(nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_weights_rsc_dat[323:0]),
      .biases_rsc_dat(nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_biases_rsc_dat[53:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_relu_layer4_t_layer5_t_relu_config5  nnet_relu_layer4_t_layer5_t_relu_config5_cmp
      (
      .data_rsc_dat(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_layer3_t_layer4_t_config4  nnet_dense_large_layer3_t_layer4_t_config4_cmp
      (
      .data_rsc_dat(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z),
      .res_rsc_z(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .weights_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_weights_rsc_dat[2591:0]),
      .biases_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_biases_rsc_dat[107:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_relu_layer2_t_layer3_t_relu_config3  nnet_relu_layer2_t_layer3_t_relu_config3_cmp
      (
      .data_rsc_dat(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_input_t_layer2_t_config2  nnet_dense_large_input_t_layer2_t_config2_cmp
      (
      .data_rsc_dat(input_48_rsci_idat_mxwt),
      .res_rsc_z(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .weights_rsc_dat(w2_rsci_idat_mxwt),
      .biases_rsc_dat(b2_rsci_idat_mxwt),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  econV0_core_input_48_rsci econV0_core_input_48_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_48_rsc_dat(input_48_rsc_dat),
      .input_48_rsc_vld(input_48_rsc_vld),
      .input_48_rsc_rdy(input_48_rsc_rdy),
      .core_wen(core_wen),
      .input_48_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .input_48_rsci_idat_mxwt(input_48_rsci_idat_mxwt)
    );
  econV0_core_layer7_out_rsci econV0_core_layer7_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_idat(layer7_out_rsci_idat)
    );
  econV0_core_const_size_in_1_rsci econV0_core_const_size_in_1_rsci_inst (
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_out_1_rsci econV0_core_const_size_out_1_rsci_inst (
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_w2_rsci econV0_core_w2_rsci_inst (
      .clk(clk),
      .rst(rst),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_rdy(w2_rsc_rdy),
      .core_wen(core_wen),
      .w2_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt)
    );
  econV0_core_b2_rsci econV0_core_b2_rsci_inst (
      .clk(clk),
      .rst(rst),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_rdy(b2_rsc_rdy),
      .core_wen(core_wen),
      .b2_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt)
    );
  econV0_core_w4_rsci econV0_core_w4_rsci_inst (
      .clk(clk),
      .rst(rst),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_rdy(w4_rsc_rdy),
      .core_wen(core_wen),
      .w4_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt)
    );
  econV0_core_b4_rsci econV0_core_b4_rsci_inst (
      .clk(clk),
      .rst(rst),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_rdy(b4_rsc_rdy),
      .core_wen(core_wen),
      .b4_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt)
    );
  econV0_core_w6_rsci econV0_core_w6_rsci_inst (
      .clk(clk),
      .rst(rst),
      .w6_rsc_dat(w6_rsc_dat),
      .w6_rsc_vld(w6_rsc_vld),
      .w6_rsc_rdy(w6_rsc_rdy),
      .core_wen(core_wen),
      .w6_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .w6_rsci_wen_comp(w6_rsci_wen_comp),
      .w6_rsci_idat_mxwt(w6_rsci_idat_mxwt)
    );
  econV0_core_b6_rsci econV0_core_b6_rsci_inst (
      .clk(clk),
      .rst(rst),
      .b6_rsc_dat(b6_rsc_dat),
      .b6_rsc_vld(b6_rsc_vld),
      .b6_rsc_rdy(b6_rsc_rdy),
      .core_wen(core_wen),
      .b6_rsci_oswt(reg_b6_rsc_triosy_obj_ld_core_psct_cse),
      .b6_rsci_wen_comp(b6_rsci_wen_comp),
      .b6_rsci_idat_mxwt(b6_rsci_idat_mxwt)
    );
  econV0_core_input_48_rsc_triosy_obj econV0_core_input_48_rsc_triosy_obj_inst (
      .input_48_rsc_triosy_lz(input_48_rsc_triosy_lz),
      .core_wten(core_wten),
      .input_48_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_layer7_out_rsc_triosy_obj econV0_core_layer7_out_rsc_triosy_obj_inst
      (
      .layer7_out_rsc_triosy_lz(layer7_out_rsc_triosy_lz),
      .core_wten(core_wten),
      .layer7_out_rsc_triosy_obj_iswt0(reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_in_1_rsc_triosy_obj econV0_core_const_size_in_1_rsc_triosy_obj_inst
      (
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_out_1_rsc_triosy_obj econV0_core_const_size_out_1_rsc_triosy_obj_inst
      (
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_w2_rsc_triosy_obj econV0_core_w2_rsc_triosy_obj_inst (
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_b2_rsc_triosy_obj econV0_core_b2_rsc_triosy_obj_inst (
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_w4_rsc_triosy_obj econV0_core_w4_rsc_triosy_obj_inst (
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_b4_rsc_triosy_obj econV0_core_b4_rsc_triosy_obj_inst (
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz),
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_w6_rsc_triosy_obj econV0_core_w6_rsc_triosy_obj_inst (
      .w6_rsc_triosy_lz(w6_rsc_triosy_lz),
      .core_wten(core_wten),
      .w6_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_b6_rsc_triosy_obj econV0_core_b6_rsc_triosy_obj_inst (
      .b6_rsc_triosy_lz(b6_rsc_triosy_lz),
      .core_wten(core_wten),
      .b6_rsc_triosy_obj_iswt0(reg_b6_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_staller econV0_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .w6_rsci_wen_comp(w6_rsci_wen_comp),
      .b6_rsci_wen_comp(b6_rsci_wen_comp)
    );
  econV0_core_core_fsm econV0_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_cse = core_wen & (fsm_output[1]);
  always @(posedge clk) begin
    if ( rst ) begin
      reg_b6_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_b6_rsc_triosy_obj_ld_core_psct_cse <= (fsm_output[8]) | (fsm_output[0]);
      reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse <= fsm_output[7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat <= 54'b000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (fsm_output[7]) ) begin
      layer7_out_rsci_idat <= nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_dense_large_layer5_t_layer6_t_config6_b6_sva <= 54'b000000000000000000000000000000000000000000000000000000;
      nnet_dense_large_layer5_t_layer6_t_config6_w6_sva <= 324'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nnet_dense_large_layer3_t_layer4_t_config4_b4_sva <= 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nnet_dense_large_layer3_t_layer4_t_config4_w4_sva <= {648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( and_cse ) begin
      nnet_dense_large_layer5_t_layer6_t_config6_b6_sva <= b6_rsci_idat_mxwt;
      nnet_dense_large_layer5_t_layer6_t_config6_w6_sva <= w6_rsci_idat_mxwt;
      nnet_dense_large_layer3_t_layer4_t_config4_b4_sva <= b4_rsci_idat_mxwt;
      nnet_dense_large_layer3_t_layer4_t_config4_w4_sva <= w4_rsci_idat_mxwt;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0
// ------------------------------------------------------------------


module econV0 (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, input_48_rsc_triosy_lz,
      layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, layer7_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_triosy_lz,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_triosy_lz,
      w2_rsc_dat, w2_rsc_vld, w2_rsc_rdy, w2_rsc_triosy_lz, b2_rsc_dat, b2_rsc_vld,
      b2_rsc_rdy, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, w4_rsc_triosy_lz,
      b4_rsc_dat, b4_rsc_vld, b4_rsc_rdy, b4_rsc_triosy_lz, w6_rsc_dat, w6_rsc_vld,
      w6_rsc_rdy, w6_rsc_triosy_lz, b6_rsc_dat, b6_rsc_vld, b6_rsc_rdy, b6_rsc_triosy_lz
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  output input_48_rsc_triosy_lz;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output layer7_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [20735:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  output w2_rsc_triosy_lz;
  input [431:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  output b2_rsc_triosy_lz;
  input [2591:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  output w4_rsc_triosy_lz;
  input [107:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  output b4_rsc_triosy_lz;
  input [323:0] w6_rsc_dat;
  input w6_rsc_vld;
  output w6_rsc_rdy;
  output w6_rsc_triosy_lz;
  input [53:0] b6_rsc_dat;
  input b6_rsc_vld;
  output b6_rsc_rdy;
  output b6_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  econV0_core econV0_core_inst (
      .clk(clk),
      .rst(rst),
      .input_48_rsc_dat(input_48_rsc_dat),
      .input_48_rsc_vld(input_48_rsc_vld),
      .input_48_rsc_rdy(input_48_rsc_rdy),
      .input_48_rsc_triosy_lz(input_48_rsc_triosy_lz),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .layer7_out_rsc_triosy_lz(layer7_out_rsc_triosy_lz),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_rdy(w2_rsc_rdy),
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_rdy(b2_rsc_rdy),
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_rdy(w4_rsc_rdy),
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_rdy(b4_rsc_rdy),
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz),
      .w6_rsc_dat(w6_rsc_dat),
      .w6_rsc_vld(w6_rsc_vld),
      .w6_rsc_rdy(w6_rsc_rdy),
      .w6_rsc_triosy_lz(w6_rsc_triosy_lz),
      .b6_rsc_dat(b6_rsc_dat),
      .b6_rsc_vld(b6_rsc_vld),
      .b6_rsc_rdy(b6_rsc_rdy),
      .b6_rsc_triosy_lz(b6_rsc_triosy_lz)
    );
endmodule



