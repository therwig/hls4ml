
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5/861329 Production Release
//  HLS Date:       Wed Mar  4 15:45:36 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Mar 13 15:33:17 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module econ_4x4_d10_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for econ_4x4_d10_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : econ_4x4_d10_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_staller
// ------------------------------------------------------------------


module econ_4x4_d10_core_staller (
  clk, rst, core_wen, core_wten, input_1_rsci_wen_comp, layer5_out_rsci_wen_comp,
      const_size_in_1_rsci_wen_comp, const_size_out_1_rsci_wen_comp, w2_rsci_wen_comp,
      b2_rsci_wen_comp, w4_rsci_wen_comp, b4_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_1_rsci_wen_comp;
  input layer5_out_rsci_wen_comp;
  input const_size_in_1_rsci_wen_comp;
  input const_size_out_1_rsci_wen_comp;
  input w2_rsci_wen_comp;
  input b2_rsci_wen_comp;
  input w4_rsci_wen_comp;
  input b4_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_1_rsci_wen_comp & layer5_out_rsci_wen_comp & const_size_in_1_rsci_wen_comp
      & const_size_out_1_rsci_wen_comp & w2_rsci_wen_comp & b2_rsci_wen_comp & w4_rsci_wen_comp
      & b4_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl (
  core_wten, b4_rsc_triosy_obj_iswt0, b4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;
  output b4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b4_rsc_triosy_obj_ld_core_sct = b4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl (
  core_wten, w4_rsc_triosy_obj_iswt0, w4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;
  output w4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w4_rsc_triosy_obj_ld_core_sct = w4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl (
  core_wten, b2_rsc_triosy_obj_iswt0, b2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;
  output b2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b2_rsc_triosy_obj_ld_core_sct = b2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl (
  core_wten, w2_rsc_triosy_obj_iswt0, w2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;
  output w2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w2_rsc_triosy_obj_ld_core_sct = w2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_out_1_rsc_triosy_obj_iswt0, const_size_out_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;
  output const_size_out_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsc_triosy_obj_ld_core_sct = const_size_out_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_in_1_rsc_triosy_obj_iswt0, const_size_in_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;
  output const_size_in_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsc_triosy_obj_ld_core_sct = const_size_in_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
    (
  core_wten, layer5_out_rsc_triosy_obj_iswt0, layer5_out_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;
  output layer5_out_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsc_triosy_obj_ld_core_sct = layer5_out_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl (
  core_wten, input_1_rsc_triosy_obj_iswt0, input_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;
  output input_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsc_triosy_obj_ld_core_sct = input_1_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsci_b4_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsci_b4_rsc_wait_dp (
  clk, rst, b4_rsci_oswt, b4_rsci_wen_comp, b4_rsci_idat_mxwt, b4_rsci_biwt, b4_rsci_bdwt,
      b4_rsci_bcwt, b4_rsci_idat
);
  input clk;
  input rst;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [69:0] b4_rsci_idat_mxwt;
  input b4_rsci_biwt;
  input b4_rsci_bdwt;
  output b4_rsci_bcwt;
  reg b4_rsci_bcwt;
  input [79:0] b4_rsci_idat;


  // Interconnect Declarations
  wire [78:0] b4_rsci_idat_mxwt_pconst;
  reg [78:0] b4_rsci_idat_bfwt_79_1;


  // Interconnect Declarations for Component Instantiations 
  assign b4_rsci_wen_comp = (~ b4_rsci_oswt) | b4_rsci_biwt | b4_rsci_bcwt;
  assign b4_rsci_idat_mxwt_pconst = MUX_v_79_2_2((b4_rsci_idat[79:1]), b4_rsci_idat_bfwt_79_1,
      b4_rsci_bcwt);
  assign b4_rsci_idat_mxwt = {(b4_rsci_idat_mxwt_pconst[78:72]) , (b4_rsci_idat_mxwt_pconst[70:64])
      , (b4_rsci_idat_mxwt_pconst[62:56]) , (b4_rsci_idat_mxwt_pconst[54:48]) , (b4_rsci_idat_mxwt_pconst[46:40])
      , (b4_rsci_idat_mxwt_pconst[38:32]) , (b4_rsci_idat_mxwt_pconst[30:24]) , (b4_rsci_idat_mxwt_pconst[22:16])
      , (b4_rsci_idat_mxwt_pconst[14:8]) , (b4_rsci_idat_mxwt_pconst[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      b4_rsci_bcwt <= 1'b0;
    end
    else begin
      b4_rsci_bcwt <= ~((~(b4_rsci_bcwt | b4_rsci_biwt)) | b4_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      b4_rsci_idat_bfwt_79_1 <= 79'b0000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( b4_rsci_biwt ) begin
      b4_rsci_idat_bfwt_79_1 <= b4_rsci_idat[79:1];
    end
  end

  function automatic [78:0] MUX_v_79_2_2;
    input [78:0] input_0;
    input [78:0] input_1;
    input [0:0] sel;
    reg [78:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_79_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsci_b4_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsci_b4_rsc_wait_ctrl (
  core_wen, b4_rsci_oswt, b4_rsci_biwt, b4_rsci_bdwt, b4_rsci_bcwt, b4_rsci_irdy_core_sct,
      b4_rsci_ivld
);
  input core_wen;
  input b4_rsci_oswt;
  output b4_rsci_biwt;
  output b4_rsci_bdwt;
  input b4_rsci_bcwt;
  output b4_rsci_irdy_core_sct;
  input b4_rsci_ivld;


  // Interconnect Declarations
  wire b4_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b4_rsci_bdwt = b4_rsci_oswt & core_wen;
  assign b4_rsci_biwt = b4_rsci_ogwt & b4_rsci_ivld;
  assign b4_rsci_ogwt = b4_rsci_oswt & (~ b4_rsci_bcwt);
  assign b4_rsci_irdy_core_sct = b4_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsci_w4_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsci_w4_rsc_wait_dp (
  clk, rst, w4_rsci_oswt, w4_rsci_wen_comp, w4_rsci_idat_mxwt, w4_rsci_biwt, w4_rsci_bdwt,
      w4_rsci_bcwt, w4_rsci_idat
);
  input clk;
  input rst;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [10239:0] w4_rsci_idat_mxwt;
  input w4_rsci_biwt;
  input w4_rsci_bdwt;
  output w4_rsci_bcwt;
  reg w4_rsci_bcwt;
  input [10239:0] w4_rsci_idat;


  // Interconnect Declarations
  reg [10239:0] w4_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w4_rsci_wen_comp = (~ w4_rsci_oswt) | w4_rsci_biwt | w4_rsci_bcwt;
  assign w4_rsci_idat_mxwt = MUX_v_10240_2_2(w4_rsci_idat, w4_rsci_idat_bfwt, w4_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_bcwt <= 1'b0;
    end
    else begin
      w4_rsci_bcwt <= ~((~(w4_rsci_bcwt | w4_rsci_biwt)) | w4_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w4_rsci_idat_bfwt <= {640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( w4_rsci_biwt ) begin
      w4_rsci_idat_bfwt <= w4_rsci_idat;
    end
  end

  function automatic [10239:0] MUX_v_10240_2_2;
    input [10239:0] input_0;
    input [10239:0] input_1;
    input [0:0] sel;
    reg [10239:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10240_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsci_w4_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsci_w4_rsc_wait_ctrl (
  core_wen, w4_rsci_oswt, w4_rsci_biwt, w4_rsci_bdwt, w4_rsci_bcwt, w4_rsci_irdy_core_sct,
      w4_rsci_ivld
);
  input core_wen;
  input w4_rsci_oswt;
  output w4_rsci_biwt;
  output w4_rsci_bdwt;
  input w4_rsci_bcwt;
  output w4_rsci_irdy_core_sct;
  input w4_rsci_ivld;


  // Interconnect Declarations
  wire w4_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w4_rsci_bdwt = w4_rsci_oswt & core_wen;
  assign w4_rsci_biwt = w4_rsci_ogwt & w4_rsci_ivld;
  assign w4_rsci_ogwt = w4_rsci_oswt & (~ w4_rsci_bcwt);
  assign w4_rsci_irdy_core_sct = w4_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsci_b2_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsci_b2_rsc_wait_dp (
  clk, rst, b2_rsci_oswt, b2_rsci_wen_comp, b2_rsci_idat_mxwt, b2_rsci_biwt, b2_rsci_bdwt,
      b2_rsci_bcwt, b2_rsci_idat
);
  input clk;
  input rst;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [55:0] b2_rsci_idat_mxwt;
  input b2_rsci_biwt;
  input b2_rsci_bdwt;
  output b2_rsci_bcwt;
  reg b2_rsci_bcwt;
  input [63:0] b2_rsci_idat;


  // Interconnect Declarations
  wire [62:0] b2_rsci_idat_mxwt_pconst;
  reg [62:0] b2_rsci_idat_bfwt_63_1;


  // Interconnect Declarations for Component Instantiations 
  assign b2_rsci_wen_comp = (~ b2_rsci_oswt) | b2_rsci_biwt | b2_rsci_bcwt;
  assign b2_rsci_idat_mxwt_pconst = MUX_v_63_2_2((b2_rsci_idat[63:1]), b2_rsci_idat_bfwt_63_1,
      b2_rsci_bcwt);
  assign b2_rsci_idat_mxwt = {(b2_rsci_idat_mxwt_pconst[62:56]) , (b2_rsci_idat_mxwt_pconst[54:48])
      , (b2_rsci_idat_mxwt_pconst[46:40]) , (b2_rsci_idat_mxwt_pconst[38:32]) , (b2_rsci_idat_mxwt_pconst[30:24])
      , (b2_rsci_idat_mxwt_pconst[22:16]) , (b2_rsci_idat_mxwt_pconst[14:8]) , (b2_rsci_idat_mxwt_pconst[6:0])};
  always @(posedge clk) begin
    if ( rst ) begin
      b2_rsci_bcwt <= 1'b0;
    end
    else begin
      b2_rsci_bcwt <= ~((~(b2_rsci_bcwt | b2_rsci_biwt)) | b2_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      b2_rsci_idat_bfwt_63_1 <= 63'b000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( b2_rsci_biwt ) begin
      b2_rsci_idat_bfwt_63_1 <= b2_rsci_idat[63:1];
    end
  end

  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsci_b2_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsci_b2_rsc_wait_ctrl (
  core_wen, b2_rsci_oswt, b2_rsci_biwt, b2_rsci_bdwt, b2_rsci_bcwt, b2_rsci_irdy_core_sct,
      b2_rsci_ivld
);
  input core_wen;
  input b2_rsci_oswt;
  output b2_rsci_biwt;
  output b2_rsci_bdwt;
  input b2_rsci_bcwt;
  output b2_rsci_irdy_core_sct;
  input b2_rsci_ivld;


  // Interconnect Declarations
  wire b2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b2_rsci_bdwt = b2_rsci_oswt & core_wen;
  assign b2_rsci_biwt = b2_rsci_ogwt & b2_rsci_ivld;
  assign b2_rsci_ogwt = b2_rsci_oswt & (~ b2_rsci_bcwt);
  assign b2_rsci_irdy_core_sct = b2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsci_w2_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsci_w2_rsc_wait_dp (
  clk, rst, w2_rsci_oswt, w2_rsci_wen_comp, w2_rsci_idat_mxwt, w2_rsci_biwt, w2_rsci_bdwt,
      w2_rsci_bcwt, w2_rsci_idat
);
  input clk;
  input rst;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [1727:0] w2_rsci_idat_mxwt;
  input w2_rsci_biwt;
  input w2_rsci_bdwt;
  output w2_rsci_bcwt;
  reg w2_rsci_bcwt;
  input [1727:0] w2_rsci_idat;


  // Interconnect Declarations
  reg [1727:0] w2_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign w2_rsci_wen_comp = (~ w2_rsci_oswt) | w2_rsci_biwt | w2_rsci_bcwt;
  assign w2_rsci_idat_mxwt = MUX_v_1728_2_2(w2_rsci_idat, w2_rsci_idat_bfwt, w2_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_bcwt <= 1'b0;
    end
    else begin
      w2_rsci_bcwt <= ~((~(w2_rsci_bcwt | w2_rsci_biwt)) | w2_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      w2_rsci_idat_bfwt <= {864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
    end
    else if ( w2_rsci_biwt ) begin
      w2_rsci_idat_bfwt <= w2_rsci_idat;
    end
  end

  function automatic [1727:0] MUX_v_1728_2_2;
    input [1727:0] input_0;
    input [1727:0] input_1;
    input [0:0] sel;
    reg [1727:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1728_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsci_w2_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsci_w2_rsc_wait_ctrl (
  core_wen, w2_rsci_oswt, w2_rsci_biwt, w2_rsci_bdwt, w2_rsci_bcwt, w2_rsci_irdy_core_sct,
      w2_rsci_ivld
);
  input core_wen;
  input w2_rsci_oswt;
  output w2_rsci_biwt;
  output w2_rsci_bdwt;
  input w2_rsci_bcwt;
  output w2_rsci_irdy_core_sct;
  input w2_rsci_ivld;


  // Interconnect Declarations
  wire w2_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign w2_rsci_bdwt = w2_rsci_oswt & core_wen;
  assign w2_rsci_biwt = w2_rsci_ogwt & w2_rsci_ivld;
  assign w2_rsci_ogwt = w2_rsci_oswt & (~ w2_rsci_bcwt);
  assign w2_rsci_irdy_core_sct = w2_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp (
  clk, rst, const_size_out_1_rsci_oswt, const_size_out_1_rsci_wen_comp, const_size_out_1_rsci_biwt,
      const_size_out_1_rsci_bdwt, const_size_out_1_rsci_bcwt
);
  input clk;
  input rst;
  input const_size_out_1_rsci_oswt;
  output const_size_out_1_rsci_wen_comp;
  input const_size_out_1_rsci_biwt;
  input const_size_out_1_rsci_bdwt;
  output const_size_out_1_rsci_bcwt;
  reg const_size_out_1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_wen_comp = (~ const_size_out_1_rsci_oswt) | const_size_out_1_rsci_biwt
      | const_size_out_1_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      const_size_out_1_rsci_bcwt <= 1'b0;
    end
    else begin
      const_size_out_1_rsci_bcwt <= ~((~(const_size_out_1_rsci_bcwt | const_size_out_1_rsci_biwt))
          | const_size_out_1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wen, const_size_out_1_rsci_oswt, const_size_out_1_rsci_irdy, const_size_out_1_rsci_biwt,
      const_size_out_1_rsci_bdwt, const_size_out_1_rsci_bcwt, const_size_out_1_rsci_ivld_core_sct
);
  input core_wen;
  input const_size_out_1_rsci_oswt;
  input const_size_out_1_rsci_irdy;
  output const_size_out_1_rsci_biwt;
  output const_size_out_1_rsci_bdwt;
  input const_size_out_1_rsci_bcwt;
  output const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_bdwt = const_size_out_1_rsci_oswt & core_wen;
  assign const_size_out_1_rsci_biwt = const_size_out_1_rsci_ogwt & const_size_out_1_rsci_irdy;
  assign const_size_out_1_rsci_ogwt = const_size_out_1_rsci_oswt & (~ const_size_out_1_rsci_bcwt);
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp (
  clk, rst, const_size_in_1_rsci_oswt, const_size_in_1_rsci_wen_comp, const_size_in_1_rsci_biwt,
      const_size_in_1_rsci_bdwt, const_size_in_1_rsci_bcwt
);
  input clk;
  input rst;
  input const_size_in_1_rsci_oswt;
  output const_size_in_1_rsci_wen_comp;
  input const_size_in_1_rsci_biwt;
  input const_size_in_1_rsci_bdwt;
  output const_size_in_1_rsci_bcwt;
  reg const_size_in_1_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_wen_comp = (~ const_size_in_1_rsci_oswt) | const_size_in_1_rsci_biwt
      | const_size_in_1_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      const_size_in_1_rsci_bcwt <= 1'b0;
    end
    else begin
      const_size_in_1_rsci_bcwt <= ~((~(const_size_in_1_rsci_bcwt | const_size_in_1_rsci_biwt))
          | const_size_in_1_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wen, const_size_in_1_rsci_oswt, const_size_in_1_rsci_irdy, const_size_in_1_rsci_biwt,
      const_size_in_1_rsci_bdwt, const_size_in_1_rsci_bcwt, const_size_in_1_rsci_ivld_core_sct
);
  input core_wen;
  input const_size_in_1_rsci_oswt;
  input const_size_in_1_rsci_irdy;
  output const_size_in_1_rsci_biwt;
  output const_size_in_1_rsci_bdwt;
  input const_size_in_1_rsci_bcwt;
  output const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_bdwt = const_size_in_1_rsci_oswt & core_wen;
  assign const_size_in_1_rsci_biwt = const_size_in_1_rsci_ogwt & const_size_in_1_rsci_irdy;
  assign const_size_in_1_rsci_ogwt = const_size_in_1_rsci_oswt & (~ const_size_in_1_rsci_bcwt);
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_dp (
  clk, rst, layer5_out_rsci_oswt, layer5_out_rsci_wen_comp, layer5_out_rsci_biwt,
      layer5_out_rsci_bdwt, layer5_out_rsci_bcwt
);
  input clk;
  input rst;
  input layer5_out_rsci_oswt;
  output layer5_out_rsci_wen_comp;
  input layer5_out_rsci_biwt;
  input layer5_out_rsci_bdwt;
  output layer5_out_rsci_bcwt;
  reg layer5_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_wen_comp = (~ layer5_out_rsci_oswt) | layer5_out_rsci_biwt
      | layer5_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_bcwt <= 1'b0;
    end
    else begin
      layer5_out_rsci_bcwt <= ~((~(layer5_out_rsci_bcwt | layer5_out_rsci_biwt))
          | layer5_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl (
  core_wen, layer5_out_rsci_oswt, layer5_out_rsci_irdy, layer5_out_rsci_biwt, layer5_out_rsci_bdwt,
      layer5_out_rsci_bcwt, layer5_out_rsci_ivld_core_sct
);
  input core_wen;
  input layer5_out_rsci_oswt;
  input layer5_out_rsci_irdy;
  output layer5_out_rsci_biwt;
  output layer5_out_rsci_bdwt;
  input layer5_out_rsci_bcwt;
  output layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire layer5_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_bdwt = layer5_out_rsci_oswt & core_wen;
  assign layer5_out_rsci_biwt = layer5_out_rsci_ogwt & layer5_out_rsci_irdy;
  assign layer5_out_rsci_ogwt = layer5_out_rsci_oswt & (~ layer5_out_rsci_bcwt);
  assign layer5_out_rsci_ivld_core_sct = layer5_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_dp
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_dp (
  clk, rst, input_1_rsci_oswt, input_1_rsci_wen_comp, input_1_rsci_idat_mxwt, input_1_rsci_biwt,
      input_1_rsci_bdwt, input_1_rsci_bcwt, input_1_rsci_idat
);
  input clk;
  input rst;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [383:0] input_1_rsci_idat_mxwt;
  input input_1_rsci_biwt;
  input input_1_rsci_bdwt;
  output input_1_rsci_bcwt;
  reg input_1_rsci_bcwt;
  input [383:0] input_1_rsci_idat;


  // Interconnect Declarations
  reg [383:0] input_1_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsci_wen_comp = (~ input_1_rsci_oswt) | input_1_rsci_biwt | input_1_rsci_bcwt;
  assign input_1_rsci_idat_mxwt = MUX_v_384_2_2(input_1_rsci_idat, input_1_rsci_idat_bfwt,
      input_1_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input_1_rsci_bcwt <= 1'b0;
    end
    else begin
      input_1_rsci_bcwt <= ~((~(input_1_rsci_bcwt | input_1_rsci_biwt)) | input_1_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_1_rsci_idat_bfwt <= 384'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( input_1_rsci_biwt ) begin
      input_1_rsci_idat_bfwt <= input_1_rsci_idat;
    end
  end

  function automatic [383:0] MUX_v_384_2_2;
    input [383:0] input_0;
    input [383:0] input_1;
    input [0:0] sel;
    reg [383:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_384_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_ctrl (
  core_wen, input_1_rsci_oswt, input_1_rsci_biwt, input_1_rsci_bdwt, input_1_rsci_bcwt,
      input_1_rsci_irdy_core_sct, input_1_rsci_ivld
);
  input core_wen;
  input input_1_rsci_oswt;
  output input_1_rsci_biwt;
  output input_1_rsci_bdwt;
  input input_1_rsci_bcwt;
  output input_1_rsci_irdy_core_sct;
  input input_1_rsci_ivld;


  // Interconnect Declarations
  wire input_1_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsci_bdwt = input_1_rsci_oswt & core_wen;
  assign input_1_rsci_biwt = input_1_rsci_ogwt & input_1_rsci_ivld;
  assign input_1_rsci_ogwt = input_1_rsci_oswt & (~ input_1_rsci_bcwt);
  assign input_1_rsci_irdy_core_sct = input_1_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj (
  b4_rsc_triosy_lz, core_wten, b4_rsc_triosy_obj_iswt0
);
  output b4_rsc_triosy_lz;
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b4_rsc_triosy_obj (
      .ld(b4_rsc_triosy_obj_ld_core_sct),
      .lz(b4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(b4_rsc_triosy_obj_iswt0),
      .b4_rsc_triosy_obj_ld_core_sct(b4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj (
  w4_rsc_triosy_lz, core_wten, w4_rsc_triosy_obj_iswt0
);
  output w4_rsc_triosy_lz;
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w4_rsc_triosy_obj (
      .ld(w4_rsc_triosy_obj_ld_core_sct),
      .lz(w4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(w4_rsc_triosy_obj_iswt0),
      .w4_rsc_triosy_obj_ld_core_sct(w4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj (
  b2_rsc_triosy_lz, core_wten, b2_rsc_triosy_obj_iswt0
);
  output b2_rsc_triosy_lz;
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b2_rsc_triosy_obj (
      .ld(b2_rsc_triosy_obj_ld_core_sct),
      .lz(b2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(b2_rsc_triosy_obj_iswt0),
      .b2_rsc_triosy_obj_ld_core_sct(b2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj (
  w2_rsc_triosy_lz, core_wten, w2_rsc_triosy_obj_iswt0
);
  output w2_rsc_triosy_lz;
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w2_rsc_triosy_obj (
      .ld(w2_rsc_triosy_obj_ld_core_sct),
      .lz(w2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(w2_rsc_triosy_obj_iswt0),
      .w2_rsc_triosy_obj_ld_core_sct(w2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj (
  const_size_out_1_rsc_triosy_lz, core_wten, const_size_out_1_rsc_triosy_obj_iswt0
);
  output const_size_out_1_rsc_triosy_lz;
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_out_1_rsc_triosy_obj (
      .ld(const_size_out_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_out_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(const_size_out_1_rsc_triosy_obj_iswt0),
      .const_size_out_1_rsc_triosy_obj_ld_core_sct(const_size_out_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj (
  const_size_in_1_rsc_triosy_lz, core_wten, const_size_in_1_rsc_triosy_obj_iswt0
);
  output const_size_in_1_rsc_triosy_lz;
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_in_1_rsc_triosy_obj (
      .ld(const_size_in_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_in_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(const_size_in_1_rsc_triosy_obj_iswt0),
      .const_size_in_1_rsc_triosy_obj_ld_core_sct(const_size_in_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj (
  layer5_out_rsc_triosy_lz, core_wten, layer5_out_rsc_triosy_obj_iswt0
);
  output layer5_out_rsc_triosy_lz;
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire layer5_out_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) layer5_out_rsc_triosy_obj (
      .ld(layer5_out_rsc_triosy_obj_ld_core_sct),
      .lz(layer5_out_rsc_triosy_lz)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(layer5_out_rsc_triosy_obj_iswt0),
      .layer5_out_rsc_triosy_obj_ld_core_sct(layer5_out_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj (
  input_1_rsc_triosy_lz, core_wten, input_1_rsc_triosy_obj_iswt0
);
  output input_1_rsc_triosy_lz;
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire input_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) input_1_rsc_triosy_obj (
      .ld(input_1_rsc_triosy_obj_ld_core_sct),
      .lz(input_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(input_1_rsc_triosy_obj_iswt0),
      .input_1_rsc_triosy_obj_ld_core_sct(input_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsci (
  clk, rst, b4_rsc_dat, b4_rsc_vld, b4_rsc_rdy, core_wen, b4_rsci_oswt, b4_rsci_wen_comp,
      b4_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  input core_wen;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [69:0] b4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b4_rsci_biwt;
  wire b4_rsci_bdwt;
  wire b4_rsci_bcwt;
  wire b4_rsci_irdy_core_sct;
  wire b4_rsci_ivld;
  wire [79:0] b4_rsci_idat;
  wire [69:0] b4_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd8),
  .width(32'sd80)) b4_rsci (
      .rdy(b4_rsc_rdy),
      .vld(b4_rsc_vld),
      .dat(b4_rsc_dat),
      .irdy(b4_rsci_irdy_core_sct),
      .ivld(b4_rsci_ivld),
      .idat(b4_rsci_idat)
    );
  econ_4x4_d10_core_b4_rsci_b4_rsc_wait_ctrl econ_4x4_d10_core_b4_rsci_b4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .b4_rsci_oswt(b4_rsci_oswt),
      .b4_rsci_biwt(b4_rsci_biwt),
      .b4_rsci_bdwt(b4_rsci_bdwt),
      .b4_rsci_bcwt(b4_rsci_bcwt),
      .b4_rsci_irdy_core_sct(b4_rsci_irdy_core_sct),
      .b4_rsci_ivld(b4_rsci_ivld)
    );
  econ_4x4_d10_core_b4_rsci_b4_rsc_wait_dp econ_4x4_d10_core_b4_rsci_b4_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .b4_rsci_oswt(b4_rsci_oswt),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt_pconst),
      .b4_rsci_biwt(b4_rsci_biwt),
      .b4_rsci_bdwt(b4_rsci_bdwt),
      .b4_rsci_bcwt(b4_rsci_bcwt),
      .b4_rsci_idat(b4_rsci_idat)
    );
  assign b4_rsci_idat_mxwt = b4_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsci (
  clk, rst, w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, core_wen, w4_rsci_oswt, w4_rsci_wen_comp,
      w4_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  input core_wen;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [10239:0] w4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w4_rsci_biwt;
  wire w4_rsci_bdwt;
  wire w4_rsci_bcwt;
  wire w4_rsci_irdy_core_sct;
  wire w4_rsci_ivld;
  wire [10239:0] w4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd10240)) w4_rsci (
      .rdy(w4_rsc_rdy),
      .vld(w4_rsc_vld),
      .dat(w4_rsc_dat),
      .irdy(w4_rsci_irdy_core_sct),
      .ivld(w4_rsci_ivld),
      .idat(w4_rsci_idat)
    );
  econ_4x4_d10_core_w4_rsci_w4_rsc_wait_ctrl econ_4x4_d10_core_w4_rsci_w4_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .w4_rsci_oswt(w4_rsci_oswt),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_bcwt(w4_rsci_bcwt),
      .w4_rsci_irdy_core_sct(w4_rsci_irdy_core_sct),
      .w4_rsci_ivld(w4_rsci_ivld)
    );
  econ_4x4_d10_core_w4_rsci_w4_rsc_wait_dp econ_4x4_d10_core_w4_rsci_w4_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .w4_rsci_oswt(w4_rsci_oswt),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt),
      .w4_rsci_biwt(w4_rsci_biwt),
      .w4_rsci_bdwt(w4_rsci_bdwt),
      .w4_rsci_bcwt(w4_rsci_bcwt),
      .w4_rsci_idat(w4_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsci (
  clk, rst, b2_rsc_dat, b2_rsc_vld, b2_rsc_rdy, core_wen, b2_rsci_oswt, b2_rsci_wen_comp,
      b2_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  input core_wen;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [55:0] b2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b2_rsci_biwt;
  wire b2_rsci_bdwt;
  wire b2_rsci_bcwt;
  wire b2_rsci_irdy_core_sct;
  wire b2_rsci_ivld;
  wire [63:0] b2_rsci_idat;
  wire [55:0] b2_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd64)) b2_rsci (
      .rdy(b2_rsc_rdy),
      .vld(b2_rsc_vld),
      .dat(b2_rsc_dat),
      .irdy(b2_rsci_irdy_core_sct),
      .ivld(b2_rsci_ivld),
      .idat(b2_rsci_idat)
    );
  econ_4x4_d10_core_b2_rsci_b2_rsc_wait_ctrl econ_4x4_d10_core_b2_rsci_b2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .b2_rsci_oswt(b2_rsci_oswt),
      .b2_rsci_biwt(b2_rsci_biwt),
      .b2_rsci_bdwt(b2_rsci_bdwt),
      .b2_rsci_bcwt(b2_rsci_bcwt),
      .b2_rsci_irdy_core_sct(b2_rsci_irdy_core_sct),
      .b2_rsci_ivld(b2_rsci_ivld)
    );
  econ_4x4_d10_core_b2_rsci_b2_rsc_wait_dp econ_4x4_d10_core_b2_rsci_b2_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .b2_rsci_oswt(b2_rsci_oswt),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt_pconst),
      .b2_rsci_biwt(b2_rsci_biwt),
      .b2_rsci_bdwt(b2_rsci_bdwt),
      .b2_rsci_bcwt(b2_rsci_bcwt),
      .b2_rsci_idat(b2_rsci_idat)
    );
  assign b2_rsci_idat_mxwt = b2_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsci (
  clk, rst, w2_rsc_dat, w2_rsc_vld, w2_rsc_rdy, core_wen, w2_rsci_oswt, w2_rsci_wen_comp,
      w2_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  input core_wen;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [1727:0] w2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w2_rsci_biwt;
  wire w2_rsci_bdwt;
  wire w2_rsci_bcwt;
  wire w2_rsci_irdy_core_sct;
  wire w2_rsci_ivld;
  wire [1727:0] w2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd1728)) w2_rsci (
      .rdy(w2_rsc_rdy),
      .vld(w2_rsc_vld),
      .dat(w2_rsc_dat),
      .irdy(w2_rsci_irdy_core_sct),
      .ivld(w2_rsci_ivld),
      .idat(w2_rsci_idat)
    );
  econ_4x4_d10_core_w2_rsci_w2_rsc_wait_ctrl econ_4x4_d10_core_w2_rsci_w2_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .w2_rsci_oswt(w2_rsci_oswt),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_bcwt(w2_rsci_bcwt),
      .w2_rsci_irdy_core_sct(w2_rsci_irdy_core_sct),
      .w2_rsci_ivld(w2_rsci_ivld)
    );
  econ_4x4_d10_core_w2_rsci_w2_rsc_wait_dp econ_4x4_d10_core_w2_rsci_w2_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .w2_rsci_oswt(w2_rsci_oswt),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt),
      .w2_rsci_biwt(w2_rsci_biwt),
      .w2_rsci_bdwt(w2_rsci_bdwt),
      .w2_rsci_bcwt(w2_rsci_bcwt),
      .w2_rsci_idat(w2_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci (
  clk, rst, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_rdy,
      core_wen, const_size_out_1_rsci_oswt, const_size_out_1_rsci_wen_comp
);
  input clk;
  input rst;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  input core_wen;
  input const_size_out_1_rsci_oswt;
  output const_size_out_1_rsci_wen_comp;


  // Interconnect Declarations
  wire const_size_out_1_rsci_irdy;
  wire const_size_out_1_rsci_biwt;
  wire const_size_out_1_rsci_bdwt;
  wire const_size_out_1_rsci_bcwt;
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd16)) const_size_out_1_rsci (
      .irdy(const_size_out_1_rsci_irdy),
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000001010),
      .rdy(const_size_out_1_rsc_rdy),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .const_size_out_1_rsci_oswt(const_size_out_1_rsci_oswt),
      .const_size_out_1_rsci_irdy(const_size_out_1_rsci_irdy),
      .const_size_out_1_rsci_biwt(const_size_out_1_rsci_biwt),
      .const_size_out_1_rsci_bdwt(const_size_out_1_rsci_bdwt),
      .const_size_out_1_rsci_bcwt(const_size_out_1_rsci_bcwt),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
  econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_out_1_rsci_oswt(const_size_out_1_rsci_oswt),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp),
      .const_size_out_1_rsci_biwt(const_size_out_1_rsci_biwt),
      .const_size_out_1_rsci_bdwt(const_size_out_1_rsci_bdwt),
      .const_size_out_1_rsci_bcwt(const_size_out_1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci (
  clk, rst, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
      core_wen, const_size_in_1_rsci_oswt, const_size_in_1_rsci_wen_comp
);
  input clk;
  input rst;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  input core_wen;
  input const_size_in_1_rsci_oswt;
  output const_size_in_1_rsci_wen_comp;


  // Interconnect Declarations
  wire const_size_in_1_rsci_irdy;
  wire const_size_in_1_rsci_biwt;
  wire const_size_in_1_rsci_bdwt;
  wire const_size_in_1_rsci_bcwt;
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd16)) const_size_in_1_rsci (
      .irdy(const_size_in_1_rsci_irdy),
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000110000),
      .rdy(const_size_in_1_rsc_rdy),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .const_size_in_1_rsci_oswt(const_size_in_1_rsci_oswt),
      .const_size_in_1_rsci_irdy(const_size_in_1_rsci_irdy),
      .const_size_in_1_rsci_biwt(const_size_in_1_rsci_biwt),
      .const_size_in_1_rsci_bdwt(const_size_in_1_rsci_bdwt),
      .const_size_in_1_rsci_bcwt(const_size_in_1_rsci_bcwt),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
  econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_in_1_rsci_oswt(const_size_in_1_rsci_oswt),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp),
      .const_size_in_1_rsci_biwt(const_size_in_1_rsci_biwt),
      .const_size_in_1_rsci_bdwt(const_size_in_1_rsci_bdwt),
      .const_size_in_1_rsci_bcwt(const_size_in_1_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci (
  clk, rst, layer5_out_rsc_dat, layer5_out_rsc_vld, layer5_out_rsc_rdy, core_wen,
      layer5_out_rsci_oswt, layer5_out_rsci_wen_comp, layer5_out_rsci_idat
);
  input clk;
  input rst;
  output [79:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  input core_wen;
  input layer5_out_rsci_oswt;
  output layer5_out_rsci_wen_comp;
  input [79:0] layer5_out_rsci_idat;


  // Interconnect Declarations
  wire layer5_out_rsci_irdy;
  wire layer5_out_rsci_biwt;
  wire layer5_out_rsci_bdwt;
  wire layer5_out_rsci_bcwt;
  wire layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [79:0] nl_layer5_out_rsci_idat;
  assign nl_layer5_out_rsci_idat = {1'b0 , (layer5_out_rsci_idat[78:72]) , 1'b0 ,
      (layer5_out_rsci_idat[70:64]) , 1'b0 , (layer5_out_rsci_idat[62:56]) , 1'b0
      , (layer5_out_rsci_idat[54:48]) , 1'b0 , (layer5_out_rsci_idat[46:40]) , 1'b0
      , (layer5_out_rsci_idat[38:32]) , 1'b0 , (layer5_out_rsci_idat[30:24]) , 1'b0
      , (layer5_out_rsci_idat[22:16]) , 1'b0 , (layer5_out_rsci_idat[14:8]) , 1'b0
      , (layer5_out_rsci_idat[6:0])};
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd80)) layer5_out_rsci (
      .irdy(layer5_out_rsci_irdy),
      .ivld(layer5_out_rsci_ivld_core_sct),
      .idat(nl_layer5_out_rsci_idat[79:0]),
      .rdy(layer5_out_rsc_rdy),
      .vld(layer5_out_rsc_vld),
      .dat(layer5_out_rsc_dat)
    );
  econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .layer5_out_rsci_oswt(layer5_out_rsci_oswt),
      .layer5_out_rsci_irdy(layer5_out_rsci_irdy),
      .layer5_out_rsci_biwt(layer5_out_rsci_biwt),
      .layer5_out_rsci_bdwt(layer5_out_rsci_bdwt),
      .layer5_out_rsci_bcwt(layer5_out_rsci_bcwt),
      .layer5_out_rsci_ivld_core_sct(layer5_out_rsci_ivld_core_sct)
    );
  econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_dp econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer5_out_rsci_oswt(layer5_out_rsci_oswt),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp),
      .layer5_out_rsci_biwt(layer5_out_rsci_biwt),
      .layer5_out_rsci_bdwt(layer5_out_rsci_bdwt),
      .layer5_out_rsci_bcwt(layer5_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsci (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, core_wen, input_1_rsci_oswt,
      input_1_rsci_wen_comp, input_1_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [383:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  input core_wen;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [383:0] input_1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_1_rsci_biwt;
  wire input_1_rsci_bdwt;
  wire input_1_rsci_bcwt;
  wire input_1_rsci_irdy_core_sct;
  wire input_1_rsci_ivld;
  wire [383:0] input_1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd384)) input_1_rsci (
      .rdy(input_1_rsc_rdy),
      .vld(input_1_rsc_vld),
      .dat(input_1_rsc_dat),
      .irdy(input_1_rsci_irdy_core_sct),
      .ivld(input_1_rsci_ivld),
      .idat(input_1_rsci_idat)
    );
  econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_ctrl econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .input_1_rsci_oswt(input_1_rsci_oswt),
      .input_1_rsci_biwt(input_1_rsci_biwt),
      .input_1_rsci_bdwt(input_1_rsci_bdwt),
      .input_1_rsci_bcwt(input_1_rsci_bcwt),
      .input_1_rsci_irdy_core_sct(input_1_rsci_irdy_core_sct),
      .input_1_rsci_ivld(input_1_rsci_ivld)
    );
  econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_dp econ_4x4_d10_core_input_1_rsci_input_1_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_1_rsci_oswt(input_1_rsci_oswt),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt),
      .input_1_rsci_biwt(input_1_rsci_biwt),
      .input_1_rsci_bdwt(input_1_rsci_bdwt),
      .input_1_rsci_bcwt(input_1_rsci_bcwt),
      .input_1_rsci_idat(input_1_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core
// ------------------------------------------------------------------


module econ_4x4_d10_core (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, input_1_rsc_triosy_lz,
      layer5_out_rsc_dat, layer5_out_rsc_vld, layer5_out_rsc_rdy, layer5_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_rdy, const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld,
      w2_rsc_rdy, w2_rsc_triosy_lz, b2_rsc_dat, b2_rsc_vld, b2_rsc_rdy, b2_rsc_triosy_lz,
      w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, w4_rsc_triosy_lz, b4_rsc_dat, b4_rsc_vld,
      b4_rsc_rdy, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [383:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  output input_1_rsc_triosy_lz;
  output [79:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  output b4_rsc_triosy_lz;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_1_rsci_wen_comp;
  wire [383:0] input_1_rsci_idat_mxwt;
  wire layer5_out_rsci_wen_comp;
  wire const_size_in_1_rsci_wen_comp;
  wire const_size_out_1_rsci_wen_comp;
  wire w2_rsci_wen_comp;
  wire [1727:0] w2_rsci_idat_mxwt;
  wire b2_rsci_wen_comp;
  wire [55:0] b2_rsci_idat_mxwt;
  wire w4_rsci_wen_comp;
  wire [10239:0] w4_rsci_idat_mxwt;
  wire b4_rsci_wen_comp;
  wire [69:0] b4_rsci_idat_mxwt;
  reg [6:0] layer5_out_rsci_idat_78_72;
  reg [6:0] layer5_out_rsci_idat_70_64;
  reg [6:0] layer5_out_rsci_idat_62_56;
  reg [6:0] layer5_out_rsci_idat_54_48;
  reg [6:0] layer5_out_rsci_idat_46_40;
  reg [6:0] layer5_out_rsci_idat_38_32;
  reg [6:0] layer5_out_rsci_idat_30_24;
  reg [6:0] layer5_out_rsci_idat_22_16;
  reg [6:0] layer5_out_rsci_idat_14_8;
  reg [6:0] layer5_out_rsci_idat_6_0;
  wire [1:0] fsm_output;
  wire [7:0] layer4_out_0_sva_1;
  wire [8:0] nl_layer4_out_0_sva_1;
  wire [7:0] MultLoop_1280_MultLoop_acc_3_ncse_sva_1;
  wire [8:0] nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1;
  wire [7:0] nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1;
  wire [8:0] nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [11:0] nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [12:0] nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1;
  wire [12:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1;
  wire [7:0] nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1;
  wire [11:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1;
  wire nnet_relu_layer4_t_result_t_relu_config5_for_if_and_cse;
  reg reg_b4_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1;
  wire [6:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289;

  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[8:0] nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[9:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[7:0] MultLoop_acc_1270_nl;
  wire[8:0] nl_MultLoop_acc_1270_nl;
  wire[7:0] MultLoop_acc_1268_nl;
  wire[8:0] nl_MultLoop_acc_1268_nl;
  wire[7:0] MultLoop_acc_1264_nl;
  wire[8:0] nl_MultLoop_acc_1264_nl;
  wire[7:0] MultLoop_acc_1256_nl;
  wire[8:0] nl_MultLoop_acc_1256_nl;
  wire[7:0] MultLoop_acc_1240_nl;
  wire[8:0] nl_MultLoop_acc_1240_nl;
  wire[7:0] MultLoop_acc_1208_nl;
  wire[8:0] nl_MultLoop_acc_1208_nl;
  wire[7:0] MultLoop_acc_1144_nl;
  wire[8:0] nl_MultLoop_acc_1144_nl;
  wire[14:0] MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1207_nl;
  wire[8:0] nl_MultLoop_acc_1207_nl;
  wire[14:0] MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1239_nl;
  wire[8:0] nl_MultLoop_acc_1239_nl;
  wire[7:0] MultLoop_acc_1206_nl;
  wire[8:0] nl_MultLoop_acc_1206_nl;
  wire[14:0] MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1205_nl;
  wire[8:0] nl_MultLoop_acc_1205_nl;
  wire[14:0] MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1255_nl;
  wire[9:0] nl_MultLoop_acc_1255_nl;
  wire[7:0] MultLoop_acc_1204_nl;
  wire[8:0] nl_MultLoop_acc_1204_nl;
  wire[14:0] MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1203_nl;
  wire[8:0] nl_MultLoop_acc_1203_nl;
  wire[14:0] MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1202_nl;
  wire[8:0] nl_MultLoop_acc_1202_nl;
  wire[14:0] MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1201_nl;
  wire[8:0] nl_MultLoop_acc_1201_nl;
  wire[14:0] MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1263_nl;
  wire[10:0] nl_MultLoop_acc_1263_nl;
  wire[7:0] MultLoop_acc_1196_nl;
  wire[8:0] nl_MultLoop_acc_1196_nl;
  wire[14:0] MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1195_nl;
  wire[8:0] nl_MultLoop_acc_1195_nl;
  wire[14:0] MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1200_nl;
  wire[8:0] nl_MultLoop_acc_1200_nl;
  wire[14:0] MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1199_nl;
  wire[8:0] nl_MultLoop_acc_1199_nl;
  wire[14:0] MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1198_nl;
  wire[8:0] nl_MultLoop_acc_1198_nl;
  wire[14:0] MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1197_nl;
  wire[8:0] nl_MultLoop_acc_1197_nl;
  wire[14:0] MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1194_nl;
  wire[8:0] nl_MultLoop_acc_1194_nl;
  wire[14:0] MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1193_nl;
  wire[8:0] nl_MultLoop_acc_1193_nl;
  wire[14:0] MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1267_nl;
  wire[11:0] nl_MultLoop_acc_1267_nl;
  wire[7:0] MultLoop_acc_1192_nl;
  wire[8:0] nl_MultLoop_acc_1192_nl;
  wire[14:0] MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1191_nl;
  wire[8:0] nl_MultLoop_acc_1191_nl;
  wire[14:0] MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1190_nl;
  wire[8:0] nl_MultLoop_acc_1190_nl;
  wire[14:0] MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1189_nl;
  wire[8:0] nl_MultLoop_acc_1189_nl;
  wire[14:0] MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1188_nl;
  wire[8:0] nl_MultLoop_acc_1188_nl;
  wire[14:0] MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1187_nl;
  wire[8:0] nl_MultLoop_acc_1187_nl;
  wire[14:0] MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1186_nl;
  wire[8:0] nl_MultLoop_acc_1186_nl;
  wire[14:0] MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1185_nl;
  wire[8:0] nl_MultLoop_acc_1185_nl;
  wire[14:0] MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1180_nl;
  wire[8:0] nl_MultLoop_acc_1180_nl;
  wire[14:0] MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1179_nl;
  wire[8:0] nl_MultLoop_acc_1179_nl;
  wire[14:0] MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1178_nl;
  wire[8:0] nl_MultLoop_acc_1178_nl;
  wire[14:0] MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1177_nl;
  wire[8:0] nl_MultLoop_acc_1177_nl;
  wire[14:0] MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1184_nl;
  wire[8:0] nl_MultLoop_acc_1184_nl;
  wire[14:0] MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1183_nl;
  wire[8:0] nl_MultLoop_acc_1183_nl;
  wire[14:0] MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1182_nl;
  wire[8:0] nl_MultLoop_acc_1182_nl;
  wire[14:0] MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1181_nl;
  wire[8:0] nl_MultLoop_acc_1181_nl;
  wire[14:0] MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1269_nl;
  wire[12:0] nl_MultLoop_acc_1269_nl;
  wire[7:0] MultLoop_acc_1172_nl;
  wire[8:0] nl_MultLoop_acc_1172_nl;
  wire[14:0] MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1171_nl;
  wire[8:0] nl_MultLoop_acc_1171_nl;
  wire[14:0] MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1164_nl;
  wire[8:0] nl_MultLoop_acc_1164_nl;
  wire[14:0] MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1163_nl;
  wire[8:0] nl_MultLoop_acc_1163_nl;
  wire[14:0] MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1168_nl;
  wire[8:0] nl_MultLoop_acc_1168_nl;
  wire[14:0] MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1167_nl;
  wire[8:0] nl_MultLoop_acc_1167_nl;
  wire[14:0] MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1148_nl;
  wire[8:0] nl_MultLoop_acc_1148_nl;
  wire[14:0] MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1147_nl;
  wire[8:0] nl_MultLoop_acc_1147_nl;
  wire[14:0] MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1152_nl;
  wire[8:0] nl_MultLoop_acc_1152_nl;
  wire[14:0] MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1151_nl;
  wire[8:0] nl_MultLoop_acc_1151_nl;
  wire[14:0] MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1150_nl;
  wire[8:0] nl_MultLoop_acc_1150_nl;
  wire[14:0] MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1149_nl;
  wire[8:0] nl_MultLoop_acc_1149_nl;
  wire[14:0] MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1160_nl;
  wire[8:0] nl_MultLoop_acc_1160_nl;
  wire[14:0] MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1159_nl;
  wire[8:0] nl_MultLoop_acc_1159_nl;
  wire[14:0] MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1158_nl;
  wire[8:0] nl_MultLoop_acc_1158_nl;
  wire[14:0] MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1157_nl;
  wire[8:0] nl_MultLoop_acc_1157_nl;
  wire[14:0] MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1156_nl;
  wire[8:0] nl_MultLoop_acc_1156_nl;
  wire[14:0] MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1155_nl;
  wire[8:0] nl_MultLoop_acc_1155_nl;
  wire[14:0] MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1154_nl;
  wire[8:0] nl_MultLoop_acc_1154_nl;
  wire[14:0] MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1153_nl;
  wire[8:0] nl_MultLoop_acc_1153_nl;
  wire[14:0] MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1176_nl;
  wire[8:0] nl_MultLoop_acc_1176_nl;
  wire[14:0] MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1175_nl;
  wire[8:0] nl_MultLoop_acc_1175_nl;
  wire[14:0] MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1174_nl;
  wire[8:0] nl_MultLoop_acc_1174_nl;
  wire[14:0] MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1173_nl;
  wire[8:0] nl_MultLoop_acc_1173_nl;
  wire[14:0] MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1170_nl;
  wire[8:0] nl_MultLoop_acc_1170_nl;
  wire[14:0] MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1169_nl;
  wire[8:0] nl_MultLoop_acc_1169_nl;
  wire[14:0] MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1166_nl;
  wire[8:0] nl_MultLoop_acc_1166_nl;
  wire[14:0] MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1165_nl;
  wire[8:0] nl_MultLoop_acc_1165_nl;
  wire[14:0] MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1162_nl;
  wire[8:0] nl_MultLoop_acc_1162_nl;
  wire[14:0] MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1161_nl;
  wire[8:0] nl_MultLoop_acc_1161_nl;
  wire[14:0] MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1146_nl;
  wire[8:0] nl_MultLoop_acc_1146_nl;
  wire[14:0] MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1145_nl;
  wire[8:0] nl_MultLoop_acc_1145_nl;
  wire[14:0] MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1143_nl;
  wire[8:0] nl_MultLoop_acc_1143_nl;
  wire[7:0] MultLoop_acc_1141_nl;
  wire[8:0] nl_MultLoop_acc_1141_nl;
  wire[7:0] MultLoop_acc_1137_nl;
  wire[8:0] nl_MultLoop_acc_1137_nl;
  wire[7:0] MultLoop_acc_1129_nl;
  wire[8:0] nl_MultLoop_acc_1129_nl;
  wire[7:0] MultLoop_acc_1113_nl;
  wire[8:0] nl_MultLoop_acc_1113_nl;
  wire[7:0] MultLoop_acc_1081_nl;
  wire[8:0] nl_MultLoop_acc_1081_nl;
  wire[7:0] MultLoop_acc_1017_nl;
  wire[8:0] nl_MultLoop_acc_1017_nl;
  wire[14:0] MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1080_nl;
  wire[8:0] nl_MultLoop_acc_1080_nl;
  wire[14:0] MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1112_nl;
  wire[8:0] nl_MultLoop_acc_1112_nl;
  wire[7:0] MultLoop_acc_1079_nl;
  wire[8:0] nl_MultLoop_acc_1079_nl;
  wire[14:0] MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1078_nl;
  wire[8:0] nl_MultLoop_acc_1078_nl;
  wire[14:0] MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1128_nl;
  wire[9:0] nl_MultLoop_acc_1128_nl;
  wire[7:0] MultLoop_acc_1077_nl;
  wire[8:0] nl_MultLoop_acc_1077_nl;
  wire[14:0] MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1076_nl;
  wire[8:0] nl_MultLoop_acc_1076_nl;
  wire[14:0] MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1075_nl;
  wire[8:0] nl_MultLoop_acc_1075_nl;
  wire[14:0] MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1074_nl;
  wire[8:0] nl_MultLoop_acc_1074_nl;
  wire[14:0] MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1136_nl;
  wire[10:0] nl_MultLoop_acc_1136_nl;
  wire[7:0] MultLoop_acc_1069_nl;
  wire[8:0] nl_MultLoop_acc_1069_nl;
  wire[14:0] MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1068_nl;
  wire[8:0] nl_MultLoop_acc_1068_nl;
  wire[14:0] MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1073_nl;
  wire[8:0] nl_MultLoop_acc_1073_nl;
  wire[14:0] MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1072_nl;
  wire[8:0] nl_MultLoop_acc_1072_nl;
  wire[14:0] MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1071_nl;
  wire[8:0] nl_MultLoop_acc_1071_nl;
  wire[14:0] MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1070_nl;
  wire[8:0] nl_MultLoop_acc_1070_nl;
  wire[14:0] MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1067_nl;
  wire[8:0] nl_MultLoop_acc_1067_nl;
  wire[14:0] MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1066_nl;
  wire[8:0] nl_MultLoop_acc_1066_nl;
  wire[14:0] MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1140_nl;
  wire[11:0] nl_MultLoop_acc_1140_nl;
  wire[7:0] MultLoop_acc_1065_nl;
  wire[8:0] nl_MultLoop_acc_1065_nl;
  wire[14:0] MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1064_nl;
  wire[8:0] nl_MultLoop_acc_1064_nl;
  wire[14:0] MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1063_nl;
  wire[8:0] nl_MultLoop_acc_1063_nl;
  wire[14:0] MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1062_nl;
  wire[8:0] nl_MultLoop_acc_1062_nl;
  wire[14:0] MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1061_nl;
  wire[8:0] nl_MultLoop_acc_1061_nl;
  wire[14:0] MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1060_nl;
  wire[8:0] nl_MultLoop_acc_1060_nl;
  wire[14:0] MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1059_nl;
  wire[8:0] nl_MultLoop_acc_1059_nl;
  wire[14:0] MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1058_nl;
  wire[8:0] nl_MultLoop_acc_1058_nl;
  wire[14:0] MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1053_nl;
  wire[8:0] nl_MultLoop_acc_1053_nl;
  wire[14:0] MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1052_nl;
  wire[8:0] nl_MultLoop_acc_1052_nl;
  wire[14:0] MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1051_nl;
  wire[8:0] nl_MultLoop_acc_1051_nl;
  wire[14:0] MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1050_nl;
  wire[8:0] nl_MultLoop_acc_1050_nl;
  wire[14:0] MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1057_nl;
  wire[8:0] nl_MultLoop_acc_1057_nl;
  wire[14:0] MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1056_nl;
  wire[8:0] nl_MultLoop_acc_1056_nl;
  wire[14:0] MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1055_nl;
  wire[8:0] nl_MultLoop_acc_1055_nl;
  wire[14:0] MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1054_nl;
  wire[8:0] nl_MultLoop_acc_1054_nl;
  wire[14:0] MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1142_nl;
  wire[12:0] nl_MultLoop_acc_1142_nl;
  wire[7:0] MultLoop_acc_1045_nl;
  wire[8:0] nl_MultLoop_acc_1045_nl;
  wire[14:0] MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1044_nl;
  wire[8:0] nl_MultLoop_acc_1044_nl;
  wire[14:0] MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1037_nl;
  wire[8:0] nl_MultLoop_acc_1037_nl;
  wire[14:0] MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1036_nl;
  wire[8:0] nl_MultLoop_acc_1036_nl;
  wire[14:0] MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1041_nl;
  wire[8:0] nl_MultLoop_acc_1041_nl;
  wire[14:0] MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1040_nl;
  wire[8:0] nl_MultLoop_acc_1040_nl;
  wire[14:0] MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1021_nl;
  wire[8:0] nl_MultLoop_acc_1021_nl;
  wire[14:0] MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1020_nl;
  wire[8:0] nl_MultLoop_acc_1020_nl;
  wire[14:0] MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1025_nl;
  wire[8:0] nl_MultLoop_acc_1025_nl;
  wire[14:0] MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1024_nl;
  wire[8:0] nl_MultLoop_acc_1024_nl;
  wire[14:0] MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1023_nl;
  wire[8:0] nl_MultLoop_acc_1023_nl;
  wire[14:0] MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1022_nl;
  wire[8:0] nl_MultLoop_acc_1022_nl;
  wire[14:0] MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1033_nl;
  wire[8:0] nl_MultLoop_acc_1033_nl;
  wire[14:0] MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1032_nl;
  wire[8:0] nl_MultLoop_acc_1032_nl;
  wire[14:0] MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1031_nl;
  wire[8:0] nl_MultLoop_acc_1031_nl;
  wire[14:0] MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1030_nl;
  wire[8:0] nl_MultLoop_acc_1030_nl;
  wire[14:0] MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1029_nl;
  wire[8:0] nl_MultLoop_acc_1029_nl;
  wire[14:0] MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1028_nl;
  wire[8:0] nl_MultLoop_acc_1028_nl;
  wire[14:0] MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1027_nl;
  wire[8:0] nl_MultLoop_acc_1027_nl;
  wire[14:0] MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1026_nl;
  wire[8:0] nl_MultLoop_acc_1026_nl;
  wire[14:0] MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1049_nl;
  wire[8:0] nl_MultLoop_acc_1049_nl;
  wire[14:0] MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1048_nl;
  wire[8:0] nl_MultLoop_acc_1048_nl;
  wire[14:0] MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1047_nl;
  wire[8:0] nl_MultLoop_acc_1047_nl;
  wire[14:0] MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1046_nl;
  wire[8:0] nl_MultLoop_acc_1046_nl;
  wire[14:0] MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1043_nl;
  wire[8:0] nl_MultLoop_acc_1043_nl;
  wire[14:0] MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1042_nl;
  wire[8:0] nl_MultLoop_acc_1042_nl;
  wire[14:0] MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1039_nl;
  wire[8:0] nl_MultLoop_acc_1039_nl;
  wire[14:0] MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1038_nl;
  wire[8:0] nl_MultLoop_acc_1038_nl;
  wire[14:0] MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1035_nl;
  wire[8:0] nl_MultLoop_acc_1035_nl;
  wire[14:0] MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1034_nl;
  wire[8:0] nl_MultLoop_acc_1034_nl;
  wire[14:0] MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1019_nl;
  wire[8:0] nl_MultLoop_acc_1019_nl;
  wire[14:0] MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1018_nl;
  wire[8:0] nl_MultLoop_acc_1018_nl;
  wire[14:0] MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_nl;
  wire[8:0] nl_MultLoop_acc_nl;
  wire[7:0] MultLoop_acc_127_nl;
  wire[8:0] nl_MultLoop_acc_127_nl;
  wire[7:0] MultLoop_acc_125_nl;
  wire[8:0] nl_MultLoop_acc_125_nl;
  wire[7:0] MultLoop_acc_121_nl;
  wire[8:0] nl_MultLoop_acc_121_nl;
  wire[7:0] MultLoop_acc_113_nl;
  wire[8:0] nl_MultLoop_acc_113_nl;
  wire[7:0] MultLoop_acc_97_nl;
  wire[8:0] nl_MultLoop_acc_97_nl;
  wire[7:0] MultLoop_acc_65_nl;
  wire[8:0] nl_MultLoop_acc_65_nl;
  wire[14:0] MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_64_nl;
  wire[8:0] nl_MultLoop_acc_64_nl;
  wire[14:0] MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_96_nl;
  wire[8:0] nl_MultLoop_acc_96_nl;
  wire[7:0] MultLoop_acc_63_nl;
  wire[8:0] nl_MultLoop_acc_63_nl;
  wire[14:0] MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_62_nl;
  wire[8:0] nl_MultLoop_acc_62_nl;
  wire[14:0] MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_112_nl;
  wire[9:0] nl_MultLoop_acc_112_nl;
  wire[7:0] MultLoop_acc_61_nl;
  wire[8:0] nl_MultLoop_acc_61_nl;
  wire[14:0] MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_60_nl;
  wire[8:0] nl_MultLoop_acc_60_nl;
  wire[14:0] MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_59_nl;
  wire[8:0] nl_MultLoop_acc_59_nl;
  wire[14:0] MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_58_nl;
  wire[8:0] nl_MultLoop_acc_58_nl;
  wire[14:0] MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_120_nl;
  wire[10:0] nl_MultLoop_acc_120_nl;
  wire[7:0] MultLoop_acc_53_nl;
  wire[8:0] nl_MultLoop_acc_53_nl;
  wire[14:0] MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_52_nl;
  wire[8:0] nl_MultLoop_acc_52_nl;
  wire[14:0] MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_57_nl;
  wire[8:0] nl_MultLoop_acc_57_nl;
  wire[14:0] MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_56_nl;
  wire[8:0] nl_MultLoop_acc_56_nl;
  wire[14:0] MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_55_nl;
  wire[8:0] nl_MultLoop_acc_55_nl;
  wire[14:0] MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_54_nl;
  wire[8:0] nl_MultLoop_acc_54_nl;
  wire[14:0] MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_51_nl;
  wire[8:0] nl_MultLoop_acc_51_nl;
  wire[14:0] MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_50_nl;
  wire[8:0] nl_MultLoop_acc_50_nl;
  wire[14:0] MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_124_nl;
  wire[11:0] nl_MultLoop_acc_124_nl;
  wire[7:0] MultLoop_acc_49_nl;
  wire[8:0] nl_MultLoop_acc_49_nl;
  wire[14:0] MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_48_nl;
  wire[8:0] nl_MultLoop_acc_48_nl;
  wire[14:0] MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_47_nl;
  wire[8:0] nl_MultLoop_acc_47_nl;
  wire[14:0] MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_46_nl;
  wire[8:0] nl_MultLoop_acc_46_nl;
  wire[14:0] MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_45_nl;
  wire[8:0] nl_MultLoop_acc_45_nl;
  wire[14:0] MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_44_nl;
  wire[8:0] nl_MultLoop_acc_44_nl;
  wire[14:0] MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_43_nl;
  wire[8:0] nl_MultLoop_acc_43_nl;
  wire[14:0] MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_42_nl;
  wire[8:0] nl_MultLoop_acc_42_nl;
  wire[14:0] MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_37_nl;
  wire[8:0] nl_MultLoop_acc_37_nl;
  wire[14:0] MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_36_nl;
  wire[8:0] nl_MultLoop_acc_36_nl;
  wire[14:0] MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_35_nl;
  wire[8:0] nl_MultLoop_acc_35_nl;
  wire[14:0] MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_34_nl;
  wire[8:0] nl_MultLoop_acc_34_nl;
  wire[14:0] MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_41_nl;
  wire[8:0] nl_MultLoop_acc_41_nl;
  wire[14:0] MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_40_nl;
  wire[8:0] nl_MultLoop_acc_40_nl;
  wire[14:0] MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_39_nl;
  wire[8:0] nl_MultLoop_acc_39_nl;
  wire[14:0] MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_38_nl;
  wire[8:0] nl_MultLoop_acc_38_nl;
  wire[14:0] MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_126_nl;
  wire[12:0] nl_MultLoop_acc_126_nl;
  wire[7:0] MultLoop_acc_29_nl;
  wire[8:0] nl_MultLoop_acc_29_nl;
  wire[14:0] MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_28_nl;
  wire[8:0] nl_MultLoop_acc_28_nl;
  wire[14:0] MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_21_nl;
  wire[8:0] nl_MultLoop_acc_21_nl;
  wire[14:0] MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_20_nl;
  wire[8:0] nl_MultLoop_acc_20_nl;
  wire[14:0] MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_25_nl;
  wire[8:0] nl_MultLoop_acc_25_nl;
  wire[14:0] MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_24_nl;
  wire[8:0] nl_MultLoop_acc_24_nl;
  wire[14:0] MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_5_nl;
  wire[8:0] nl_MultLoop_acc_5_nl;
  wire[14:0] MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_4_nl;
  wire[8:0] nl_MultLoop_acc_4_nl;
  wire[14:0] MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_9_nl;
  wire[8:0] nl_MultLoop_acc_9_nl;
  wire[14:0] MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_8_nl;
  wire[8:0] nl_MultLoop_acc_8_nl;
  wire[14:0] MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_7_nl;
  wire[8:0] nl_MultLoop_acc_7_nl;
  wire[14:0] MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_6_nl;
  wire[8:0] nl_MultLoop_acc_6_nl;
  wire[14:0] MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_17_nl;
  wire[8:0] nl_MultLoop_acc_17_nl;
  wire[14:0] MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_16_nl;
  wire[8:0] nl_MultLoop_acc_16_nl;
  wire[14:0] MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_15_nl;
  wire[8:0] nl_MultLoop_acc_15_nl;
  wire[14:0] MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_14_nl;
  wire[8:0] nl_MultLoop_acc_14_nl;
  wire[14:0] MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_13_nl;
  wire[8:0] nl_MultLoop_acc_13_nl;
  wire[14:0] MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_12_nl;
  wire[8:0] nl_MultLoop_acc_12_nl;
  wire[14:0] MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_11_nl;
  wire[8:0] nl_MultLoop_acc_11_nl;
  wire[14:0] MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_10_nl;
  wire[8:0] nl_MultLoop_acc_10_nl;
  wire[14:0] MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_33_nl;
  wire[8:0] nl_MultLoop_acc_33_nl;
  wire[14:0] MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_32_nl;
  wire[8:0] nl_MultLoop_acc_32_nl;
  wire[14:0] MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_31_nl;
  wire[8:0] nl_MultLoop_acc_31_nl;
  wire[14:0] MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_30_nl;
  wire[8:0] nl_MultLoop_acc_30_nl;
  wire[14:0] MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_27_nl;
  wire[8:0] nl_MultLoop_acc_27_nl;
  wire[14:0] MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_26_nl;
  wire[8:0] nl_MultLoop_acc_26_nl;
  wire[14:0] MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_23_nl;
  wire[8:0] nl_MultLoop_acc_23_nl;
  wire[14:0] MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_22_nl;
  wire[8:0] nl_MultLoop_acc_22_nl;
  wire[14:0] MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_19_nl;
  wire[8:0] nl_MultLoop_acc_19_nl;
  wire[14:0] MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_18_nl;
  wire[8:0] nl_MultLoop_acc_18_nl;
  wire[14:0] MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_3_nl;
  wire[8:0] nl_MultLoop_acc_3_nl;
  wire[14:0] MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_2_nl;
  wire[8:0] nl_MultLoop_acc_2_nl;
  wire[14:0] MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1016_nl;
  wire[8:0] nl_MultLoop_acc_1016_nl;
  wire[7:0] MultLoop_acc_1014_nl;
  wire[8:0] nl_MultLoop_acc_1014_nl;
  wire[7:0] MultLoop_acc_1010_nl;
  wire[8:0] nl_MultLoop_acc_1010_nl;
  wire[7:0] MultLoop_acc_1002_nl;
  wire[8:0] nl_MultLoop_acc_1002_nl;
  wire[7:0] MultLoop_acc_986_nl;
  wire[8:0] nl_MultLoop_acc_986_nl;
  wire[7:0] MultLoop_acc_954_nl;
  wire[8:0] nl_MultLoop_acc_954_nl;
  wire[7:0] MultLoop_acc_890_nl;
  wire[8:0] nl_MultLoop_acc_890_nl;
  wire[14:0] MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_953_nl;
  wire[8:0] nl_MultLoop_acc_953_nl;
  wire[14:0] MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_985_nl;
  wire[8:0] nl_MultLoop_acc_985_nl;
  wire[7:0] MultLoop_acc_952_nl;
  wire[8:0] nl_MultLoop_acc_952_nl;
  wire[14:0] MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_951_nl;
  wire[8:0] nl_MultLoop_acc_951_nl;
  wire[14:0] MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1001_nl;
  wire[9:0] nl_MultLoop_acc_1001_nl;
  wire[7:0] MultLoop_acc_950_nl;
  wire[8:0] nl_MultLoop_acc_950_nl;
  wire[14:0] MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_949_nl;
  wire[8:0] nl_MultLoop_acc_949_nl;
  wire[14:0] MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_948_nl;
  wire[8:0] nl_MultLoop_acc_948_nl;
  wire[14:0] MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_947_nl;
  wire[8:0] nl_MultLoop_acc_947_nl;
  wire[14:0] MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1009_nl;
  wire[10:0] nl_MultLoop_acc_1009_nl;
  wire[7:0] MultLoop_acc_942_nl;
  wire[8:0] nl_MultLoop_acc_942_nl;
  wire[14:0] MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_941_nl;
  wire[8:0] nl_MultLoop_acc_941_nl;
  wire[14:0] MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_946_nl;
  wire[8:0] nl_MultLoop_acc_946_nl;
  wire[14:0] MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_945_nl;
  wire[8:0] nl_MultLoop_acc_945_nl;
  wire[14:0] MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_944_nl;
  wire[8:0] nl_MultLoop_acc_944_nl;
  wire[14:0] MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_943_nl;
  wire[8:0] nl_MultLoop_acc_943_nl;
  wire[14:0] MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_940_nl;
  wire[8:0] nl_MultLoop_acc_940_nl;
  wire[14:0] MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_939_nl;
  wire[8:0] nl_MultLoop_acc_939_nl;
  wire[14:0] MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1013_nl;
  wire[11:0] nl_MultLoop_acc_1013_nl;
  wire[7:0] MultLoop_acc_938_nl;
  wire[8:0] nl_MultLoop_acc_938_nl;
  wire[14:0] MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_937_nl;
  wire[8:0] nl_MultLoop_acc_937_nl;
  wire[14:0] MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_936_nl;
  wire[8:0] nl_MultLoop_acc_936_nl;
  wire[14:0] MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_935_nl;
  wire[8:0] nl_MultLoop_acc_935_nl;
  wire[14:0] MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_934_nl;
  wire[8:0] nl_MultLoop_acc_934_nl;
  wire[14:0] MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_933_nl;
  wire[8:0] nl_MultLoop_acc_933_nl;
  wire[14:0] MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_932_nl;
  wire[8:0] nl_MultLoop_acc_932_nl;
  wire[14:0] MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_931_nl;
  wire[8:0] nl_MultLoop_acc_931_nl;
  wire[14:0] MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_926_nl;
  wire[8:0] nl_MultLoop_acc_926_nl;
  wire[14:0] MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_925_nl;
  wire[8:0] nl_MultLoop_acc_925_nl;
  wire[14:0] MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_924_nl;
  wire[8:0] nl_MultLoop_acc_924_nl;
  wire[14:0] MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_923_nl;
  wire[8:0] nl_MultLoop_acc_923_nl;
  wire[14:0] MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_930_nl;
  wire[8:0] nl_MultLoop_acc_930_nl;
  wire[14:0] MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_929_nl;
  wire[8:0] nl_MultLoop_acc_929_nl;
  wire[14:0] MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_928_nl;
  wire[8:0] nl_MultLoop_acc_928_nl;
  wire[14:0] MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_927_nl;
  wire[8:0] nl_MultLoop_acc_927_nl;
  wire[14:0] MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_1015_nl;
  wire[12:0] nl_MultLoop_acc_1015_nl;
  wire[7:0] MultLoop_acc_918_nl;
  wire[8:0] nl_MultLoop_acc_918_nl;
  wire[14:0] MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_917_nl;
  wire[8:0] nl_MultLoop_acc_917_nl;
  wire[14:0] MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_910_nl;
  wire[8:0] nl_MultLoop_acc_910_nl;
  wire[14:0] MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_909_nl;
  wire[8:0] nl_MultLoop_acc_909_nl;
  wire[14:0] MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_914_nl;
  wire[8:0] nl_MultLoop_acc_914_nl;
  wire[14:0] MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_913_nl;
  wire[8:0] nl_MultLoop_acc_913_nl;
  wire[14:0] MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_894_nl;
  wire[8:0] nl_MultLoop_acc_894_nl;
  wire[14:0] MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_893_nl;
  wire[8:0] nl_MultLoop_acc_893_nl;
  wire[14:0] MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_898_nl;
  wire[8:0] nl_MultLoop_acc_898_nl;
  wire[14:0] MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_897_nl;
  wire[8:0] nl_MultLoop_acc_897_nl;
  wire[14:0] MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_896_nl;
  wire[8:0] nl_MultLoop_acc_896_nl;
  wire[14:0] MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_895_nl;
  wire[8:0] nl_MultLoop_acc_895_nl;
  wire[14:0] MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_906_nl;
  wire[8:0] nl_MultLoop_acc_906_nl;
  wire[14:0] MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_905_nl;
  wire[8:0] nl_MultLoop_acc_905_nl;
  wire[14:0] MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_904_nl;
  wire[8:0] nl_MultLoop_acc_904_nl;
  wire[14:0] MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_903_nl;
  wire[8:0] nl_MultLoop_acc_903_nl;
  wire[14:0] MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_902_nl;
  wire[8:0] nl_MultLoop_acc_902_nl;
  wire[14:0] MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_901_nl;
  wire[8:0] nl_MultLoop_acc_901_nl;
  wire[14:0] MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_900_nl;
  wire[8:0] nl_MultLoop_acc_900_nl;
  wire[14:0] MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_899_nl;
  wire[8:0] nl_MultLoop_acc_899_nl;
  wire[14:0] MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_922_nl;
  wire[8:0] nl_MultLoop_acc_922_nl;
  wire[14:0] MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_921_nl;
  wire[8:0] nl_MultLoop_acc_921_nl;
  wire[14:0] MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_920_nl;
  wire[8:0] nl_MultLoop_acc_920_nl;
  wire[14:0] MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_919_nl;
  wire[8:0] nl_MultLoop_acc_919_nl;
  wire[14:0] MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_916_nl;
  wire[8:0] nl_MultLoop_acc_916_nl;
  wire[14:0] MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_915_nl;
  wire[8:0] nl_MultLoop_acc_915_nl;
  wire[14:0] MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_912_nl;
  wire[8:0] nl_MultLoop_acc_912_nl;
  wire[14:0] MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_911_nl;
  wire[8:0] nl_MultLoop_acc_911_nl;
  wire[14:0] MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_908_nl;
  wire[8:0] nl_MultLoop_acc_908_nl;
  wire[14:0] MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_907_nl;
  wire[8:0] nl_MultLoop_acc_907_nl;
  wire[14:0] MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_892_nl;
  wire[8:0] nl_MultLoop_acc_892_nl;
  wire[14:0] MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_891_nl;
  wire[8:0] nl_MultLoop_acc_891_nl;
  wire[14:0] MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_254_nl;
  wire[8:0] nl_MultLoop_acc_254_nl;
  wire[7:0] MultLoop_acc_252_nl;
  wire[8:0] nl_MultLoop_acc_252_nl;
  wire[7:0] MultLoop_acc_248_nl;
  wire[8:0] nl_MultLoop_acc_248_nl;
  wire[7:0] MultLoop_acc_240_nl;
  wire[8:0] nl_MultLoop_acc_240_nl;
  wire[7:0] MultLoop_acc_224_nl;
  wire[8:0] nl_MultLoop_acc_224_nl;
  wire[7:0] MultLoop_acc_192_nl;
  wire[8:0] nl_MultLoop_acc_192_nl;
  wire[7:0] MultLoop_acc_128_nl;
  wire[8:0] nl_MultLoop_acc_128_nl;
  wire[14:0] MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_191_nl;
  wire[8:0] nl_MultLoop_acc_191_nl;
  wire[14:0] MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_223_nl;
  wire[8:0] nl_MultLoop_acc_223_nl;
  wire[7:0] MultLoop_acc_190_nl;
  wire[8:0] nl_MultLoop_acc_190_nl;
  wire[14:0] MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_189_nl;
  wire[8:0] nl_MultLoop_acc_189_nl;
  wire[14:0] MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_239_nl;
  wire[9:0] nl_MultLoop_acc_239_nl;
  wire[7:0] MultLoop_acc_188_nl;
  wire[8:0] nl_MultLoop_acc_188_nl;
  wire[14:0] MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_187_nl;
  wire[8:0] nl_MultLoop_acc_187_nl;
  wire[14:0] MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_186_nl;
  wire[8:0] nl_MultLoop_acc_186_nl;
  wire[14:0] MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_185_nl;
  wire[8:0] nl_MultLoop_acc_185_nl;
  wire[14:0] MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_247_nl;
  wire[10:0] nl_MultLoop_acc_247_nl;
  wire[7:0] MultLoop_acc_180_nl;
  wire[8:0] nl_MultLoop_acc_180_nl;
  wire[14:0] MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_179_nl;
  wire[8:0] nl_MultLoop_acc_179_nl;
  wire[14:0] MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_184_nl;
  wire[8:0] nl_MultLoop_acc_184_nl;
  wire[14:0] MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_183_nl;
  wire[8:0] nl_MultLoop_acc_183_nl;
  wire[14:0] MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_182_nl;
  wire[8:0] nl_MultLoop_acc_182_nl;
  wire[14:0] MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_181_nl;
  wire[8:0] nl_MultLoop_acc_181_nl;
  wire[14:0] MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_178_nl;
  wire[8:0] nl_MultLoop_acc_178_nl;
  wire[14:0] MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_177_nl;
  wire[8:0] nl_MultLoop_acc_177_nl;
  wire[14:0] MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_251_nl;
  wire[11:0] nl_MultLoop_acc_251_nl;
  wire[7:0] MultLoop_acc_176_nl;
  wire[8:0] nl_MultLoop_acc_176_nl;
  wire[14:0] MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_175_nl;
  wire[8:0] nl_MultLoop_acc_175_nl;
  wire[14:0] MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_174_nl;
  wire[8:0] nl_MultLoop_acc_174_nl;
  wire[14:0] MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_173_nl;
  wire[8:0] nl_MultLoop_acc_173_nl;
  wire[14:0] MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_172_nl;
  wire[8:0] nl_MultLoop_acc_172_nl;
  wire[14:0] MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_171_nl;
  wire[8:0] nl_MultLoop_acc_171_nl;
  wire[14:0] MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_170_nl;
  wire[8:0] nl_MultLoop_acc_170_nl;
  wire[14:0] MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_169_nl;
  wire[8:0] nl_MultLoop_acc_169_nl;
  wire[14:0] MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_164_nl;
  wire[8:0] nl_MultLoop_acc_164_nl;
  wire[14:0] MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_163_nl;
  wire[8:0] nl_MultLoop_acc_163_nl;
  wire[14:0] MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_162_nl;
  wire[8:0] nl_MultLoop_acc_162_nl;
  wire[14:0] MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_161_nl;
  wire[8:0] nl_MultLoop_acc_161_nl;
  wire[14:0] MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_168_nl;
  wire[8:0] nl_MultLoop_acc_168_nl;
  wire[14:0] MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_167_nl;
  wire[8:0] nl_MultLoop_acc_167_nl;
  wire[14:0] MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_166_nl;
  wire[8:0] nl_MultLoop_acc_166_nl;
  wire[14:0] MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_165_nl;
  wire[8:0] nl_MultLoop_acc_165_nl;
  wire[14:0] MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_253_nl;
  wire[12:0] nl_MultLoop_acc_253_nl;
  wire[7:0] MultLoop_acc_156_nl;
  wire[8:0] nl_MultLoop_acc_156_nl;
  wire[14:0] MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_155_nl;
  wire[8:0] nl_MultLoop_acc_155_nl;
  wire[14:0] MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_148_nl;
  wire[8:0] nl_MultLoop_acc_148_nl;
  wire[14:0] MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_147_nl;
  wire[8:0] nl_MultLoop_acc_147_nl;
  wire[14:0] MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_152_nl;
  wire[8:0] nl_MultLoop_acc_152_nl;
  wire[14:0] MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_151_nl;
  wire[8:0] nl_MultLoop_acc_151_nl;
  wire[14:0] MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_132_nl;
  wire[8:0] nl_MultLoop_acc_132_nl;
  wire[14:0] MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_131_nl;
  wire[8:0] nl_MultLoop_acc_131_nl;
  wire[14:0] MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_136_nl;
  wire[8:0] nl_MultLoop_acc_136_nl;
  wire[14:0] MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_135_nl;
  wire[8:0] nl_MultLoop_acc_135_nl;
  wire[14:0] MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_134_nl;
  wire[8:0] nl_MultLoop_acc_134_nl;
  wire[14:0] MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_133_nl;
  wire[8:0] nl_MultLoop_acc_133_nl;
  wire[14:0] MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_144_nl;
  wire[8:0] nl_MultLoop_acc_144_nl;
  wire[14:0] MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_143_nl;
  wire[8:0] nl_MultLoop_acc_143_nl;
  wire[14:0] MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_142_nl;
  wire[8:0] nl_MultLoop_acc_142_nl;
  wire[14:0] MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_141_nl;
  wire[8:0] nl_MultLoop_acc_141_nl;
  wire[14:0] MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_140_nl;
  wire[8:0] nl_MultLoop_acc_140_nl;
  wire[14:0] MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_139_nl;
  wire[8:0] nl_MultLoop_acc_139_nl;
  wire[14:0] MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_138_nl;
  wire[8:0] nl_MultLoop_acc_138_nl;
  wire[14:0] MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_137_nl;
  wire[8:0] nl_MultLoop_acc_137_nl;
  wire[14:0] MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_160_nl;
  wire[8:0] nl_MultLoop_acc_160_nl;
  wire[14:0] MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_159_nl;
  wire[8:0] nl_MultLoop_acc_159_nl;
  wire[14:0] MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_158_nl;
  wire[8:0] nl_MultLoop_acc_158_nl;
  wire[14:0] MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_157_nl;
  wire[8:0] nl_MultLoop_acc_157_nl;
  wire[14:0] MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_154_nl;
  wire[8:0] nl_MultLoop_acc_154_nl;
  wire[14:0] MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_153_nl;
  wire[8:0] nl_MultLoop_acc_153_nl;
  wire[14:0] MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_150_nl;
  wire[8:0] nl_MultLoop_acc_150_nl;
  wire[14:0] MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_149_nl;
  wire[8:0] nl_MultLoop_acc_149_nl;
  wire[14:0] MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_146_nl;
  wire[8:0] nl_MultLoop_acc_146_nl;
  wire[14:0] MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_145_nl;
  wire[8:0] nl_MultLoop_acc_145_nl;
  wire[14:0] MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_130_nl;
  wire[8:0] nl_MultLoop_acc_130_nl;
  wire[14:0] MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_129_nl;
  wire[8:0] nl_MultLoop_acc_129_nl;
  wire[14:0] MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_889_nl;
  wire[8:0] nl_MultLoop_acc_889_nl;
  wire[7:0] MultLoop_acc_887_nl;
  wire[8:0] nl_MultLoop_acc_887_nl;
  wire[7:0] MultLoop_acc_883_nl;
  wire[8:0] nl_MultLoop_acc_883_nl;
  wire[7:0] MultLoop_acc_875_nl;
  wire[8:0] nl_MultLoop_acc_875_nl;
  wire[7:0] MultLoop_acc_859_nl;
  wire[8:0] nl_MultLoop_acc_859_nl;
  wire[7:0] MultLoop_acc_827_nl;
  wire[8:0] nl_MultLoop_acc_827_nl;
  wire[7:0] MultLoop_acc_763_nl;
  wire[8:0] nl_MultLoop_acc_763_nl;
  wire[14:0] MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_826_nl;
  wire[8:0] nl_MultLoop_acc_826_nl;
  wire[14:0] MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_858_nl;
  wire[8:0] nl_MultLoop_acc_858_nl;
  wire[7:0] MultLoop_acc_825_nl;
  wire[8:0] nl_MultLoop_acc_825_nl;
  wire[14:0] MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_824_nl;
  wire[8:0] nl_MultLoop_acc_824_nl;
  wire[14:0] MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_874_nl;
  wire[9:0] nl_MultLoop_acc_874_nl;
  wire[7:0] MultLoop_acc_823_nl;
  wire[8:0] nl_MultLoop_acc_823_nl;
  wire[14:0] MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_822_nl;
  wire[8:0] nl_MultLoop_acc_822_nl;
  wire[14:0] MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_821_nl;
  wire[8:0] nl_MultLoop_acc_821_nl;
  wire[14:0] MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_820_nl;
  wire[8:0] nl_MultLoop_acc_820_nl;
  wire[14:0] MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_882_nl;
  wire[10:0] nl_MultLoop_acc_882_nl;
  wire[7:0] MultLoop_acc_815_nl;
  wire[8:0] nl_MultLoop_acc_815_nl;
  wire[14:0] MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_814_nl;
  wire[8:0] nl_MultLoop_acc_814_nl;
  wire[14:0] MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_819_nl;
  wire[8:0] nl_MultLoop_acc_819_nl;
  wire[14:0] MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_818_nl;
  wire[8:0] nl_MultLoop_acc_818_nl;
  wire[14:0] MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_817_nl;
  wire[8:0] nl_MultLoop_acc_817_nl;
  wire[14:0] MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_816_nl;
  wire[8:0] nl_MultLoop_acc_816_nl;
  wire[14:0] MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_813_nl;
  wire[8:0] nl_MultLoop_acc_813_nl;
  wire[14:0] MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_812_nl;
  wire[8:0] nl_MultLoop_acc_812_nl;
  wire[14:0] MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_886_nl;
  wire[11:0] nl_MultLoop_acc_886_nl;
  wire[7:0] MultLoop_acc_811_nl;
  wire[8:0] nl_MultLoop_acc_811_nl;
  wire[14:0] MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_810_nl;
  wire[8:0] nl_MultLoop_acc_810_nl;
  wire[14:0] MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_809_nl;
  wire[8:0] nl_MultLoop_acc_809_nl;
  wire[14:0] MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_808_nl;
  wire[8:0] nl_MultLoop_acc_808_nl;
  wire[14:0] MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_807_nl;
  wire[8:0] nl_MultLoop_acc_807_nl;
  wire[14:0] MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_806_nl;
  wire[8:0] nl_MultLoop_acc_806_nl;
  wire[14:0] MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_805_nl;
  wire[8:0] nl_MultLoop_acc_805_nl;
  wire[14:0] MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_804_nl;
  wire[8:0] nl_MultLoop_acc_804_nl;
  wire[14:0] MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_799_nl;
  wire[8:0] nl_MultLoop_acc_799_nl;
  wire[14:0] MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_798_nl;
  wire[8:0] nl_MultLoop_acc_798_nl;
  wire[14:0] MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_797_nl;
  wire[8:0] nl_MultLoop_acc_797_nl;
  wire[14:0] MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_796_nl;
  wire[8:0] nl_MultLoop_acc_796_nl;
  wire[14:0] MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_803_nl;
  wire[8:0] nl_MultLoop_acc_803_nl;
  wire[14:0] MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_802_nl;
  wire[8:0] nl_MultLoop_acc_802_nl;
  wire[14:0] MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_801_nl;
  wire[8:0] nl_MultLoop_acc_801_nl;
  wire[14:0] MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_800_nl;
  wire[8:0] nl_MultLoop_acc_800_nl;
  wire[14:0] MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_888_nl;
  wire[12:0] nl_MultLoop_acc_888_nl;
  wire[7:0] MultLoop_acc_791_nl;
  wire[8:0] nl_MultLoop_acc_791_nl;
  wire[14:0] MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_790_nl;
  wire[8:0] nl_MultLoop_acc_790_nl;
  wire[14:0] MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_783_nl;
  wire[8:0] nl_MultLoop_acc_783_nl;
  wire[14:0] MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_782_nl;
  wire[8:0] nl_MultLoop_acc_782_nl;
  wire[14:0] MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_787_nl;
  wire[8:0] nl_MultLoop_acc_787_nl;
  wire[14:0] MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_786_nl;
  wire[8:0] nl_MultLoop_acc_786_nl;
  wire[14:0] MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_767_nl;
  wire[8:0] nl_MultLoop_acc_767_nl;
  wire[14:0] MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_766_nl;
  wire[8:0] nl_MultLoop_acc_766_nl;
  wire[14:0] MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_771_nl;
  wire[8:0] nl_MultLoop_acc_771_nl;
  wire[14:0] MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_770_nl;
  wire[8:0] nl_MultLoop_acc_770_nl;
  wire[14:0] MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_769_nl;
  wire[8:0] nl_MultLoop_acc_769_nl;
  wire[14:0] MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_768_nl;
  wire[8:0] nl_MultLoop_acc_768_nl;
  wire[14:0] MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_779_nl;
  wire[8:0] nl_MultLoop_acc_779_nl;
  wire[14:0] MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_778_nl;
  wire[8:0] nl_MultLoop_acc_778_nl;
  wire[14:0] MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_777_nl;
  wire[8:0] nl_MultLoop_acc_777_nl;
  wire[14:0] MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_776_nl;
  wire[8:0] nl_MultLoop_acc_776_nl;
  wire[14:0] MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_775_nl;
  wire[8:0] nl_MultLoop_acc_775_nl;
  wire[14:0] MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_774_nl;
  wire[8:0] nl_MultLoop_acc_774_nl;
  wire[14:0] MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_773_nl;
  wire[8:0] nl_MultLoop_acc_773_nl;
  wire[14:0] MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_772_nl;
  wire[8:0] nl_MultLoop_acc_772_nl;
  wire[14:0] MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_795_nl;
  wire[8:0] nl_MultLoop_acc_795_nl;
  wire[14:0] MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_794_nl;
  wire[8:0] nl_MultLoop_acc_794_nl;
  wire[14:0] MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_793_nl;
  wire[8:0] nl_MultLoop_acc_793_nl;
  wire[14:0] MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_792_nl;
  wire[8:0] nl_MultLoop_acc_792_nl;
  wire[14:0] MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_789_nl;
  wire[8:0] nl_MultLoop_acc_789_nl;
  wire[14:0] MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_788_nl;
  wire[8:0] nl_MultLoop_acc_788_nl;
  wire[14:0] MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_785_nl;
  wire[8:0] nl_MultLoop_acc_785_nl;
  wire[14:0] MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_784_nl;
  wire[8:0] nl_MultLoop_acc_784_nl;
  wire[14:0] MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_781_nl;
  wire[8:0] nl_MultLoop_acc_781_nl;
  wire[14:0] MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_780_nl;
  wire[8:0] nl_MultLoop_acc_780_nl;
  wire[14:0] MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_765_nl;
  wire[8:0] nl_MultLoop_acc_765_nl;
  wire[14:0] MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_764_nl;
  wire[8:0] nl_MultLoop_acc_764_nl;
  wire[14:0] MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_381_nl;
  wire[8:0] nl_MultLoop_acc_381_nl;
  wire[7:0] MultLoop_acc_379_nl;
  wire[8:0] nl_MultLoop_acc_379_nl;
  wire[7:0] MultLoop_acc_375_nl;
  wire[8:0] nl_MultLoop_acc_375_nl;
  wire[7:0] MultLoop_acc_367_nl;
  wire[8:0] nl_MultLoop_acc_367_nl;
  wire[7:0] MultLoop_acc_351_nl;
  wire[8:0] nl_MultLoop_acc_351_nl;
  wire[7:0] MultLoop_acc_319_nl;
  wire[8:0] nl_MultLoop_acc_319_nl;
  wire[7:0] MultLoop_acc_255_nl;
  wire[8:0] nl_MultLoop_acc_255_nl;
  wire[14:0] MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_318_nl;
  wire[8:0] nl_MultLoop_acc_318_nl;
  wire[14:0] MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_350_nl;
  wire[8:0] nl_MultLoop_acc_350_nl;
  wire[7:0] MultLoop_acc_317_nl;
  wire[8:0] nl_MultLoop_acc_317_nl;
  wire[14:0] MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_316_nl;
  wire[8:0] nl_MultLoop_acc_316_nl;
  wire[14:0] MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_366_nl;
  wire[9:0] nl_MultLoop_acc_366_nl;
  wire[7:0] MultLoop_acc_315_nl;
  wire[8:0] nl_MultLoop_acc_315_nl;
  wire[14:0] MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_314_nl;
  wire[8:0] nl_MultLoop_acc_314_nl;
  wire[14:0] MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_313_nl;
  wire[8:0] nl_MultLoop_acc_313_nl;
  wire[14:0] MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_312_nl;
  wire[8:0] nl_MultLoop_acc_312_nl;
  wire[14:0] MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_374_nl;
  wire[10:0] nl_MultLoop_acc_374_nl;
  wire[7:0] MultLoop_acc_307_nl;
  wire[8:0] nl_MultLoop_acc_307_nl;
  wire[14:0] MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_306_nl;
  wire[8:0] nl_MultLoop_acc_306_nl;
  wire[14:0] MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_311_nl;
  wire[8:0] nl_MultLoop_acc_311_nl;
  wire[14:0] MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_310_nl;
  wire[8:0] nl_MultLoop_acc_310_nl;
  wire[14:0] MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_309_nl;
  wire[8:0] nl_MultLoop_acc_309_nl;
  wire[14:0] MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_308_nl;
  wire[8:0] nl_MultLoop_acc_308_nl;
  wire[14:0] MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_305_nl;
  wire[8:0] nl_MultLoop_acc_305_nl;
  wire[14:0] MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_304_nl;
  wire[8:0] nl_MultLoop_acc_304_nl;
  wire[14:0] MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_378_nl;
  wire[11:0] nl_MultLoop_acc_378_nl;
  wire[7:0] MultLoop_acc_303_nl;
  wire[8:0] nl_MultLoop_acc_303_nl;
  wire[14:0] MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_302_nl;
  wire[8:0] nl_MultLoop_acc_302_nl;
  wire[14:0] MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_301_nl;
  wire[8:0] nl_MultLoop_acc_301_nl;
  wire[14:0] MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_300_nl;
  wire[8:0] nl_MultLoop_acc_300_nl;
  wire[14:0] MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_299_nl;
  wire[8:0] nl_MultLoop_acc_299_nl;
  wire[14:0] MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_298_nl;
  wire[8:0] nl_MultLoop_acc_298_nl;
  wire[14:0] MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_297_nl;
  wire[8:0] nl_MultLoop_acc_297_nl;
  wire[14:0] MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_296_nl;
  wire[8:0] nl_MultLoop_acc_296_nl;
  wire[14:0] MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_291_nl;
  wire[8:0] nl_MultLoop_acc_291_nl;
  wire[14:0] MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_290_nl;
  wire[8:0] nl_MultLoop_acc_290_nl;
  wire[14:0] MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_289_nl;
  wire[8:0] nl_MultLoop_acc_289_nl;
  wire[14:0] MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_288_nl;
  wire[8:0] nl_MultLoop_acc_288_nl;
  wire[14:0] MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_295_nl;
  wire[8:0] nl_MultLoop_acc_295_nl;
  wire[14:0] MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_294_nl;
  wire[8:0] nl_MultLoop_acc_294_nl;
  wire[14:0] MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_293_nl;
  wire[8:0] nl_MultLoop_acc_293_nl;
  wire[14:0] MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_292_nl;
  wire[8:0] nl_MultLoop_acc_292_nl;
  wire[14:0] MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_380_nl;
  wire[12:0] nl_MultLoop_acc_380_nl;
  wire[7:0] MultLoop_acc_283_nl;
  wire[8:0] nl_MultLoop_acc_283_nl;
  wire[14:0] MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_282_nl;
  wire[8:0] nl_MultLoop_acc_282_nl;
  wire[14:0] MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_275_nl;
  wire[8:0] nl_MultLoop_acc_275_nl;
  wire[14:0] MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_274_nl;
  wire[8:0] nl_MultLoop_acc_274_nl;
  wire[14:0] MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_279_nl;
  wire[8:0] nl_MultLoop_acc_279_nl;
  wire[14:0] MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_278_nl;
  wire[8:0] nl_MultLoop_acc_278_nl;
  wire[14:0] MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_259_nl;
  wire[8:0] nl_MultLoop_acc_259_nl;
  wire[14:0] MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_258_nl;
  wire[8:0] nl_MultLoop_acc_258_nl;
  wire[14:0] MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_263_nl;
  wire[8:0] nl_MultLoop_acc_263_nl;
  wire[14:0] MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_262_nl;
  wire[8:0] nl_MultLoop_acc_262_nl;
  wire[14:0] MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_261_nl;
  wire[8:0] nl_MultLoop_acc_261_nl;
  wire[14:0] MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_260_nl;
  wire[8:0] nl_MultLoop_acc_260_nl;
  wire[14:0] MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_271_nl;
  wire[8:0] nl_MultLoop_acc_271_nl;
  wire[14:0] MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_270_nl;
  wire[8:0] nl_MultLoop_acc_270_nl;
  wire[14:0] MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_269_nl;
  wire[8:0] nl_MultLoop_acc_269_nl;
  wire[14:0] MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_268_nl;
  wire[8:0] nl_MultLoop_acc_268_nl;
  wire[14:0] MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_267_nl;
  wire[8:0] nl_MultLoop_acc_267_nl;
  wire[14:0] MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_266_nl;
  wire[8:0] nl_MultLoop_acc_266_nl;
  wire[14:0] MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_265_nl;
  wire[8:0] nl_MultLoop_acc_265_nl;
  wire[14:0] MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_264_nl;
  wire[8:0] nl_MultLoop_acc_264_nl;
  wire[14:0] MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_287_nl;
  wire[8:0] nl_MultLoop_acc_287_nl;
  wire[14:0] MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_286_nl;
  wire[8:0] nl_MultLoop_acc_286_nl;
  wire[14:0] MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_285_nl;
  wire[8:0] nl_MultLoop_acc_285_nl;
  wire[14:0] MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_284_nl;
  wire[8:0] nl_MultLoop_acc_284_nl;
  wire[14:0] MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_281_nl;
  wire[8:0] nl_MultLoop_acc_281_nl;
  wire[14:0] MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_280_nl;
  wire[8:0] nl_MultLoop_acc_280_nl;
  wire[14:0] MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_277_nl;
  wire[8:0] nl_MultLoop_acc_277_nl;
  wire[14:0] MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_276_nl;
  wire[8:0] nl_MultLoop_acc_276_nl;
  wire[14:0] MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_273_nl;
  wire[8:0] nl_MultLoop_acc_273_nl;
  wire[14:0] MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_272_nl;
  wire[8:0] nl_MultLoop_acc_272_nl;
  wire[14:0] MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_257_nl;
  wire[8:0] nl_MultLoop_acc_257_nl;
  wire[14:0] MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_256_nl;
  wire[8:0] nl_MultLoop_acc_256_nl;
  wire[14:0] MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_762_nl;
  wire[8:0] nl_MultLoop_acc_762_nl;
  wire[7:0] MultLoop_acc_760_nl;
  wire[8:0] nl_MultLoop_acc_760_nl;
  wire[7:0] MultLoop_acc_756_nl;
  wire[8:0] nl_MultLoop_acc_756_nl;
  wire[7:0] MultLoop_acc_748_nl;
  wire[8:0] nl_MultLoop_acc_748_nl;
  wire[7:0] MultLoop_acc_732_nl;
  wire[8:0] nl_MultLoop_acc_732_nl;
  wire[7:0] MultLoop_acc_700_nl;
  wire[8:0] nl_MultLoop_acc_700_nl;
  wire[7:0] MultLoop_acc_636_nl;
  wire[8:0] nl_MultLoop_acc_636_nl;
  wire[14:0] MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_699_nl;
  wire[8:0] nl_MultLoop_acc_699_nl;
  wire[14:0] MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_731_nl;
  wire[8:0] nl_MultLoop_acc_731_nl;
  wire[7:0] MultLoop_acc_698_nl;
  wire[8:0] nl_MultLoop_acc_698_nl;
  wire[14:0] MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_697_nl;
  wire[8:0] nl_MultLoop_acc_697_nl;
  wire[14:0] MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_747_nl;
  wire[9:0] nl_MultLoop_acc_747_nl;
  wire[7:0] MultLoop_acc_696_nl;
  wire[8:0] nl_MultLoop_acc_696_nl;
  wire[14:0] MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_695_nl;
  wire[8:0] nl_MultLoop_acc_695_nl;
  wire[14:0] MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_694_nl;
  wire[8:0] nl_MultLoop_acc_694_nl;
  wire[14:0] MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_693_nl;
  wire[8:0] nl_MultLoop_acc_693_nl;
  wire[14:0] MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_755_nl;
  wire[10:0] nl_MultLoop_acc_755_nl;
  wire[7:0] MultLoop_acc_688_nl;
  wire[8:0] nl_MultLoop_acc_688_nl;
  wire[14:0] MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_687_nl;
  wire[8:0] nl_MultLoop_acc_687_nl;
  wire[14:0] MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_692_nl;
  wire[8:0] nl_MultLoop_acc_692_nl;
  wire[14:0] MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_691_nl;
  wire[8:0] nl_MultLoop_acc_691_nl;
  wire[14:0] MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_690_nl;
  wire[8:0] nl_MultLoop_acc_690_nl;
  wire[14:0] MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_689_nl;
  wire[8:0] nl_MultLoop_acc_689_nl;
  wire[14:0] MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_686_nl;
  wire[8:0] nl_MultLoop_acc_686_nl;
  wire[14:0] MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_685_nl;
  wire[8:0] nl_MultLoop_acc_685_nl;
  wire[14:0] MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_759_nl;
  wire[11:0] nl_MultLoop_acc_759_nl;
  wire[7:0] MultLoop_acc_684_nl;
  wire[8:0] nl_MultLoop_acc_684_nl;
  wire[14:0] MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_683_nl;
  wire[8:0] nl_MultLoop_acc_683_nl;
  wire[14:0] MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_682_nl;
  wire[8:0] nl_MultLoop_acc_682_nl;
  wire[14:0] MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_681_nl;
  wire[8:0] nl_MultLoop_acc_681_nl;
  wire[14:0] MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_680_nl;
  wire[8:0] nl_MultLoop_acc_680_nl;
  wire[14:0] MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_679_nl;
  wire[8:0] nl_MultLoop_acc_679_nl;
  wire[14:0] MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_678_nl;
  wire[8:0] nl_MultLoop_acc_678_nl;
  wire[14:0] MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_677_nl;
  wire[8:0] nl_MultLoop_acc_677_nl;
  wire[14:0] MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_672_nl;
  wire[8:0] nl_MultLoop_acc_672_nl;
  wire[14:0] MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_671_nl;
  wire[8:0] nl_MultLoop_acc_671_nl;
  wire[14:0] MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_670_nl;
  wire[8:0] nl_MultLoop_acc_670_nl;
  wire[14:0] MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_669_nl;
  wire[8:0] nl_MultLoop_acc_669_nl;
  wire[14:0] MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_676_nl;
  wire[8:0] nl_MultLoop_acc_676_nl;
  wire[14:0] MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_675_nl;
  wire[8:0] nl_MultLoop_acc_675_nl;
  wire[14:0] MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_674_nl;
  wire[8:0] nl_MultLoop_acc_674_nl;
  wire[14:0] MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_673_nl;
  wire[8:0] nl_MultLoop_acc_673_nl;
  wire[14:0] MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_761_nl;
  wire[12:0] nl_MultLoop_acc_761_nl;
  wire[7:0] MultLoop_acc_664_nl;
  wire[8:0] nl_MultLoop_acc_664_nl;
  wire[14:0] MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_663_nl;
  wire[8:0] nl_MultLoop_acc_663_nl;
  wire[14:0] MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_656_nl;
  wire[8:0] nl_MultLoop_acc_656_nl;
  wire[14:0] MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_655_nl;
  wire[8:0] nl_MultLoop_acc_655_nl;
  wire[14:0] MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_660_nl;
  wire[8:0] nl_MultLoop_acc_660_nl;
  wire[14:0] MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_659_nl;
  wire[8:0] nl_MultLoop_acc_659_nl;
  wire[14:0] MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_640_nl;
  wire[8:0] nl_MultLoop_acc_640_nl;
  wire[14:0] MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_639_nl;
  wire[8:0] nl_MultLoop_acc_639_nl;
  wire[14:0] MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_644_nl;
  wire[8:0] nl_MultLoop_acc_644_nl;
  wire[14:0] MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_643_nl;
  wire[8:0] nl_MultLoop_acc_643_nl;
  wire[14:0] MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_642_nl;
  wire[8:0] nl_MultLoop_acc_642_nl;
  wire[14:0] MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_641_nl;
  wire[8:0] nl_MultLoop_acc_641_nl;
  wire[14:0] MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_652_nl;
  wire[8:0] nl_MultLoop_acc_652_nl;
  wire[14:0] MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_651_nl;
  wire[8:0] nl_MultLoop_acc_651_nl;
  wire[14:0] MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_650_nl;
  wire[8:0] nl_MultLoop_acc_650_nl;
  wire[14:0] MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_649_nl;
  wire[8:0] nl_MultLoop_acc_649_nl;
  wire[14:0] MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_648_nl;
  wire[8:0] nl_MultLoop_acc_648_nl;
  wire[14:0] MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_647_nl;
  wire[8:0] nl_MultLoop_acc_647_nl;
  wire[14:0] MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_646_nl;
  wire[8:0] nl_MultLoop_acc_646_nl;
  wire[14:0] MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_645_nl;
  wire[8:0] nl_MultLoop_acc_645_nl;
  wire[14:0] MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_668_nl;
  wire[8:0] nl_MultLoop_acc_668_nl;
  wire[14:0] MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_667_nl;
  wire[8:0] nl_MultLoop_acc_667_nl;
  wire[14:0] MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_666_nl;
  wire[8:0] nl_MultLoop_acc_666_nl;
  wire[14:0] MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_665_nl;
  wire[8:0] nl_MultLoop_acc_665_nl;
  wire[14:0] MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_662_nl;
  wire[8:0] nl_MultLoop_acc_662_nl;
  wire[14:0] MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_661_nl;
  wire[8:0] nl_MultLoop_acc_661_nl;
  wire[14:0] MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_658_nl;
  wire[8:0] nl_MultLoop_acc_658_nl;
  wire[14:0] MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_657_nl;
  wire[8:0] nl_MultLoop_acc_657_nl;
  wire[14:0] MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_654_nl;
  wire[8:0] nl_MultLoop_acc_654_nl;
  wire[14:0] MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_653_nl;
  wire[8:0] nl_MultLoop_acc_653_nl;
  wire[14:0] MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_638_nl;
  wire[8:0] nl_MultLoop_acc_638_nl;
  wire[14:0] MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_637_nl;
  wire[8:0] nl_MultLoop_acc_637_nl;
  wire[14:0] MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_508_nl;
  wire[8:0] nl_MultLoop_acc_508_nl;
  wire[7:0] MultLoop_acc_506_nl;
  wire[8:0] nl_MultLoop_acc_506_nl;
  wire[7:0] MultLoop_acc_502_nl;
  wire[8:0] nl_MultLoop_acc_502_nl;
  wire[7:0] MultLoop_acc_494_nl;
  wire[8:0] nl_MultLoop_acc_494_nl;
  wire[7:0] MultLoop_acc_478_nl;
  wire[8:0] nl_MultLoop_acc_478_nl;
  wire[7:0] MultLoop_acc_446_nl;
  wire[8:0] nl_MultLoop_acc_446_nl;
  wire[7:0] MultLoop_acc_382_nl;
  wire[8:0] nl_MultLoop_acc_382_nl;
  wire[14:0] MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_445_nl;
  wire[8:0] nl_MultLoop_acc_445_nl;
  wire[14:0] MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_477_nl;
  wire[8:0] nl_MultLoop_acc_477_nl;
  wire[7:0] MultLoop_acc_444_nl;
  wire[8:0] nl_MultLoop_acc_444_nl;
  wire[14:0] MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_443_nl;
  wire[8:0] nl_MultLoop_acc_443_nl;
  wire[14:0] MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_493_nl;
  wire[9:0] nl_MultLoop_acc_493_nl;
  wire[7:0] MultLoop_acc_442_nl;
  wire[8:0] nl_MultLoop_acc_442_nl;
  wire[14:0] MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_441_nl;
  wire[8:0] nl_MultLoop_acc_441_nl;
  wire[14:0] MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_440_nl;
  wire[8:0] nl_MultLoop_acc_440_nl;
  wire[14:0] MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_439_nl;
  wire[8:0] nl_MultLoop_acc_439_nl;
  wire[14:0] MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_501_nl;
  wire[10:0] nl_MultLoop_acc_501_nl;
  wire[7:0] MultLoop_acc_434_nl;
  wire[8:0] nl_MultLoop_acc_434_nl;
  wire[14:0] MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_433_nl;
  wire[8:0] nl_MultLoop_acc_433_nl;
  wire[14:0] MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_438_nl;
  wire[8:0] nl_MultLoop_acc_438_nl;
  wire[14:0] MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_437_nl;
  wire[8:0] nl_MultLoop_acc_437_nl;
  wire[14:0] MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_436_nl;
  wire[8:0] nl_MultLoop_acc_436_nl;
  wire[14:0] MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_435_nl;
  wire[8:0] nl_MultLoop_acc_435_nl;
  wire[14:0] MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_432_nl;
  wire[8:0] nl_MultLoop_acc_432_nl;
  wire[14:0] MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_431_nl;
  wire[8:0] nl_MultLoop_acc_431_nl;
  wire[14:0] MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_505_nl;
  wire[11:0] nl_MultLoop_acc_505_nl;
  wire[7:0] MultLoop_acc_430_nl;
  wire[8:0] nl_MultLoop_acc_430_nl;
  wire[14:0] MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_429_nl;
  wire[8:0] nl_MultLoop_acc_429_nl;
  wire[14:0] MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_428_nl;
  wire[8:0] nl_MultLoop_acc_428_nl;
  wire[14:0] MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_427_nl;
  wire[8:0] nl_MultLoop_acc_427_nl;
  wire[14:0] MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_426_nl;
  wire[8:0] nl_MultLoop_acc_426_nl;
  wire[14:0] MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_425_nl;
  wire[8:0] nl_MultLoop_acc_425_nl;
  wire[14:0] MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_424_nl;
  wire[8:0] nl_MultLoop_acc_424_nl;
  wire[14:0] MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_423_nl;
  wire[8:0] nl_MultLoop_acc_423_nl;
  wire[14:0] MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_418_nl;
  wire[8:0] nl_MultLoop_acc_418_nl;
  wire[14:0] MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_417_nl;
  wire[8:0] nl_MultLoop_acc_417_nl;
  wire[14:0] MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_416_nl;
  wire[8:0] nl_MultLoop_acc_416_nl;
  wire[14:0] MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_415_nl;
  wire[8:0] nl_MultLoop_acc_415_nl;
  wire[14:0] MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_422_nl;
  wire[8:0] nl_MultLoop_acc_422_nl;
  wire[14:0] MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_421_nl;
  wire[8:0] nl_MultLoop_acc_421_nl;
  wire[14:0] MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_420_nl;
  wire[8:0] nl_MultLoop_acc_420_nl;
  wire[14:0] MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_419_nl;
  wire[8:0] nl_MultLoop_acc_419_nl;
  wire[14:0] MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_507_nl;
  wire[12:0] nl_MultLoop_acc_507_nl;
  wire[7:0] MultLoop_acc_410_nl;
  wire[8:0] nl_MultLoop_acc_410_nl;
  wire[14:0] MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_409_nl;
  wire[8:0] nl_MultLoop_acc_409_nl;
  wire[14:0] MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_402_nl;
  wire[8:0] nl_MultLoop_acc_402_nl;
  wire[14:0] MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_401_nl;
  wire[8:0] nl_MultLoop_acc_401_nl;
  wire[14:0] MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_406_nl;
  wire[8:0] nl_MultLoop_acc_406_nl;
  wire[14:0] MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_405_nl;
  wire[8:0] nl_MultLoop_acc_405_nl;
  wire[14:0] MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_386_nl;
  wire[8:0] nl_MultLoop_acc_386_nl;
  wire[14:0] MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_385_nl;
  wire[8:0] nl_MultLoop_acc_385_nl;
  wire[14:0] MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_390_nl;
  wire[8:0] nl_MultLoop_acc_390_nl;
  wire[14:0] MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_389_nl;
  wire[8:0] nl_MultLoop_acc_389_nl;
  wire[14:0] MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_388_nl;
  wire[8:0] nl_MultLoop_acc_388_nl;
  wire[14:0] MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_387_nl;
  wire[8:0] nl_MultLoop_acc_387_nl;
  wire[14:0] MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_398_nl;
  wire[8:0] nl_MultLoop_acc_398_nl;
  wire[14:0] MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_397_nl;
  wire[8:0] nl_MultLoop_acc_397_nl;
  wire[14:0] MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_396_nl;
  wire[8:0] nl_MultLoop_acc_396_nl;
  wire[14:0] MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_395_nl;
  wire[8:0] nl_MultLoop_acc_395_nl;
  wire[14:0] MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_394_nl;
  wire[8:0] nl_MultLoop_acc_394_nl;
  wire[14:0] MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_393_nl;
  wire[8:0] nl_MultLoop_acc_393_nl;
  wire[14:0] MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_392_nl;
  wire[8:0] nl_MultLoop_acc_392_nl;
  wire[14:0] MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_391_nl;
  wire[8:0] nl_MultLoop_acc_391_nl;
  wire[14:0] MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_414_nl;
  wire[8:0] nl_MultLoop_acc_414_nl;
  wire[14:0] MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_413_nl;
  wire[8:0] nl_MultLoop_acc_413_nl;
  wire[14:0] MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_412_nl;
  wire[8:0] nl_MultLoop_acc_412_nl;
  wire[14:0] MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_411_nl;
  wire[8:0] nl_MultLoop_acc_411_nl;
  wire[14:0] MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_408_nl;
  wire[8:0] nl_MultLoop_acc_408_nl;
  wire[14:0] MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_407_nl;
  wire[8:0] nl_MultLoop_acc_407_nl;
  wire[14:0] MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_404_nl;
  wire[8:0] nl_MultLoop_acc_404_nl;
  wire[14:0] MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_403_nl;
  wire[8:0] nl_MultLoop_acc_403_nl;
  wire[14:0] MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_400_nl;
  wire[8:0] nl_MultLoop_acc_400_nl;
  wire[14:0] MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_399_nl;
  wire[8:0] nl_MultLoop_acc_399_nl;
  wire[14:0] MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_384_nl;
  wire[8:0] nl_MultLoop_acc_384_nl;
  wire[14:0] MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_383_nl;
  wire[8:0] nl_MultLoop_acc_383_nl;
  wire[14:0] MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_635_nl;
  wire[8:0] nl_MultLoop_acc_635_nl;
  wire[7:0] MultLoop_acc_633_nl;
  wire[8:0] nl_MultLoop_acc_633_nl;
  wire[7:0] MultLoop_acc_629_nl;
  wire[8:0] nl_MultLoop_acc_629_nl;
  wire[7:0] MultLoop_acc_621_nl;
  wire[8:0] nl_MultLoop_acc_621_nl;
  wire[7:0] MultLoop_acc_605_nl;
  wire[8:0] nl_MultLoop_acc_605_nl;
  wire[7:0] MultLoop_acc_573_nl;
  wire[8:0] nl_MultLoop_acc_573_nl;
  wire[7:0] MultLoop_acc_509_nl;
  wire[8:0] nl_MultLoop_acc_509_nl;
  wire[14:0] MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_572_nl;
  wire[8:0] nl_MultLoop_acc_572_nl;
  wire[14:0] MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_604_nl;
  wire[8:0] nl_MultLoop_acc_604_nl;
  wire[7:0] MultLoop_acc_571_nl;
  wire[8:0] nl_MultLoop_acc_571_nl;
  wire[14:0] MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_570_nl;
  wire[8:0] nl_MultLoop_acc_570_nl;
  wire[14:0] MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_620_nl;
  wire[9:0] nl_MultLoop_acc_620_nl;
  wire[7:0] MultLoop_acc_569_nl;
  wire[8:0] nl_MultLoop_acc_569_nl;
  wire[14:0] MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_568_nl;
  wire[8:0] nl_MultLoop_acc_568_nl;
  wire[14:0] MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_567_nl;
  wire[8:0] nl_MultLoop_acc_567_nl;
  wire[14:0] MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_566_nl;
  wire[8:0] nl_MultLoop_acc_566_nl;
  wire[14:0] MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_628_nl;
  wire[10:0] nl_MultLoop_acc_628_nl;
  wire[7:0] MultLoop_acc_561_nl;
  wire[8:0] nl_MultLoop_acc_561_nl;
  wire[14:0] MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_560_nl;
  wire[8:0] nl_MultLoop_acc_560_nl;
  wire[14:0] MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_565_nl;
  wire[8:0] nl_MultLoop_acc_565_nl;
  wire[14:0] MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_564_nl;
  wire[8:0] nl_MultLoop_acc_564_nl;
  wire[14:0] MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_563_nl;
  wire[8:0] nl_MultLoop_acc_563_nl;
  wire[14:0] MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_562_nl;
  wire[8:0] nl_MultLoop_acc_562_nl;
  wire[14:0] MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_559_nl;
  wire[8:0] nl_MultLoop_acc_559_nl;
  wire[14:0] MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_558_nl;
  wire[8:0] nl_MultLoop_acc_558_nl;
  wire[14:0] MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_632_nl;
  wire[11:0] nl_MultLoop_acc_632_nl;
  wire[7:0] MultLoop_acc_557_nl;
  wire[8:0] nl_MultLoop_acc_557_nl;
  wire[14:0] MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_556_nl;
  wire[8:0] nl_MultLoop_acc_556_nl;
  wire[14:0] MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_555_nl;
  wire[8:0] nl_MultLoop_acc_555_nl;
  wire[14:0] MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_554_nl;
  wire[8:0] nl_MultLoop_acc_554_nl;
  wire[14:0] MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_553_nl;
  wire[8:0] nl_MultLoop_acc_553_nl;
  wire[14:0] MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_552_nl;
  wire[8:0] nl_MultLoop_acc_552_nl;
  wire[14:0] MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_551_nl;
  wire[8:0] nl_MultLoop_acc_551_nl;
  wire[14:0] MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_550_nl;
  wire[8:0] nl_MultLoop_acc_550_nl;
  wire[14:0] MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_545_nl;
  wire[8:0] nl_MultLoop_acc_545_nl;
  wire[14:0] MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_544_nl;
  wire[8:0] nl_MultLoop_acc_544_nl;
  wire[14:0] MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_543_nl;
  wire[8:0] nl_MultLoop_acc_543_nl;
  wire[14:0] MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_542_nl;
  wire[8:0] nl_MultLoop_acc_542_nl;
  wire[14:0] MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_549_nl;
  wire[8:0] nl_MultLoop_acc_549_nl;
  wire[14:0] MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_548_nl;
  wire[8:0] nl_MultLoop_acc_548_nl;
  wire[14:0] MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_547_nl;
  wire[8:0] nl_MultLoop_acc_547_nl;
  wire[14:0] MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_546_nl;
  wire[8:0] nl_MultLoop_acc_546_nl;
  wire[14:0] MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_634_nl;
  wire[12:0] nl_MultLoop_acc_634_nl;
  wire[7:0] MultLoop_acc_537_nl;
  wire[8:0] nl_MultLoop_acc_537_nl;
  wire[14:0] MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_536_nl;
  wire[8:0] nl_MultLoop_acc_536_nl;
  wire[14:0] MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_529_nl;
  wire[8:0] nl_MultLoop_acc_529_nl;
  wire[14:0] MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_528_nl;
  wire[8:0] nl_MultLoop_acc_528_nl;
  wire[14:0] MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_533_nl;
  wire[8:0] nl_MultLoop_acc_533_nl;
  wire[14:0] MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_532_nl;
  wire[8:0] nl_MultLoop_acc_532_nl;
  wire[14:0] MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_513_nl;
  wire[8:0] nl_MultLoop_acc_513_nl;
  wire[14:0] MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_512_nl;
  wire[8:0] nl_MultLoop_acc_512_nl;
  wire[14:0] MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_517_nl;
  wire[8:0] nl_MultLoop_acc_517_nl;
  wire[14:0] MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_516_nl;
  wire[8:0] nl_MultLoop_acc_516_nl;
  wire[14:0] MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_515_nl;
  wire[8:0] nl_MultLoop_acc_515_nl;
  wire[14:0] MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_514_nl;
  wire[8:0] nl_MultLoop_acc_514_nl;
  wire[14:0] MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_525_nl;
  wire[8:0] nl_MultLoop_acc_525_nl;
  wire[14:0] MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_524_nl;
  wire[8:0] nl_MultLoop_acc_524_nl;
  wire[14:0] MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_523_nl;
  wire[8:0] nl_MultLoop_acc_523_nl;
  wire[14:0] MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_522_nl;
  wire[8:0] nl_MultLoop_acc_522_nl;
  wire[14:0] MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_521_nl;
  wire[8:0] nl_MultLoop_acc_521_nl;
  wire[14:0] MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_520_nl;
  wire[8:0] nl_MultLoop_acc_520_nl;
  wire[14:0] MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_519_nl;
  wire[8:0] nl_MultLoop_acc_519_nl;
  wire[14:0] MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_518_nl;
  wire[8:0] nl_MultLoop_acc_518_nl;
  wire[14:0] MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_541_nl;
  wire[8:0] nl_MultLoop_acc_541_nl;
  wire[14:0] MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_540_nl;
  wire[8:0] nl_MultLoop_acc_540_nl;
  wire[14:0] MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_539_nl;
  wire[8:0] nl_MultLoop_acc_539_nl;
  wire[14:0] MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_538_nl;
  wire[8:0] nl_MultLoop_acc_538_nl;
  wire[14:0] MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_535_nl;
  wire[8:0] nl_MultLoop_acc_535_nl;
  wire[14:0] MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_534_nl;
  wire[8:0] nl_MultLoop_acc_534_nl;
  wire[14:0] MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_531_nl;
  wire[8:0] nl_MultLoop_acc_531_nl;
  wire[14:0] MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_530_nl;
  wire[8:0] nl_MultLoop_acc_530_nl;
  wire[14:0] MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_527_nl;
  wire[8:0] nl_MultLoop_acc_527_nl;
  wire[14:0] MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_526_nl;
  wire[8:0] nl_MultLoop_acc_526_nl;
  wire[14:0] MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_511_nl;
  wire[8:0] nl_MultLoop_acc_511_nl;
  wire[14:0] MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[7:0] MultLoop_acc_510_nl;
  wire[8:0] nl_MultLoop_acc_510_nl;
  wire[14:0] MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[14:0] MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [15:0] nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] AccumDotWidth_acc_2262_nl;
  wire[8:0] nl_AccumDotWidth_acc_2262_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2251_nl;
  wire[8:0] nl_AccumDotWidth_acc_2251_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2240_nl;
  wire[8:0] nl_AccumDotWidth_acc_2240_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2229_nl;
  wire[8:0] nl_AccumDotWidth_acc_2229_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2218_nl;
  wire[8:0] nl_AccumDotWidth_acc_2218_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2207_nl;
  wire[8:0] nl_AccumDotWidth_acc_2207_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2196_nl;
  wire[8:0] nl_AccumDotWidth_acc_2196_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2185_nl;
  wire[8:0] nl_AccumDotWidth_acc_2185_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2168_nl;
  wire[8:0] nl_AccumDotWidth_acc_2168_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2151_nl;
  wire[8:0] nl_AccumDotWidth_acc_2151_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2134_nl;
  wire[8:0] nl_AccumDotWidth_acc_2134_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2117_nl;
  wire[8:0] nl_AccumDotWidth_acc_2117_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2100_nl;
  wire[8:0] nl_AccumDotWidth_acc_2100_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2083_nl;
  wire[8:0] nl_AccumDotWidth_acc_2083_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2066_nl;
  wire[8:0] nl_AccumDotWidth_acc_2066_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2049_nl;
  wire[8:0] nl_AccumDotWidth_acc_2049_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2032_nl;
  wire[8:0] nl_AccumDotWidth_acc_2032_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_2015_nl;
  wire[8:0] nl_AccumDotWidth_acc_2015_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1998_nl;
  wire[8:0] nl_AccumDotWidth_acc_1998_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1981_nl;
  wire[8:0] nl_AccumDotWidth_acc_1981_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1964_nl;
  wire[8:0] nl_AccumDotWidth_acc_1964_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1947_nl;
  wire[8:0] nl_AccumDotWidth_acc_1947_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1930_nl;
  wire[8:0] nl_AccumDotWidth_acc_1930_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1913_nl;
  wire[8:0] nl_AccumDotWidth_acc_1913_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1902_nl;
  wire[8:0] nl_AccumDotWidth_acc_1902_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1891_nl;
  wire[8:0] nl_AccumDotWidth_acc_1891_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1880_nl;
  wire[8:0] nl_AccumDotWidth_acc_1880_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1869_nl;
  wire[8:0] nl_AccumDotWidth_acc_1869_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1858_nl;
  wire[8:0] nl_AccumDotWidth_acc_1858_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1847_nl;
  wire[8:0] nl_AccumDotWidth_acc_1847_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1836_nl;
  wire[8:0] nl_AccumDotWidth_acc_1836_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1825_nl;
  wire[8:0] nl_AccumDotWidth_acc_1825_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1808_nl;
  wire[8:0] nl_AccumDotWidth_acc_1808_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1791_nl;
  wire[8:0] nl_AccumDotWidth_acc_1791_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1774_nl;
  wire[8:0] nl_AccumDotWidth_acc_1774_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1757_nl;
  wire[8:0] nl_AccumDotWidth_acc_1757_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1740_nl;
  wire[8:0] nl_AccumDotWidth_acc_1740_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1723_nl;
  wire[8:0] nl_AccumDotWidth_acc_1723_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1706_nl;
  wire[8:0] nl_AccumDotWidth_acc_1706_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1689_nl;
  wire[8:0] nl_AccumDotWidth_acc_1689_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1663_nl;
  wire[8:0] nl_AccumDotWidth_acc_1663_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1637_nl;
  wire[8:0] nl_AccumDotWidth_acc_1637_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1611_nl;
  wire[8:0] nl_AccumDotWidth_acc_1611_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1585_nl;
  wire[8:0] nl_AccumDotWidth_acc_1585_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1559_nl;
  wire[8:0] nl_AccumDotWidth_acc_1559_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1533_nl;
  wire[8:0] nl_AccumDotWidth_acc_1533_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1507_nl;
  wire[8:0] nl_AccumDotWidth_acc_1507_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1481_nl;
  wire[8:0] nl_AccumDotWidth_acc_1481_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1455_nl;
  wire[8:0] nl_AccumDotWidth_acc_1455_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1429_nl;
  wire[8:0] nl_AccumDotWidth_acc_1429_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1403_nl;
  wire[8:0] nl_AccumDotWidth_acc_1403_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1377_nl;
  wire[8:0] nl_AccumDotWidth_acc_1377_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1351_nl;
  wire[8:0] nl_AccumDotWidth_acc_1351_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1325_nl;
  wire[8:0] nl_AccumDotWidth_acc_1325_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1299_nl;
  wire[8:0] nl_AccumDotWidth_acc_1299_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1273_nl;
  wire[8:0] nl_AccumDotWidth_acc_1273_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1256_nl;
  wire[8:0] nl_AccumDotWidth_acc_1256_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1239_nl;
  wire[8:0] nl_AccumDotWidth_acc_1239_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1222_nl;
  wire[8:0] nl_AccumDotWidth_acc_1222_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1205_nl;
  wire[8:0] nl_AccumDotWidth_acc_1205_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1188_nl;
  wire[8:0] nl_AccumDotWidth_acc_1188_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1171_nl;
  wire[8:0] nl_AccumDotWidth_acc_1171_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1154_nl;
  wire[8:0] nl_AccumDotWidth_acc_1154_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1137_nl;
  wire[8:0] nl_AccumDotWidth_acc_1137_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1120_nl;
  wire[8:0] nl_AccumDotWidth_acc_1120_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1103_nl;
  wire[8:0] nl_AccumDotWidth_acc_1103_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1086_nl;
  wire[8:0] nl_AccumDotWidth_acc_1086_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1069_nl;
  wire[8:0] nl_AccumDotWidth_acc_1069_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1052_nl;
  wire[8:0] nl_AccumDotWidth_acc_1052_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1035_nl;
  wire[8:0] nl_AccumDotWidth_acc_1035_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1018_nl;
  wire[8:0] nl_AccumDotWidth_acc_1018_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_1001_nl;
  wire[8:0] nl_AccumDotWidth_acc_1001_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_975_nl;
  wire[8:0] nl_AccumDotWidth_acc_975_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_949_nl;
  wire[8:0] nl_AccumDotWidth_acc_949_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_923_nl;
  wire[8:0] nl_AccumDotWidth_acc_923_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_897_nl;
  wire[8:0] nl_AccumDotWidth_acc_897_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_871_nl;
  wire[8:0] nl_AccumDotWidth_acc_871_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_845_nl;
  wire[8:0] nl_AccumDotWidth_acc_845_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_819_nl;
  wire[8:0] nl_AccumDotWidth_acc_819_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_793_nl;
  wire[8:0] nl_AccumDotWidth_acc_793_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_767_nl;
  wire[8:0] nl_AccumDotWidth_acc_767_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_741_nl;
  wire[8:0] nl_AccumDotWidth_acc_741_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_715_nl;
  wire[8:0] nl_AccumDotWidth_acc_715_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_689_nl;
  wire[8:0] nl_AccumDotWidth_acc_689_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_663_nl;
  wire[8:0] nl_AccumDotWidth_acc_663_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_637_nl;
  wire[8:0] nl_AccumDotWidth_acc_637_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_611_nl;
  wire[8:0] nl_AccumDotWidth_acc_611_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_585_nl;
  wire[8:0] nl_AccumDotWidth_acc_585_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_568_nl;
  wire[8:0] nl_AccumDotWidth_acc_568_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_551_nl;
  wire[8:0] nl_AccumDotWidth_acc_551_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_534_nl;
  wire[8:0] nl_AccumDotWidth_acc_534_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_517_nl;
  wire[8:0] nl_AccumDotWidth_acc_517_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_500_nl;
  wire[8:0] nl_AccumDotWidth_acc_500_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_483_nl;
  wire[8:0] nl_AccumDotWidth_acc_483_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_466_nl;
  wire[8:0] nl_AccumDotWidth_acc_466_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_449_nl;
  wire[8:0] nl_AccumDotWidth_acc_449_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_438_nl;
  wire[8:0] nl_AccumDotWidth_acc_438_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_427_nl;
  wire[8:0] nl_AccumDotWidth_acc_427_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_416_nl;
  wire[8:0] nl_AccumDotWidth_acc_416_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_405_nl;
  wire[8:0] nl_AccumDotWidth_acc_405_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_394_nl;
  wire[8:0] nl_AccumDotWidth_acc_394_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_383_nl;
  wire[8:0] nl_AccumDotWidth_acc_383_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_372_nl;
  wire[8:0] nl_AccumDotWidth_acc_372_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_361_nl;
  wire[8:0] nl_AccumDotWidth_acc_361_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_344_nl;
  wire[8:0] nl_AccumDotWidth_acc_344_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_327_nl;
  wire[8:0] nl_AccumDotWidth_acc_327_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_310_nl;
  wire[8:0] nl_AccumDotWidth_acc_310_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_293_nl;
  wire[8:0] nl_AccumDotWidth_acc_293_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_276_nl;
  wire[8:0] nl_AccumDotWidth_acc_276_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_259_nl;
  wire[8:0] nl_AccumDotWidth_acc_259_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_242_nl;
  wire[8:0] nl_AccumDotWidth_acc_242_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_225_nl;
  wire[8:0] nl_AccumDotWidth_acc_225_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_208_nl;
  wire[8:0] nl_AccumDotWidth_acc_208_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_191_nl;
  wire[8:0] nl_AccumDotWidth_acc_191_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_174_nl;
  wire[8:0] nl_AccumDotWidth_acc_174_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_157_nl;
  wire[8:0] nl_AccumDotWidth_acc_157_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_140_nl;
  wire[8:0] nl_AccumDotWidth_acc_140_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_123_nl;
  wire[8:0] nl_AccumDotWidth_acc_123_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_106_nl;
  wire[8:0] nl_AccumDotWidth_acc_106_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_89_nl;
  wire[8:0] nl_AccumDotWidth_acc_89_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_78_nl;
  wire[8:0] nl_AccumDotWidth_acc_78_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_67_nl;
  wire[8:0] nl_AccumDotWidth_acc_67_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_56_nl;
  wire[8:0] nl_AccumDotWidth_acc_56_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_45_nl;
  wire[8:0] nl_AccumDotWidth_acc_45_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_34_nl;
  wire[8:0] nl_AccumDotWidth_acc_34_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_23_nl;
  wire[8:0] nl_AccumDotWidth_acc_23_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_12_nl;
  wire[8:0] nl_AccumDotWidth_acc_12_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[7:0] AccumDotWidth_acc_7_nl;
  wire[8:0] nl_AccumDotWidth_acc_7_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl;
  wire[14:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire signed [15:0] nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl;
  wire[8:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;
  wire[9:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [79:0] nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat;
  assign nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat = {1'b0 ,
      layer5_out_rsci_idat_78_72 , 1'b0 , layer5_out_rsci_idat_70_64 , 1'b0 , layer5_out_rsci_idat_62_56
      , 1'b0 , layer5_out_rsci_idat_54_48 , 1'b0 , layer5_out_rsci_idat_46_40 , 1'b0
      , layer5_out_rsci_idat_38_32 , 1'b0 , layer5_out_rsci_idat_30_24 , 1'b0 , layer5_out_rsci_idat_22_16
      , 1'b0 , layer5_out_rsci_idat_14_8 , 1'b0 , layer5_out_rsci_idat_6_0};
  econ_4x4_d10_core_input_1_rsci econ_4x4_d10_core_input_1_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_rdy(input_1_rsc_rdy),
      .core_wen(core_wen),
      .input_1_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_layer5_out_rsci econ_4x4_d10_core_layer5_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_rdy(layer5_out_rsc_rdy),
      .core_wen(core_wen),
      .layer5_out_rsci_oswt(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp),
      .layer5_out_rsci_idat(nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat[79:0])
    );
  econ_4x4_d10_core_const_size_in_1_rsci econ_4x4_d10_core_const_size_in_1_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_rdy(const_size_in_1_rsc_rdy),
      .core_wen(core_wen),
      .const_size_in_1_rsci_oswt(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp)
    );
  econ_4x4_d10_core_const_size_out_1_rsci econ_4x4_d10_core_const_size_out_1_rsci_inst
      (
      .clk(clk),
      .rst(rst),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_rdy(const_size_out_1_rsc_rdy),
      .core_wen(core_wen),
      .const_size_out_1_rsci_oswt(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp)
    );
  econ_4x4_d10_core_w2_rsci econ_4x4_d10_core_w2_rsci_inst (
      .clk(clk),
      .rst(rst),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_rdy(w2_rsc_rdy),
      .core_wen(core_wen),
      .w2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b2_rsci econ_4x4_d10_core_b2_rsci_inst (
      .clk(clk),
      .rst(rst),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_rdy(b2_rsc_rdy),
      .core_wen(core_wen),
      .b2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_w4_rsci econ_4x4_d10_core_w4_rsci_inst (
      .clk(clk),
      .rst(rst),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_rdy(w4_rsc_rdy),
      .core_wen(core_wen),
      .w4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b4_rsci econ_4x4_d10_core_b4_rsci_inst (
      .clk(clk),
      .rst(rst),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_rdy(b4_rsc_rdy),
      .core_wen(core_wen),
      .b4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj econ_4x4_d10_core_input_1_rsc_triosy_obj_inst
      (
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj econ_4x4_d10_core_layer5_out_rsc_triosy_obj_inst
      (
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_inst
      (
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_inst
      (
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj econ_4x4_d10_core_w2_rsc_triosy_obj_inst (
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj econ_4x4_d10_core_b2_rsc_triosy_obj_inst (
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj econ_4x4_d10_core_w4_rsc_triosy_obj_inst (
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj econ_4x4_d10_core_b4_rsc_triosy_obj_inst (
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz),
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_staller econ_4x4_d10_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .layer5_out_rsci_wen_comp(layer5_out_rsci_wen_comp),
      .const_size_in_1_rsci_wen_comp(const_size_in_1_rsci_wen_comp),
      .const_size_out_1_rsci_wen_comp(const_size_out_1_rsci_wen_comp),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .b4_rsci_wen_comp(b4_rsci_wen_comp)
    );
  econ_4x4_d10_core_core_fsm econ_4x4_d10_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign nnet_relu_layer4_t_result_t_relu_config5_for_if_and_cse = core_wen & (~
      (fsm_output[0]));
  assign nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1023:1016]));
  assign MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1144_nl = (readslicef_15_8_7(MultLoop_128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[6:0]);
  assign MultLoop_acc_1144_nl = nl_MultLoop_acc_1144_nl[7:0];
  assign nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[7:0]));
  assign MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1208_nl = MultLoop_acc_1144_nl + (readslicef_15_8_7(MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1208_nl = nl_MultLoop_acc_1208_nl[7:0];
  assign nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[15:8]));
  assign MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[23:16]));
  assign MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1207_nl = (readslicef_15_8_7(MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1207_nl = nl_MultLoop_acc_1207_nl[7:0];
  assign nl_MultLoop_acc_1240_nl = MultLoop_acc_1208_nl + MultLoop_acc_1207_nl;
  assign MultLoop_acc_1240_nl = nl_MultLoop_acc_1240_nl[7:0];
  assign nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[31:24]));
  assign MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[39:32]));
  assign MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1206_nl = (readslicef_15_8_7(MultLoop_4_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_5_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1206_nl = nl_MultLoop_acc_1206_nl[7:0];
  assign nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[47:40]));
  assign MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[55:48]));
  assign MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1205_nl = (readslicef_15_8_7(MultLoop_6_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_7_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1205_nl = nl_MultLoop_acc_1205_nl[7:0];
  assign nl_MultLoop_acc_1239_nl = MultLoop_acc_1206_nl + MultLoop_acc_1205_nl;
  assign MultLoop_acc_1239_nl = nl_MultLoop_acc_1239_nl[7:0];
  assign nl_MultLoop_acc_1256_nl = MultLoop_acc_1240_nl + MultLoop_acc_1239_nl;
  assign MultLoop_acc_1256_nl = nl_MultLoop_acc_1256_nl[7:0];
  assign nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[63:56]));
  assign MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[71:64]));
  assign MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1204_nl = (readslicef_15_8_7(MultLoop_8_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_9_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1204_nl = nl_MultLoop_acc_1204_nl[7:0];
  assign nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[79:72]));
  assign MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[87:80]));
  assign MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1203_nl = (readslicef_15_8_7(MultLoop_10_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_11_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1203_nl = nl_MultLoop_acc_1203_nl[7:0];
  assign nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[95:88]));
  assign MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[103:96]));
  assign MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1202_nl = (readslicef_15_8_7(MultLoop_12_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_13_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1202_nl = nl_MultLoop_acc_1202_nl[7:0];
  assign nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[111:104]));
  assign MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[119:112]));
  assign MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1201_nl = (readslicef_15_8_7(MultLoop_14_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_15_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1201_nl = nl_MultLoop_acc_1201_nl[7:0];
  assign nl_MultLoop_acc_1255_nl = MultLoop_acc_1204_nl + MultLoop_acc_1203_nl +
      MultLoop_acc_1202_nl + MultLoop_acc_1201_nl;
  assign MultLoop_acc_1255_nl = nl_MultLoop_acc_1255_nl[7:0];
  assign nl_MultLoop_acc_1264_nl = MultLoop_acc_1256_nl + MultLoop_acc_1255_nl;
  assign MultLoop_acc_1264_nl = nl_MultLoop_acc_1264_nl[7:0];
  assign nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[191:184]));
  assign MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[199:192]));
  assign MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1196_nl = (readslicef_15_8_7(MultLoop_24_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_25_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1196_nl = nl_MultLoop_acc_1196_nl[7:0];
  assign nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[207:200]));
  assign MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[215:208]));
  assign MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1195_nl = (readslicef_15_8_7(MultLoop_26_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_27_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1195_nl = nl_MultLoop_acc_1195_nl[7:0];
  assign nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[127:120]));
  assign MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[135:128]));
  assign MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1200_nl = (readslicef_15_8_7(MultLoop_16_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_17_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1200_nl = nl_MultLoop_acc_1200_nl[7:0];
  assign nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[143:136]));
  assign MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[151:144]));
  assign MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1199_nl = (readslicef_15_8_7(MultLoop_18_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_19_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1199_nl = nl_MultLoop_acc_1199_nl[7:0];
  assign nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[159:152]));
  assign MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[167:160]));
  assign MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1198_nl = (readslicef_15_8_7(MultLoop_20_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_21_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1198_nl = nl_MultLoop_acc_1198_nl[7:0];
  assign nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[175:168]));
  assign MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[183:176]));
  assign MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1197_nl = (readslicef_15_8_7(MultLoop_22_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_23_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1197_nl = nl_MultLoop_acc_1197_nl[7:0];
  assign nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[223:216]));
  assign MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[231:224]));
  assign MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1194_nl = (readslicef_15_8_7(MultLoop_28_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_29_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1194_nl = nl_MultLoop_acc_1194_nl[7:0];
  assign nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[239:232]));
  assign MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[247:240]));
  assign MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1193_nl = (readslicef_15_8_7(MultLoop_30_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_31_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1193_nl = nl_MultLoop_acc_1193_nl[7:0];
  assign nl_MultLoop_acc_1263_nl = MultLoop_acc_1196_nl + MultLoop_acc_1195_nl +
      MultLoop_acc_1200_nl + MultLoop_acc_1199_nl + MultLoop_acc_1198_nl + MultLoop_acc_1197_nl
      + MultLoop_acc_1194_nl + MultLoop_acc_1193_nl;
  assign MultLoop_acc_1263_nl = nl_MultLoop_acc_1263_nl[7:0];
  assign nl_MultLoop_acc_1268_nl = MultLoop_acc_1264_nl + MultLoop_acc_1263_nl;
  assign MultLoop_acc_1268_nl = nl_MultLoop_acc_1268_nl[7:0];
  assign nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[255:248]));
  assign MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[263:256]));
  assign MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1192_nl = (readslicef_15_8_7(MultLoop_32_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_33_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1192_nl = nl_MultLoop_acc_1192_nl[7:0];
  assign nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[271:264]));
  assign MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[279:272]));
  assign MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1191_nl = (readslicef_15_8_7(MultLoop_34_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_35_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1191_nl = nl_MultLoop_acc_1191_nl[7:0];
  assign nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[287:280]));
  assign MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[295:288]));
  assign MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1190_nl = (readslicef_15_8_7(MultLoop_36_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_37_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1190_nl = nl_MultLoop_acc_1190_nl[7:0];
  assign nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[303:296]));
  assign MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[311:304]));
  assign MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1189_nl = (readslicef_15_8_7(MultLoop_38_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_39_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1189_nl = nl_MultLoop_acc_1189_nl[7:0];
  assign nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[319:312]));
  assign MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[327:320]));
  assign MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1188_nl = (readslicef_15_8_7(MultLoop_40_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_41_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1188_nl = nl_MultLoop_acc_1188_nl[7:0];
  assign nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[335:328]));
  assign MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[343:336]));
  assign MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1187_nl = (readslicef_15_8_7(MultLoop_42_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1187_nl = nl_MultLoop_acc_1187_nl[7:0];
  assign nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[351:344]));
  assign MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[359:352]));
  assign MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1186_nl = (readslicef_15_8_7(MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1186_nl = nl_MultLoop_acc_1186_nl[7:0];
  assign nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[367:360]));
  assign MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[375:368]));
  assign MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1185_nl = (readslicef_15_8_7(MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1185_nl = nl_MultLoop_acc_1185_nl[7:0];
  assign nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[447:440]));
  assign MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[455:448]));
  assign MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1180_nl = (readslicef_15_8_7(MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1180_nl = nl_MultLoop_acc_1180_nl[7:0];
  assign nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[463:456]));
  assign MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[471:464]));
  assign MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1179_nl = (readslicef_15_8_7(MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1179_nl = nl_MultLoop_acc_1179_nl[7:0];
  assign nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[479:472]));
  assign MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[487:480]));
  assign MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1178_nl = (readslicef_15_8_7(MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1178_nl = nl_MultLoop_acc_1178_nl[7:0];
  assign nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[495:488]));
  assign MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[503:496]));
  assign MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1177_nl = (readslicef_15_8_7(MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1177_nl = nl_MultLoop_acc_1177_nl[7:0];
  assign nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[383:376]));
  assign MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[391:384]));
  assign MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1184_nl = (readslicef_15_8_7(MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1184_nl = nl_MultLoop_acc_1184_nl[7:0];
  assign nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[399:392]));
  assign MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[407:400]));
  assign MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1183_nl = (readslicef_15_8_7(MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1183_nl = nl_MultLoop_acc_1183_nl[7:0];
  assign nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[415:408]));
  assign MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[423:416]));
  assign MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1182_nl = (readslicef_15_8_7(MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1182_nl = nl_MultLoop_acc_1182_nl[7:0];
  assign nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[431:424]));
  assign MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[439:432]));
  assign MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1181_nl = (readslicef_15_8_7(MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1181_nl = nl_MultLoop_acc_1181_nl[7:0];
  assign nl_MultLoop_acc_1267_nl = MultLoop_acc_1192_nl + MultLoop_acc_1191_nl +
      MultLoop_acc_1190_nl + MultLoop_acc_1189_nl + MultLoop_acc_1188_nl + MultLoop_acc_1187_nl
      + MultLoop_acc_1186_nl + MultLoop_acc_1185_nl + MultLoop_acc_1180_nl + MultLoop_acc_1179_nl
      + MultLoop_acc_1178_nl + MultLoop_acc_1177_nl + MultLoop_acc_1184_nl + MultLoop_acc_1183_nl
      + MultLoop_acc_1182_nl + MultLoop_acc_1181_nl;
  assign MultLoop_acc_1267_nl = nl_MultLoop_acc_1267_nl[7:0];
  assign nl_MultLoop_acc_1270_nl = MultLoop_acc_1268_nl + MultLoop_acc_1267_nl;
  assign MultLoop_acc_1270_nl = nl_MultLoop_acc_1270_nl[7:0];
  assign nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[575:568]));
  assign MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[583:576]));
  assign MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1172_nl = (readslicef_15_8_7(MultLoop_72_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_73_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1172_nl = nl_MultLoop_acc_1172_nl[7:0];
  assign nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[591:584]));
  assign MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[599:592]));
  assign MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1171_nl = (readslicef_15_8_7(MultLoop_74_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_75_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1171_nl = nl_MultLoop_acc_1171_nl[7:0];
  assign nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[703:696]));
  assign MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[711:704]));
  assign MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1164_nl = (readslicef_15_8_7(MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1164_nl = nl_MultLoop_acc_1164_nl[7:0];
  assign nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[719:712]));
  assign MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[727:720]));
  assign MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1163_nl = (readslicef_15_8_7(MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1163_nl = nl_MultLoop_acc_1163_nl[7:0];
  assign nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[639:632]));
  assign MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[647:640]));
  assign MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1168_nl = (readslicef_15_8_7(MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1168_nl = nl_MultLoop_acc_1168_nl[7:0];
  assign nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[655:648]));
  assign MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[663:656]));
  assign MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1167_nl = (readslicef_15_8_7(MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1167_nl = nl_MultLoop_acc_1167_nl[7:0];
  assign nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[959:952]));
  assign MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[967:960]));
  assign MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1148_nl = (readslicef_15_8_7(MultLoop_120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1148_nl = nl_MultLoop_acc_1148_nl[7:0];
  assign nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[975:968]));
  assign MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[983:976]));
  assign MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1147_nl = (readslicef_15_8_7(MultLoop_122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1147_nl = nl_MultLoop_acc_1147_nl[7:0];
  assign nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[895:888]));
  assign MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[903:896]));
  assign MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1152_nl = (readslicef_15_8_7(MultLoop_112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1152_nl = nl_MultLoop_acc_1152_nl[7:0];
  assign nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[911:904]));
  assign MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[919:912]));
  assign MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1151_nl = (readslicef_15_8_7(MultLoop_114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1151_nl = nl_MultLoop_acc_1151_nl[7:0];
  assign nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[927:920]));
  assign MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[935:928]));
  assign MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1150_nl = (readslicef_15_8_7(MultLoop_116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1150_nl = nl_MultLoop_acc_1150_nl[7:0];
  assign nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[943:936]));
  assign MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[951:944]));
  assign MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1149_nl = (readslicef_15_8_7(MultLoop_118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1149_nl = nl_MultLoop_acc_1149_nl[7:0];
  assign nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[767:760]));
  assign MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[775:768]));
  assign MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1160_nl = (readslicef_15_8_7(MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_97_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1160_nl = nl_MultLoop_acc_1160_nl[7:0];
  assign nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[783:776]));
  assign MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[791:784]));
  assign MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1159_nl = (readslicef_15_8_7(MultLoop_98_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1159_nl = nl_MultLoop_acc_1159_nl[7:0];
  assign nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[799:792]));
  assign MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[807:800]));
  assign MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1158_nl = (readslicef_15_8_7(MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1158_nl = nl_MultLoop_acc_1158_nl[7:0];
  assign nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[815:808]));
  assign MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[823:816]));
  assign MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1157_nl = (readslicef_15_8_7(MultLoop_102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1157_nl = nl_MultLoop_acc_1157_nl[7:0];
  assign nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[831:824]));
  assign MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[839:832]));
  assign MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1156_nl = (readslicef_15_8_7(MultLoop_104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1156_nl = nl_MultLoop_acc_1156_nl[7:0];
  assign nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[847:840]));
  assign MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[855:848]));
  assign MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1155_nl = (readslicef_15_8_7(MultLoop_106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1155_nl = nl_MultLoop_acc_1155_nl[7:0];
  assign nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[863:856]));
  assign MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[871:864]));
  assign MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1154_nl = (readslicef_15_8_7(MultLoop_108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1154_nl = nl_MultLoop_acc_1154_nl[7:0];
  assign nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[879:872]));
  assign MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[887:880]));
  assign MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1153_nl = (readslicef_15_8_7(MultLoop_110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1153_nl = nl_MultLoop_acc_1153_nl[7:0];
  assign nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[511:504]));
  assign MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[519:512]));
  assign MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1176_nl = (readslicef_15_8_7(MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1176_nl = nl_MultLoop_acc_1176_nl[7:0];
  assign nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[527:520]));
  assign MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[535:528]));
  assign MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1175_nl = (readslicef_15_8_7(MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1175_nl = nl_MultLoop_acc_1175_nl[7:0];
  assign nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[543:536]));
  assign MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[551:544]));
  assign MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1174_nl = (readslicef_15_8_7(MultLoop_68_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_69_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1174_nl = nl_MultLoop_acc_1174_nl[7:0];
  assign nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[559:552]));
  assign MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[567:560]));
  assign MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1173_nl = (readslicef_15_8_7(MultLoop_70_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_71_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1173_nl = nl_MultLoop_acc_1173_nl[7:0];
  assign nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[607:600]));
  assign MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[615:608]));
  assign MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1170_nl = (readslicef_15_8_7(MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1170_nl = nl_MultLoop_acc_1170_nl[7:0];
  assign nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[623:616]));
  assign MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[631:624]));
  assign MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1169_nl = (readslicef_15_8_7(MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1169_nl = nl_MultLoop_acc_1169_nl[7:0];
  assign nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[671:664]));
  assign MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[679:672]));
  assign MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1166_nl = (readslicef_15_8_7(MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1166_nl = nl_MultLoop_acc_1166_nl[7:0];
  assign nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[687:680]));
  assign MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[695:688]));
  assign MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1165_nl = (readslicef_15_8_7(MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1165_nl = nl_MultLoop_acc_1165_nl[7:0];
  assign nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[735:728]));
  assign MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[743:736]));
  assign MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1162_nl = (readslicef_15_8_7(MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1162_nl = nl_MultLoop_acc_1162_nl[7:0];
  assign nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[751:744]));
  assign MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[759:752]));
  assign MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1161_nl = (readslicef_15_8_7(MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1161_nl = nl_MultLoop_acc_1161_nl[7:0];
  assign nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[991:984]));
  assign MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[999:992]));
  assign MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1146_nl = (readslicef_15_8_7(MultLoop_124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1146_nl = nl_MultLoop_acc_1146_nl[7:0];
  assign nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1007:1000]));
  assign MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1015:1008]));
  assign MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1145_nl = (readslicef_15_8_7(MultLoop_126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1145_nl = nl_MultLoop_acc_1145_nl[7:0];
  assign nl_MultLoop_acc_1269_nl = MultLoop_acc_1172_nl + MultLoop_acc_1171_nl +
      MultLoop_acc_1164_nl + MultLoop_acc_1163_nl + MultLoop_acc_1168_nl + MultLoop_acc_1167_nl
      + MultLoop_acc_1148_nl + MultLoop_acc_1147_nl + MultLoop_acc_1152_nl + MultLoop_acc_1151_nl
      + MultLoop_acc_1150_nl + MultLoop_acc_1149_nl + MultLoop_acc_1160_nl + MultLoop_acc_1159_nl
      + MultLoop_acc_1158_nl + MultLoop_acc_1157_nl + MultLoop_acc_1156_nl + MultLoop_acc_1155_nl
      + MultLoop_acc_1154_nl + MultLoop_acc_1153_nl + MultLoop_acc_1176_nl + MultLoop_acc_1175_nl
      + MultLoop_acc_1174_nl + MultLoop_acc_1173_nl + MultLoop_acc_1170_nl + MultLoop_acc_1169_nl
      + MultLoop_acc_1166_nl + MultLoop_acc_1165_nl + MultLoop_acc_1162_nl + MultLoop_acc_1161_nl
      + MultLoop_acc_1146_nl + MultLoop_acc_1145_nl;
  assign MultLoop_acc_1269_nl = nl_MultLoop_acc_1269_nl[7:0];
  assign nl_layer4_out_0_sva_1 = MultLoop_acc_1270_nl + MultLoop_acc_1269_nl;
  assign layer4_out_0_sva_1 = nl_layer4_out_0_sva_1[7:0];
  assign nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10239:10232]));
  assign MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1017_nl = (readslicef_15_8_7(MultLoop_1280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[69:63]);
  assign MultLoop_acc_1017_nl = nl_MultLoop_acc_1017_nl[7:0];
  assign nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[9223:9216]));
  assign MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1081_nl = MultLoop_acc_1017_nl + (readslicef_15_8_7(MultLoop_1153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1081_nl = nl_MultLoop_acc_1081_nl[7:0];
  assign nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9231:9224]));
  assign MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9239:9232]));
  assign MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1080_nl = (readslicef_15_8_7(MultLoop_1154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1080_nl = nl_MultLoop_acc_1080_nl[7:0];
  assign nl_MultLoop_acc_1113_nl = MultLoop_acc_1081_nl + MultLoop_acc_1080_nl;
  assign MultLoop_acc_1113_nl = nl_MultLoop_acc_1113_nl[7:0];
  assign nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9247:9240]));
  assign MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9255:9248]));
  assign MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1079_nl = (readslicef_15_8_7(MultLoop_1156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1079_nl = nl_MultLoop_acc_1079_nl[7:0];
  assign nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9263:9256]));
  assign MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9271:9264]));
  assign MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1078_nl = (readslicef_15_8_7(MultLoop_1158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1078_nl = nl_MultLoop_acc_1078_nl[7:0];
  assign nl_MultLoop_acc_1112_nl = MultLoop_acc_1079_nl + MultLoop_acc_1078_nl;
  assign MultLoop_acc_1112_nl = nl_MultLoop_acc_1112_nl[7:0];
  assign nl_MultLoop_acc_1129_nl = MultLoop_acc_1113_nl + MultLoop_acc_1112_nl;
  assign MultLoop_acc_1129_nl = nl_MultLoop_acc_1129_nl[7:0];
  assign nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9279:9272]));
  assign MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9287:9280]));
  assign MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1077_nl = (readslicef_15_8_7(MultLoop_1160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1077_nl = nl_MultLoop_acc_1077_nl[7:0];
  assign nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9295:9288]));
  assign MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9303:9296]));
  assign MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1076_nl = (readslicef_15_8_7(MultLoop_1162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1076_nl = nl_MultLoop_acc_1076_nl[7:0];
  assign nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9311:9304]));
  assign MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9319:9312]));
  assign MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1075_nl = (readslicef_15_8_7(MultLoop_1164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1075_nl = nl_MultLoop_acc_1075_nl[7:0];
  assign nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9327:9320]));
  assign MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9335:9328]));
  assign MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1074_nl = (readslicef_15_8_7(MultLoop_1166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1074_nl = nl_MultLoop_acc_1074_nl[7:0];
  assign nl_MultLoop_acc_1128_nl = MultLoop_acc_1077_nl + MultLoop_acc_1076_nl +
      MultLoop_acc_1075_nl + MultLoop_acc_1074_nl;
  assign MultLoop_acc_1128_nl = nl_MultLoop_acc_1128_nl[7:0];
  assign nl_MultLoop_acc_1137_nl = MultLoop_acc_1129_nl + MultLoop_acc_1128_nl;
  assign MultLoop_acc_1137_nl = nl_MultLoop_acc_1137_nl[7:0];
  assign nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9407:9400]));
  assign MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9415:9408]));
  assign MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1069_nl = (readslicef_15_8_7(MultLoop_1176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1069_nl = nl_MultLoop_acc_1069_nl[7:0];
  assign nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9423:9416]));
  assign MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9431:9424]));
  assign MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1068_nl = (readslicef_15_8_7(MultLoop_1178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1068_nl = nl_MultLoop_acc_1068_nl[7:0];
  assign nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9343:9336]));
  assign MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9351:9344]));
  assign MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1073_nl = (readslicef_15_8_7(MultLoop_1168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1073_nl = nl_MultLoop_acc_1073_nl[7:0];
  assign nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9359:9352]));
  assign MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9367:9360]));
  assign MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1072_nl = (readslicef_15_8_7(MultLoop_1170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1072_nl = nl_MultLoop_acc_1072_nl[7:0];
  assign nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9375:9368]));
  assign MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9383:9376]));
  assign MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1071_nl = (readslicef_15_8_7(MultLoop_1172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1071_nl = nl_MultLoop_acc_1071_nl[7:0];
  assign nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9391:9384]));
  assign MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9399:9392]));
  assign MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1070_nl = (readslicef_15_8_7(MultLoop_1174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1070_nl = nl_MultLoop_acc_1070_nl[7:0];
  assign nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9439:9432]));
  assign MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9447:9440]));
  assign MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1067_nl = (readslicef_15_8_7(MultLoop_1180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1067_nl = nl_MultLoop_acc_1067_nl[7:0];
  assign nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9455:9448]));
  assign MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9463:9456]));
  assign MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1066_nl = (readslicef_15_8_7(MultLoop_1182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1066_nl = nl_MultLoop_acc_1066_nl[7:0];
  assign nl_MultLoop_acc_1136_nl = MultLoop_acc_1069_nl + MultLoop_acc_1068_nl +
      MultLoop_acc_1073_nl + MultLoop_acc_1072_nl + MultLoop_acc_1071_nl + MultLoop_acc_1070_nl
      + MultLoop_acc_1067_nl + MultLoop_acc_1066_nl;
  assign MultLoop_acc_1136_nl = nl_MultLoop_acc_1136_nl[7:0];
  assign nl_MultLoop_acc_1141_nl = MultLoop_acc_1137_nl + MultLoop_acc_1136_nl;
  assign MultLoop_acc_1141_nl = nl_MultLoop_acc_1141_nl[7:0];
  assign nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9471:9464]));
  assign MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9479:9472]));
  assign MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1065_nl = (readslicef_15_8_7(MultLoop_1184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1065_nl = nl_MultLoop_acc_1065_nl[7:0];
  assign nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9487:9480]));
  assign MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9495:9488]));
  assign MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1064_nl = (readslicef_15_8_7(MultLoop_1186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1064_nl = nl_MultLoop_acc_1064_nl[7:0];
  assign nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9503:9496]));
  assign MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9511:9504]));
  assign MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1063_nl = (readslicef_15_8_7(MultLoop_1188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1063_nl = nl_MultLoop_acc_1063_nl[7:0];
  assign nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9519:9512]));
  assign MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9527:9520]));
  assign MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1062_nl = (readslicef_15_8_7(MultLoop_1190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1062_nl = nl_MultLoop_acc_1062_nl[7:0];
  assign nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9535:9528]));
  assign MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9543:9536]));
  assign MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1061_nl = (readslicef_15_8_7(MultLoop_1192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1061_nl = nl_MultLoop_acc_1061_nl[7:0];
  assign nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9551:9544]));
  assign MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9559:9552]));
  assign MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1060_nl = (readslicef_15_8_7(MultLoop_1194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1060_nl = nl_MultLoop_acc_1060_nl[7:0];
  assign nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9567:9560]));
  assign MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9575:9568]));
  assign MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1059_nl = (readslicef_15_8_7(MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1059_nl = nl_MultLoop_acc_1059_nl[7:0];
  assign nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9583:9576]));
  assign MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9591:9584]));
  assign MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1058_nl = (readslicef_15_8_7(MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1058_nl = nl_MultLoop_acc_1058_nl[7:0];
  assign nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9663:9656]));
  assign MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9671:9664]));
  assign MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1053_nl = (readslicef_15_8_7(MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1053_nl = nl_MultLoop_acc_1053_nl[7:0];
  assign nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9679:9672]));
  assign MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9687:9680]));
  assign MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1052_nl = (readslicef_15_8_7(MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1052_nl = nl_MultLoop_acc_1052_nl[7:0];
  assign nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9695:9688]));
  assign MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9703:9696]));
  assign MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1051_nl = (readslicef_15_8_7(MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1051_nl = nl_MultLoop_acc_1051_nl[7:0];
  assign nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9711:9704]));
  assign MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9719:9712]));
  assign MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1050_nl = (readslicef_15_8_7(MultLoop_1214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1050_nl = nl_MultLoop_acc_1050_nl[7:0];
  assign nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9599:9592]));
  assign MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9607:9600]));
  assign MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1057_nl = (readslicef_15_8_7(MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1057_nl = nl_MultLoop_acc_1057_nl[7:0];
  assign nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9615:9608]));
  assign MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9623:9616]));
  assign MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1056_nl = (readslicef_15_8_7(MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1056_nl = nl_MultLoop_acc_1056_nl[7:0];
  assign nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9631:9624]));
  assign MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9639:9632]));
  assign MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1055_nl = (readslicef_15_8_7(MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1055_nl = nl_MultLoop_acc_1055_nl[7:0];
  assign nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9647:9640]));
  assign MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9655:9648]));
  assign MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1054_nl = (readslicef_15_8_7(MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1054_nl = nl_MultLoop_acc_1054_nl[7:0];
  assign nl_MultLoop_acc_1140_nl = MultLoop_acc_1065_nl + MultLoop_acc_1064_nl +
      MultLoop_acc_1063_nl + MultLoop_acc_1062_nl + MultLoop_acc_1061_nl + MultLoop_acc_1060_nl
      + MultLoop_acc_1059_nl + MultLoop_acc_1058_nl + MultLoop_acc_1053_nl + MultLoop_acc_1052_nl
      + MultLoop_acc_1051_nl + MultLoop_acc_1050_nl + MultLoop_acc_1057_nl + MultLoop_acc_1056_nl
      + MultLoop_acc_1055_nl + MultLoop_acc_1054_nl;
  assign MultLoop_acc_1140_nl = nl_MultLoop_acc_1140_nl[7:0];
  assign nl_MultLoop_acc_1143_nl = MultLoop_acc_1141_nl + MultLoop_acc_1140_nl;
  assign MultLoop_acc_1143_nl = nl_MultLoop_acc_1143_nl[7:0];
  assign nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9791:9784]));
  assign MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9799:9792]));
  assign MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1045_nl = (readslicef_15_8_7(MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1045_nl = nl_MultLoop_acc_1045_nl[7:0];
  assign nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9807:9800]));
  assign MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9815:9808]));
  assign MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1044_nl = (readslicef_15_8_7(MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1044_nl = nl_MultLoop_acc_1044_nl[7:0];
  assign nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9919:9912]));
  assign MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9927:9920]));
  assign MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1037_nl = (readslicef_15_8_7(MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1037_nl = nl_MultLoop_acc_1037_nl[7:0];
  assign nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9935:9928]));
  assign MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9943:9936]));
  assign MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1036_nl = (readslicef_15_8_7(MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1036_nl = nl_MultLoop_acc_1036_nl[7:0];
  assign nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9855:9848]));
  assign MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9863:9856]));
  assign MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1041_nl = (readslicef_15_8_7(MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1041_nl = nl_MultLoop_acc_1041_nl[7:0];
  assign nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9871:9864]));
  assign MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9879:9872]));
  assign MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1040_nl = (readslicef_15_8_7(MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1040_nl = nl_MultLoop_acc_1040_nl[7:0];
  assign nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10175:10168]));
  assign MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10183:10176]));
  assign MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1021_nl = (readslicef_15_8_7(MultLoop_1272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1021_nl = nl_MultLoop_acc_1021_nl[7:0];
  assign nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10191:10184]));
  assign MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10199:10192]));
  assign MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1020_nl = (readslicef_15_8_7(MultLoop_1274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1020_nl = nl_MultLoop_acc_1020_nl[7:0];
  assign nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10111:10104]));
  assign MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10119:10112]));
  assign MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1025_nl = (readslicef_15_8_7(MultLoop_1264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1025_nl = nl_MultLoop_acc_1025_nl[7:0];
  assign nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10127:10120]));
  assign MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10135:10128]));
  assign MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1024_nl = (readslicef_15_8_7(MultLoop_1266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1024_nl = nl_MultLoop_acc_1024_nl[7:0];
  assign nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10143:10136]));
  assign MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10151:10144]));
  assign MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1023_nl = (readslicef_15_8_7(MultLoop_1268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1023_nl = nl_MultLoop_acc_1023_nl[7:0];
  assign nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10159:10152]));
  assign MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10167:10160]));
  assign MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1022_nl = (readslicef_15_8_7(MultLoop_1270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1022_nl = nl_MultLoop_acc_1022_nl[7:0];
  assign nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9983:9976]));
  assign MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9991:9984]));
  assign MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1033_nl = (readslicef_15_8_7(MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1033_nl = nl_MultLoop_acc_1033_nl[7:0];
  assign nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9999:9992]));
  assign MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10007:10000]));
  assign MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1032_nl = (readslicef_15_8_7(MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1032_nl = nl_MultLoop_acc_1032_nl[7:0];
  assign nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10015:10008]));
  assign MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10023:10016]));
  assign MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1031_nl = (readslicef_15_8_7(MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1031_nl = nl_MultLoop_acc_1031_nl[7:0];
  assign nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10031:10024]));
  assign MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10039:10032]));
  assign MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1030_nl = (readslicef_15_8_7(MultLoop_1254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1030_nl = nl_MultLoop_acc_1030_nl[7:0];
  assign nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10047:10040]));
  assign MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10055:10048]));
  assign MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1029_nl = (readslicef_15_8_7(MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1029_nl = nl_MultLoop_acc_1029_nl[7:0];
  assign nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10063:10056]));
  assign MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10071:10064]));
  assign MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1028_nl = (readslicef_15_8_7(MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1028_nl = nl_MultLoop_acc_1028_nl[7:0];
  assign nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10079:10072]));
  assign MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10087:10080]));
  assign MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1027_nl = (readslicef_15_8_7(MultLoop_1260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1027_nl = nl_MultLoop_acc_1027_nl[7:0];
  assign nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10095:10088]));
  assign MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10103:10096]));
  assign MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1026_nl = (readslicef_15_8_7(MultLoop_1262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1026_nl = nl_MultLoop_acc_1026_nl[7:0];
  assign nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9727:9720]));
  assign MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9735:9728]));
  assign MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1049_nl = (readslicef_15_8_7(MultLoop_1216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1049_nl = nl_MultLoop_acc_1049_nl[7:0];
  assign nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9743:9736]));
  assign MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9751:9744]));
  assign MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1048_nl = (readslicef_15_8_7(MultLoop_1218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1048_nl = nl_MultLoop_acc_1048_nl[7:0];
  assign nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9759:9752]));
  assign MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9767:9760]));
  assign MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1047_nl = (readslicef_15_8_7(MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1047_nl = nl_MultLoop_acc_1047_nl[7:0];
  assign nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9775:9768]));
  assign MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9783:9776]));
  assign MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1046_nl = (readslicef_15_8_7(MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1046_nl = nl_MultLoop_acc_1046_nl[7:0];
  assign nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9823:9816]));
  assign MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9831:9824]));
  assign MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1043_nl = (readslicef_15_8_7(MultLoop_1228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1043_nl = nl_MultLoop_acc_1043_nl[7:0];
  assign nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9839:9832]));
  assign MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9847:9840]));
  assign MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1042_nl = (readslicef_15_8_7(MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1042_nl = nl_MultLoop_acc_1042_nl[7:0];
  assign nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9887:9880]));
  assign MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9895:9888]));
  assign MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1039_nl = (readslicef_15_8_7(MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1039_nl = nl_MultLoop_acc_1039_nl[7:0];
  assign nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9903:9896]));
  assign MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9911:9904]));
  assign MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1038_nl = (readslicef_15_8_7(MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1038_nl = nl_MultLoop_acc_1038_nl[7:0];
  assign nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9951:9944]));
  assign MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9959:9952]));
  assign MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1035_nl = (readslicef_15_8_7(MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1035_nl = nl_MultLoop_acc_1035_nl[7:0];
  assign nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9967:9960]));
  assign MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9975:9968]));
  assign MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1034_nl = (readslicef_15_8_7(MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1034_nl = nl_MultLoop_acc_1034_nl[7:0];
  assign nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10207:10200]));
  assign MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10215:10208]));
  assign MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1019_nl = (readslicef_15_8_7(MultLoop_1276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1019_nl = nl_MultLoop_acc_1019_nl[7:0];
  assign nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10223:10216]));
  assign MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[10231:10224]));
  assign MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_1018_nl = (readslicef_15_8_7(MultLoop_1278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_1018_nl = nl_MultLoop_acc_1018_nl[7:0];
  assign nl_MultLoop_acc_1142_nl = MultLoop_acc_1045_nl + MultLoop_acc_1044_nl +
      MultLoop_acc_1037_nl + MultLoop_acc_1036_nl + MultLoop_acc_1041_nl + MultLoop_acc_1040_nl
      + MultLoop_acc_1021_nl + MultLoop_acc_1020_nl + MultLoop_acc_1025_nl + MultLoop_acc_1024_nl
      + MultLoop_acc_1023_nl + MultLoop_acc_1022_nl + MultLoop_acc_1033_nl + MultLoop_acc_1032_nl
      + MultLoop_acc_1031_nl + MultLoop_acc_1030_nl + MultLoop_acc_1029_nl + MultLoop_acc_1028_nl
      + MultLoop_acc_1027_nl + MultLoop_acc_1026_nl + MultLoop_acc_1049_nl + MultLoop_acc_1048_nl
      + MultLoop_acc_1047_nl + MultLoop_acc_1046_nl + MultLoop_acc_1043_nl + MultLoop_acc_1042_nl
      + MultLoop_acc_1039_nl + MultLoop_acc_1038_nl + MultLoop_acc_1035_nl + MultLoop_acc_1034_nl
      + MultLoop_acc_1019_nl + MultLoop_acc_1018_nl;
  assign MultLoop_acc_1142_nl = nl_MultLoop_acc_1142_nl[7:0];
  assign nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1 = MultLoop_acc_1143_nl + MultLoop_acc_1142_nl;
  assign MultLoop_1280_MultLoop_acc_3_ncse_sva_1 = nl_MultLoop_1280_MultLoop_acc_3_ncse_sva_1[7:0];
  assign nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2047:2040]));
  assign MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_65_nl = (readslicef_15_8_7(MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[13:7]);
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[7:0];
  assign nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[1031:1024]));
  assign MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_97_nl = MultLoop_acc_65_nl + (readslicef_15_8_7(MultLoop_129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_97_nl = nl_MultLoop_acc_97_nl[7:0];
  assign nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1039:1032]));
  assign MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1047:1040]));
  assign MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_64_nl = (readslicef_15_8_7(MultLoop_130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_64_nl = nl_MultLoop_acc_64_nl[7:0];
  assign nl_MultLoop_acc_113_nl = MultLoop_acc_97_nl + MultLoop_acc_64_nl;
  assign MultLoop_acc_113_nl = nl_MultLoop_acc_113_nl[7:0];
  assign nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1055:1048]));
  assign MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1063:1056]));
  assign MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_63_nl = (readslicef_15_8_7(MultLoop_132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_63_nl = nl_MultLoop_acc_63_nl[7:0];
  assign nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1071:1064]));
  assign MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1079:1072]));
  assign MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_62_nl = (readslicef_15_8_7(MultLoop_134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_62_nl = nl_MultLoop_acc_62_nl[7:0];
  assign nl_MultLoop_acc_96_nl = MultLoop_acc_63_nl + MultLoop_acc_62_nl;
  assign MultLoop_acc_96_nl = nl_MultLoop_acc_96_nl[7:0];
  assign nl_MultLoop_acc_121_nl = MultLoop_acc_113_nl + MultLoop_acc_96_nl;
  assign MultLoop_acc_121_nl = nl_MultLoop_acc_121_nl[7:0];
  assign nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1087:1080]));
  assign MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1095:1088]));
  assign MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_61_nl = (readslicef_15_8_7(MultLoop_136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_61_nl = nl_MultLoop_acc_61_nl[7:0];
  assign nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1103:1096]));
  assign MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1111:1104]));
  assign MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_60_nl = (readslicef_15_8_7(MultLoop_138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_60_nl = nl_MultLoop_acc_60_nl[7:0];
  assign nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1119:1112]));
  assign MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1127:1120]));
  assign MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_59_nl = (readslicef_15_8_7(MultLoop_140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_59_nl = nl_MultLoop_acc_59_nl[7:0];
  assign nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1135:1128]));
  assign MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1143:1136]));
  assign MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_58_nl = (readslicef_15_8_7(MultLoop_142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_58_nl = nl_MultLoop_acc_58_nl[7:0];
  assign nl_MultLoop_acc_112_nl = MultLoop_acc_61_nl + MultLoop_acc_60_nl + MultLoop_acc_59_nl
      + MultLoop_acc_58_nl;
  assign MultLoop_acc_112_nl = nl_MultLoop_acc_112_nl[7:0];
  assign nl_MultLoop_acc_125_nl = MultLoop_acc_121_nl + MultLoop_acc_112_nl;
  assign MultLoop_acc_125_nl = nl_MultLoop_acc_125_nl[7:0];
  assign nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1215:1208]));
  assign MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1223:1216]));
  assign MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_53_nl = (readslicef_15_8_7(MultLoop_152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_153_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[7:0];
  assign nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1231:1224]));
  assign MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1239:1232]));
  assign MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_52_nl = (readslicef_15_8_7(MultLoop_154_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_155_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_52_nl = nl_MultLoop_acc_52_nl[7:0];
  assign nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1151:1144]));
  assign MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1159:1152]));
  assign MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_57_nl = (readslicef_15_8_7(MultLoop_144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_57_nl = nl_MultLoop_acc_57_nl[7:0];
  assign nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1167:1160]));
  assign MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1175:1168]));
  assign MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_56_nl = (readslicef_15_8_7(MultLoop_146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_56_nl = nl_MultLoop_acc_56_nl[7:0];
  assign nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1183:1176]));
  assign MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1191:1184]));
  assign MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_55_nl = (readslicef_15_8_7(MultLoop_148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_55_nl = nl_MultLoop_acc_55_nl[7:0];
  assign nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1199:1192]));
  assign MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1207:1200]));
  assign MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_54_nl = (readslicef_15_8_7(MultLoop_150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_54_nl = nl_MultLoop_acc_54_nl[7:0];
  assign nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1247:1240]));
  assign MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1255:1248]));
  assign MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_51_nl = (readslicef_15_8_7(MultLoop_156_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_157_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_51_nl = nl_MultLoop_acc_51_nl[7:0];
  assign nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1263:1256]));
  assign MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1271:1264]));
  assign MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_50_nl = (readslicef_15_8_7(MultLoop_158_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_159_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_50_nl = nl_MultLoop_acc_50_nl[7:0];
  assign nl_MultLoop_acc_120_nl = MultLoop_acc_53_nl + MultLoop_acc_52_nl + MultLoop_acc_57_nl
      + MultLoop_acc_56_nl + MultLoop_acc_55_nl + MultLoop_acc_54_nl + MultLoop_acc_51_nl
      + MultLoop_acc_50_nl;
  assign MultLoop_acc_120_nl = nl_MultLoop_acc_120_nl[7:0];
  assign nl_MultLoop_acc_127_nl = MultLoop_acc_125_nl + MultLoop_acc_120_nl;
  assign MultLoop_acc_127_nl = nl_MultLoop_acc_127_nl[7:0];
  assign nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1279:1272]));
  assign MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1287:1280]));
  assign MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_49_nl = (readslicef_15_8_7(MultLoop_160_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_161_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_49_nl = nl_MultLoop_acc_49_nl[7:0];
  assign nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1295:1288]));
  assign MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1303:1296]));
  assign MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_48_nl = (readslicef_15_8_7(MultLoop_162_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_163_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_48_nl = nl_MultLoop_acc_48_nl[7:0];
  assign nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1311:1304]));
  assign MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1319:1312]));
  assign MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_47_nl = (readslicef_15_8_7(MultLoop_164_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_165_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_47_nl = nl_MultLoop_acc_47_nl[7:0];
  assign nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1327:1320]));
  assign MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1335:1328]));
  assign MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_46_nl = (readslicef_15_8_7(MultLoop_166_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_167_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_46_nl = nl_MultLoop_acc_46_nl[7:0];
  assign nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1343:1336]));
  assign MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1351:1344]));
  assign MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_45_nl = (readslicef_15_8_7(MultLoop_168_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_169_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[7:0];
  assign nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1359:1352]));
  assign MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1367:1360]));
  assign MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_44_nl = (readslicef_15_8_7(MultLoop_170_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_171_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_44_nl = nl_MultLoop_acc_44_nl[7:0];
  assign nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1375:1368]));
  assign MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1383:1376]));
  assign MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_43_nl = (readslicef_15_8_7(MultLoop_172_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_173_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_43_nl = nl_MultLoop_acc_43_nl[7:0];
  assign nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1391:1384]));
  assign MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1399:1392]));
  assign MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_42_nl = (readslicef_15_8_7(MultLoop_174_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_175_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[7:0];
  assign nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1471:1464]));
  assign MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1479:1472]));
  assign MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_37_nl = (readslicef_15_8_7(MultLoop_184_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_185_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_37_nl = nl_MultLoop_acc_37_nl[7:0];
  assign nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1487:1480]));
  assign MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1495:1488]));
  assign MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_36_nl = (readslicef_15_8_7(MultLoop_186_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_187_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_36_nl = nl_MultLoop_acc_36_nl[7:0];
  assign nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1503:1496]));
  assign MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1511:1504]));
  assign MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_35_nl = (readslicef_15_8_7(MultLoop_188_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_189_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_35_nl = nl_MultLoop_acc_35_nl[7:0];
  assign nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1519:1512]));
  assign MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1527:1520]));
  assign MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_34_nl = (readslicef_15_8_7(MultLoop_190_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_191_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_34_nl = nl_MultLoop_acc_34_nl[7:0];
  assign nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1407:1400]));
  assign MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1415:1408]));
  assign MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_41_nl = (readslicef_15_8_7(MultLoop_176_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_177_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_41_nl = nl_MultLoop_acc_41_nl[7:0];
  assign nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1423:1416]));
  assign MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1431:1424]));
  assign MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_40_nl = (readslicef_15_8_7(MultLoop_178_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_179_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_40_nl = nl_MultLoop_acc_40_nl[7:0];
  assign nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1439:1432]));
  assign MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1447:1440]));
  assign MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_39_nl = (readslicef_15_8_7(MultLoop_180_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_181_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_39_nl = nl_MultLoop_acc_39_nl[7:0];
  assign nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1455:1448]));
  assign MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1463:1456]));
  assign MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_38_nl = (readslicef_15_8_7(MultLoop_182_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_183_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_38_nl = nl_MultLoop_acc_38_nl[7:0];
  assign nl_MultLoop_acc_124_nl = MultLoop_acc_49_nl + MultLoop_acc_48_nl + MultLoop_acc_47_nl
      + MultLoop_acc_46_nl + MultLoop_acc_45_nl + MultLoop_acc_44_nl + MultLoop_acc_43_nl
      + MultLoop_acc_42_nl + MultLoop_acc_37_nl + MultLoop_acc_36_nl + MultLoop_acc_35_nl
      + MultLoop_acc_34_nl + MultLoop_acc_41_nl + MultLoop_acc_40_nl + MultLoop_acc_39_nl
      + MultLoop_acc_38_nl;
  assign MultLoop_acc_124_nl = nl_MultLoop_acc_124_nl[7:0];
  assign nl_MultLoop_acc_nl = MultLoop_acc_127_nl + MultLoop_acc_124_nl;
  assign MultLoop_acc_nl = nl_MultLoop_acc_nl[7:0];
  assign nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1599:1592]));
  assign MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1607:1600]));
  assign MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_29_nl = (readslicef_15_8_7(MultLoop_200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_29_nl = nl_MultLoop_acc_29_nl[7:0];
  assign nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1615:1608]));
  assign MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1623:1616]));
  assign MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_28_nl = (readslicef_15_8_7(MultLoop_202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_28_nl = nl_MultLoop_acc_28_nl[7:0];
  assign nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1727:1720]));
  assign MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1735:1728]));
  assign MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_21_nl = (readslicef_15_8_7(MultLoop_216_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_217_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[7:0];
  assign nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1743:1736]));
  assign MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1751:1744]));
  assign MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_20_nl = (readslicef_15_8_7(MultLoop_218_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_219_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_20_nl = nl_MultLoop_acc_20_nl[7:0];
  assign nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1663:1656]));
  assign MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1671:1664]));
  assign MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_25_nl = (readslicef_15_8_7(MultLoop_208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_25_nl = nl_MultLoop_acc_25_nl[7:0];
  assign nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1679:1672]));
  assign MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1687:1680]));
  assign MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_24_nl = (readslicef_15_8_7(MultLoop_210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_24_nl = nl_MultLoop_acc_24_nl[7:0];
  assign nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1983:1976]));
  assign MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1991:1984]));
  assign MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_5_nl = (readslicef_15_8_7(MultLoop_248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_5_nl = nl_MultLoop_acc_5_nl[7:0];
  assign nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1999:1992]));
  assign MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2007:2000]));
  assign MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_4_nl = (readslicef_15_8_7(MultLoop_250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_4_nl = nl_MultLoop_acc_4_nl[7:0];
  assign nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1919:1912]));
  assign MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1927:1920]));
  assign MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_9_nl = (readslicef_15_8_7(MultLoop_240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_9_nl = nl_MultLoop_acc_9_nl[7:0];
  assign nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1935:1928]));
  assign MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1943:1936]));
  assign MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_8_nl = (readslicef_15_8_7(MultLoop_242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_8_nl = nl_MultLoop_acc_8_nl[7:0];
  assign nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1951:1944]));
  assign MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1959:1952]));
  assign MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_7_nl = (readslicef_15_8_7(MultLoop_244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_7_nl = nl_MultLoop_acc_7_nl[7:0];
  assign nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1967:1960]));
  assign MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1975:1968]));
  assign MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_6_nl = (readslicef_15_8_7(MultLoop_246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_6_nl = nl_MultLoop_acc_6_nl[7:0];
  assign nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1791:1784]));
  assign MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1799:1792]));
  assign MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_17_nl = (readslicef_15_8_7(MultLoop_224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_17_nl = nl_MultLoop_acc_17_nl[7:0];
  assign nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1807:1800]));
  assign MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1815:1808]));
  assign MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_16_nl = (readslicef_15_8_7(MultLoop_226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_16_nl = nl_MultLoop_acc_16_nl[7:0];
  assign nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1823:1816]));
  assign MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1831:1824]));
  assign MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_15_nl = (readslicef_15_8_7(MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_15_nl = nl_MultLoop_acc_15_nl[7:0];
  assign nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1839:1832]));
  assign MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1847:1840]));
  assign MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_14_nl = (readslicef_15_8_7(MultLoop_230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[7:0];
  assign nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1855:1848]));
  assign MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1863:1856]));
  assign MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_13_nl = (readslicef_15_8_7(MultLoop_232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_233_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_13_nl = nl_MultLoop_acc_13_nl[7:0];
  assign nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1871:1864]));
  assign MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1879:1872]));
  assign MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_12_nl = (readslicef_15_8_7(MultLoop_234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_12_nl = nl_MultLoop_acc_12_nl[7:0];
  assign nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1887:1880]));
  assign MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1895:1888]));
  assign MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_11_nl = (readslicef_15_8_7(MultLoop_236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_11_nl = nl_MultLoop_acc_11_nl[7:0];
  assign nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1903:1896]));
  assign MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1911:1904]));
  assign MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_10_nl = (readslicef_15_8_7(MultLoop_238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_10_nl = nl_MultLoop_acc_10_nl[7:0];
  assign nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1535:1528]));
  assign MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1543:1536]));
  assign MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_33_nl = (readslicef_15_8_7(MultLoop_192_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_33_nl = nl_MultLoop_acc_33_nl[7:0];
  assign nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1551:1544]));
  assign MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1559:1552]));
  assign MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_32_nl = (readslicef_15_8_7(MultLoop_194_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_32_nl = nl_MultLoop_acc_32_nl[7:0];
  assign nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1567:1560]));
  assign MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1575:1568]));
  assign MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_31_nl = (readslicef_15_8_7(MultLoop_196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_31_nl = nl_MultLoop_acc_31_nl[7:0];
  assign nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1583:1576]));
  assign MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1591:1584]));
  assign MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_30_nl = (readslicef_15_8_7(MultLoop_198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_30_nl = nl_MultLoop_acc_30_nl[7:0];
  assign nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1631:1624]));
  assign MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1639:1632]));
  assign MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_27_nl = (readslicef_15_8_7(MultLoop_204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_27_nl = nl_MultLoop_acc_27_nl[7:0];
  assign nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1647:1640]));
  assign MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1655:1648]));
  assign MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_26_nl = (readslicef_15_8_7(MultLoop_206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_26_nl = nl_MultLoop_acc_26_nl[7:0];
  assign nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1695:1688]));
  assign MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1703:1696]));
  assign MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_23_nl = (readslicef_15_8_7(MultLoop_212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_23_nl = nl_MultLoop_acc_23_nl[7:0];
  assign nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1711:1704]));
  assign MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1719:1712]));
  assign MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_22_nl = (readslicef_15_8_7(MultLoop_214_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_215_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_22_nl = nl_MultLoop_acc_22_nl[7:0];
  assign nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1759:1752]));
  assign MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1767:1760]));
  assign MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_19_nl = (readslicef_15_8_7(MultLoop_220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_19_nl = nl_MultLoop_acc_19_nl[7:0];
  assign nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1775:1768]));
  assign MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[1783:1776]));
  assign MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_18_nl = (readslicef_15_8_7(MultLoop_222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[7:0];
  assign nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2015:2008]));
  assign MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2023:2016]));
  assign MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_3_nl = (readslicef_15_8_7(MultLoop_252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_253_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_3_nl = nl_MultLoop_acc_3_nl[7:0];
  assign nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2031:2024]));
  assign MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2039:2032]));
  assign MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_2_nl = (readslicef_15_8_7(MultLoop_254_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_2_nl = nl_MultLoop_acc_2_nl[7:0];
  assign nl_MultLoop_acc_126_nl = MultLoop_acc_29_nl + MultLoop_acc_28_nl + MultLoop_acc_21_nl
      + MultLoop_acc_20_nl + MultLoop_acc_25_nl + MultLoop_acc_24_nl + MultLoop_acc_5_nl
      + MultLoop_acc_4_nl + MultLoop_acc_9_nl + MultLoop_acc_8_nl + MultLoop_acc_7_nl
      + MultLoop_acc_6_nl + MultLoop_acc_17_nl + MultLoop_acc_16_nl + MultLoop_acc_15_nl
      + MultLoop_acc_14_nl + MultLoop_acc_13_nl + MultLoop_acc_12_nl + MultLoop_acc_11_nl
      + MultLoop_acc_10_nl + MultLoop_acc_33_nl + MultLoop_acc_32_nl + MultLoop_acc_31_nl
      + MultLoop_acc_30_nl + MultLoop_acc_27_nl + MultLoop_acc_26_nl + MultLoop_acc_23_nl
      + MultLoop_acc_22_nl + MultLoop_acc_19_nl + MultLoop_acc_18_nl + MultLoop_acc_3_nl
      + MultLoop_acc_2_nl;
  assign MultLoop_acc_126_nl = nl_MultLoop_acc_126_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1 = MultLoop_acc_nl
      + MultLoop_acc_126_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1[7:0];
  assign nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9215:9208]));
  assign MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_890_nl = (readslicef_15_8_7(MultLoop_1152_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[62:56]);
  assign MultLoop_acc_890_nl = nl_MultLoop_acc_890_nl[7:0];
  assign nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[8199:8192]));
  assign MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_954_nl = MultLoop_acc_890_nl + (readslicef_15_8_7(MultLoop_1025_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_954_nl = nl_MultLoop_acc_954_nl[7:0];
  assign nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8207:8200]));
  assign MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8215:8208]));
  assign MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_953_nl = (readslicef_15_8_7(MultLoop_1026_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1027_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_953_nl = nl_MultLoop_acc_953_nl[7:0];
  assign nl_MultLoop_acc_986_nl = MultLoop_acc_954_nl + MultLoop_acc_953_nl;
  assign MultLoop_acc_986_nl = nl_MultLoop_acc_986_nl[7:0];
  assign nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8223:8216]));
  assign MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8231:8224]));
  assign MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_952_nl = (readslicef_15_8_7(MultLoop_1028_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1029_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_952_nl = nl_MultLoop_acc_952_nl[7:0];
  assign nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8239:8232]));
  assign MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8247:8240]));
  assign MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_951_nl = (readslicef_15_8_7(MultLoop_1030_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1031_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_951_nl = nl_MultLoop_acc_951_nl[7:0];
  assign nl_MultLoop_acc_985_nl = MultLoop_acc_952_nl + MultLoop_acc_951_nl;
  assign MultLoop_acc_985_nl = nl_MultLoop_acc_985_nl[7:0];
  assign nl_MultLoop_acc_1002_nl = MultLoop_acc_986_nl + MultLoop_acc_985_nl;
  assign MultLoop_acc_1002_nl = nl_MultLoop_acc_1002_nl[7:0];
  assign nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8255:8248]));
  assign MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8263:8256]));
  assign MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_950_nl = (readslicef_15_8_7(MultLoop_1032_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1033_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_950_nl = nl_MultLoop_acc_950_nl[7:0];
  assign nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8271:8264]));
  assign MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8279:8272]));
  assign MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_949_nl = (readslicef_15_8_7(MultLoop_1034_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1035_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_949_nl = nl_MultLoop_acc_949_nl[7:0];
  assign nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8287:8280]));
  assign MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8295:8288]));
  assign MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_948_nl = (readslicef_15_8_7(MultLoop_1036_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1037_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_948_nl = nl_MultLoop_acc_948_nl[7:0];
  assign nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8303:8296]));
  assign MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8311:8304]));
  assign MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_947_nl = (readslicef_15_8_7(MultLoop_1038_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1039_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_947_nl = nl_MultLoop_acc_947_nl[7:0];
  assign nl_MultLoop_acc_1001_nl = MultLoop_acc_950_nl + MultLoop_acc_949_nl + MultLoop_acc_948_nl
      + MultLoop_acc_947_nl;
  assign MultLoop_acc_1001_nl = nl_MultLoop_acc_1001_nl[7:0];
  assign nl_MultLoop_acc_1010_nl = MultLoop_acc_1002_nl + MultLoop_acc_1001_nl;
  assign MultLoop_acc_1010_nl = nl_MultLoop_acc_1010_nl[7:0];
  assign nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8383:8376]));
  assign MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8391:8384]));
  assign MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_942_nl = (readslicef_15_8_7(MultLoop_1048_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1049_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_942_nl = nl_MultLoop_acc_942_nl[7:0];
  assign nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8399:8392]));
  assign MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8407:8400]));
  assign MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_941_nl = (readslicef_15_8_7(MultLoop_1050_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1051_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_941_nl = nl_MultLoop_acc_941_nl[7:0];
  assign nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8319:8312]));
  assign MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8327:8320]));
  assign MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_946_nl = (readslicef_15_8_7(MultLoop_1040_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1041_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_946_nl = nl_MultLoop_acc_946_nl[7:0];
  assign nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8335:8328]));
  assign MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8343:8336]));
  assign MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_945_nl = (readslicef_15_8_7(MultLoop_1042_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1043_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_945_nl = nl_MultLoop_acc_945_nl[7:0];
  assign nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8351:8344]));
  assign MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8359:8352]));
  assign MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_944_nl = (readslicef_15_8_7(MultLoop_1044_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1045_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_944_nl = nl_MultLoop_acc_944_nl[7:0];
  assign nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8367:8360]));
  assign MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8375:8368]));
  assign MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_943_nl = (readslicef_15_8_7(MultLoop_1046_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1047_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_943_nl = nl_MultLoop_acc_943_nl[7:0];
  assign nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8415:8408]));
  assign MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8423:8416]));
  assign MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_940_nl = (readslicef_15_8_7(MultLoop_1052_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1053_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_940_nl = nl_MultLoop_acc_940_nl[7:0];
  assign nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8431:8424]));
  assign MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8439:8432]));
  assign MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_939_nl = (readslicef_15_8_7(MultLoop_1054_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1055_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_939_nl = nl_MultLoop_acc_939_nl[7:0];
  assign nl_MultLoop_acc_1009_nl = MultLoop_acc_942_nl + MultLoop_acc_941_nl + MultLoop_acc_946_nl
      + MultLoop_acc_945_nl + MultLoop_acc_944_nl + MultLoop_acc_943_nl + MultLoop_acc_940_nl
      + MultLoop_acc_939_nl;
  assign MultLoop_acc_1009_nl = nl_MultLoop_acc_1009_nl[7:0];
  assign nl_MultLoop_acc_1014_nl = MultLoop_acc_1010_nl + MultLoop_acc_1009_nl;
  assign MultLoop_acc_1014_nl = nl_MultLoop_acc_1014_nl[7:0];
  assign nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8447:8440]));
  assign MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8455:8448]));
  assign MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_938_nl = (readslicef_15_8_7(MultLoop_1056_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1057_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_938_nl = nl_MultLoop_acc_938_nl[7:0];
  assign nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8463:8456]));
  assign MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8471:8464]));
  assign MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_937_nl = (readslicef_15_8_7(MultLoop_1058_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1059_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_937_nl = nl_MultLoop_acc_937_nl[7:0];
  assign nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8479:8472]));
  assign MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8487:8480]));
  assign MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_936_nl = (readslicef_15_8_7(MultLoop_1060_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1061_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_936_nl = nl_MultLoop_acc_936_nl[7:0];
  assign nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8495:8488]));
  assign MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8503:8496]));
  assign MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_935_nl = (readslicef_15_8_7(MultLoop_1062_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1063_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_935_nl = nl_MultLoop_acc_935_nl[7:0];
  assign nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8511:8504]));
  assign MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8519:8512]));
  assign MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_934_nl = (readslicef_15_8_7(MultLoop_1064_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1065_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_934_nl = nl_MultLoop_acc_934_nl[7:0];
  assign nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8527:8520]));
  assign MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8535:8528]));
  assign MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_933_nl = (readslicef_15_8_7(MultLoop_1066_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1067_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_933_nl = nl_MultLoop_acc_933_nl[7:0];
  assign nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8543:8536]));
  assign MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8551:8544]));
  assign MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_932_nl = (readslicef_15_8_7(MultLoop_1068_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1069_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_932_nl = nl_MultLoop_acc_932_nl[7:0];
  assign nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8559:8552]));
  assign MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8567:8560]));
  assign MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_931_nl = (readslicef_15_8_7(MultLoop_1070_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1071_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_931_nl = nl_MultLoop_acc_931_nl[7:0];
  assign nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8639:8632]));
  assign MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8647:8640]));
  assign MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_926_nl = (readslicef_15_8_7(MultLoop_1080_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1081_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_926_nl = nl_MultLoop_acc_926_nl[7:0];
  assign nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8655:8648]));
  assign MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8663:8656]));
  assign MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_925_nl = (readslicef_15_8_7(MultLoop_1082_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1083_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_925_nl = nl_MultLoop_acc_925_nl[7:0];
  assign nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8671:8664]));
  assign MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8679:8672]));
  assign MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_924_nl = (readslicef_15_8_7(MultLoop_1084_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1085_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_924_nl = nl_MultLoop_acc_924_nl[7:0];
  assign nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8687:8680]));
  assign MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8695:8688]));
  assign MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_923_nl = (readslicef_15_8_7(MultLoop_1086_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1087_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_923_nl = nl_MultLoop_acc_923_nl[7:0];
  assign nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8575:8568]));
  assign MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8583:8576]));
  assign MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_930_nl = (readslicef_15_8_7(MultLoop_1072_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1073_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_930_nl = nl_MultLoop_acc_930_nl[7:0];
  assign nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8591:8584]));
  assign MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8599:8592]));
  assign MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_929_nl = (readslicef_15_8_7(MultLoop_1074_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1075_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_929_nl = nl_MultLoop_acc_929_nl[7:0];
  assign nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8607:8600]));
  assign MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8615:8608]));
  assign MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_928_nl = (readslicef_15_8_7(MultLoop_1076_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1077_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_928_nl = nl_MultLoop_acc_928_nl[7:0];
  assign nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8623:8616]));
  assign MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8631:8624]));
  assign MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_927_nl = (readslicef_15_8_7(MultLoop_1078_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1079_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_927_nl = nl_MultLoop_acc_927_nl[7:0];
  assign nl_MultLoop_acc_1013_nl = MultLoop_acc_938_nl + MultLoop_acc_937_nl + MultLoop_acc_936_nl
      + MultLoop_acc_935_nl + MultLoop_acc_934_nl + MultLoop_acc_933_nl + MultLoop_acc_932_nl
      + MultLoop_acc_931_nl + MultLoop_acc_926_nl + MultLoop_acc_925_nl + MultLoop_acc_924_nl
      + MultLoop_acc_923_nl + MultLoop_acc_930_nl + MultLoop_acc_929_nl + MultLoop_acc_928_nl
      + MultLoop_acc_927_nl;
  assign MultLoop_acc_1013_nl = nl_MultLoop_acc_1013_nl[7:0];
  assign nl_MultLoop_acc_1016_nl = MultLoop_acc_1014_nl + MultLoop_acc_1013_nl;
  assign MultLoop_acc_1016_nl = nl_MultLoop_acc_1016_nl[7:0];
  assign nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8767:8760]));
  assign MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8775:8768]));
  assign MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_918_nl = (readslicef_15_8_7(MultLoop_1096_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1097_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_918_nl = nl_MultLoop_acc_918_nl[7:0];
  assign nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8783:8776]));
  assign MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8791:8784]));
  assign MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_917_nl = (readslicef_15_8_7(MultLoop_1098_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1099_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_917_nl = nl_MultLoop_acc_917_nl[7:0];
  assign nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8895:8888]));
  assign MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8903:8896]));
  assign MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_910_nl = (readslicef_15_8_7(MultLoop_1112_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1113_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_910_nl = nl_MultLoop_acc_910_nl[7:0];
  assign nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8911:8904]));
  assign MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8919:8912]));
  assign MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_909_nl = (readslicef_15_8_7(MultLoop_1114_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1115_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_909_nl = nl_MultLoop_acc_909_nl[7:0];
  assign nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8831:8824]));
  assign MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8839:8832]));
  assign MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_914_nl = (readslicef_15_8_7(MultLoop_1104_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1105_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_914_nl = nl_MultLoop_acc_914_nl[7:0];
  assign nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8847:8840]));
  assign MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8855:8848]));
  assign MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_913_nl = (readslicef_15_8_7(MultLoop_1106_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_913_nl = nl_MultLoop_acc_913_nl[7:0];
  assign nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9151:9144]));
  assign MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9159:9152]));
  assign MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_894_nl = (readslicef_15_8_7(MultLoop_1144_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1145_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_894_nl = nl_MultLoop_acc_894_nl[7:0];
  assign nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9167:9160]));
  assign MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9175:9168]));
  assign MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_893_nl = (readslicef_15_8_7(MultLoop_1146_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1147_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_893_nl = nl_MultLoop_acc_893_nl[7:0];
  assign nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9087:9080]));
  assign MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9095:9088]));
  assign MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_898_nl = (readslicef_15_8_7(MultLoop_1136_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1137_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_898_nl = nl_MultLoop_acc_898_nl[7:0];
  assign nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9103:9096]));
  assign MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9111:9104]));
  assign MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_897_nl = (readslicef_15_8_7(MultLoop_1138_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1139_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_897_nl = nl_MultLoop_acc_897_nl[7:0];
  assign nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9119:9112]));
  assign MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9127:9120]));
  assign MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_896_nl = (readslicef_15_8_7(MultLoop_1140_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1141_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_896_nl = nl_MultLoop_acc_896_nl[7:0];
  assign nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9135:9128]));
  assign MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9143:9136]));
  assign MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_895_nl = (readslicef_15_8_7(MultLoop_1142_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1143_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_895_nl = nl_MultLoop_acc_895_nl[7:0];
  assign nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8959:8952]));
  assign MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8967:8960]));
  assign MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_906_nl = (readslicef_15_8_7(MultLoop_1120_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1121_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_906_nl = nl_MultLoop_acc_906_nl[7:0];
  assign nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8975:8968]));
  assign MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8983:8976]));
  assign MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_905_nl = (readslicef_15_8_7(MultLoop_1122_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_905_nl = nl_MultLoop_acc_905_nl[7:0];
  assign nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8991:8984]));
  assign MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8999:8992]));
  assign MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_904_nl = (readslicef_15_8_7(MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1125_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_904_nl = nl_MultLoop_acc_904_nl[7:0];
  assign nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9007:9000]));
  assign MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9015:9008]));
  assign MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_903_nl = (readslicef_15_8_7(MultLoop_1126_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1127_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_903_nl = nl_MultLoop_acc_903_nl[7:0];
  assign nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9023:9016]));
  assign MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9031:9024]));
  assign MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_902_nl = (readslicef_15_8_7(MultLoop_1128_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1129_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_902_nl = nl_MultLoop_acc_902_nl[7:0];
  assign nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9039:9032]));
  assign MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9047:9040]));
  assign MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_901_nl = (readslicef_15_8_7(MultLoop_1130_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_901_nl = nl_MultLoop_acc_901_nl[7:0];
  assign nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9055:9048]));
  assign MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9063:9056]));
  assign MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_900_nl = (readslicef_15_8_7(MultLoop_1132_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1133_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_900_nl = nl_MultLoop_acc_900_nl[7:0];
  assign nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9071:9064]));
  assign MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9079:9072]));
  assign MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_899_nl = (readslicef_15_8_7(MultLoop_1134_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1135_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_899_nl = nl_MultLoop_acc_899_nl[7:0];
  assign nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8703:8696]));
  assign MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8711:8704]));
  assign MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_922_nl = (readslicef_15_8_7(MultLoop_1088_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1089_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_922_nl = nl_MultLoop_acc_922_nl[7:0];
  assign nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8719:8712]));
  assign MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8727:8720]));
  assign MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_921_nl = (readslicef_15_8_7(MultLoop_1090_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1091_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_921_nl = nl_MultLoop_acc_921_nl[7:0];
  assign nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8735:8728]));
  assign MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8743:8736]));
  assign MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_920_nl = (readslicef_15_8_7(MultLoop_1092_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1093_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_920_nl = nl_MultLoop_acc_920_nl[7:0];
  assign nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8751:8744]));
  assign MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8759:8752]));
  assign MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_919_nl = (readslicef_15_8_7(MultLoop_1094_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1095_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_919_nl = nl_MultLoop_acc_919_nl[7:0];
  assign nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8799:8792]));
  assign MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8807:8800]));
  assign MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_916_nl = (readslicef_15_8_7(MultLoop_1100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1101_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_916_nl = nl_MultLoop_acc_916_nl[7:0];
  assign nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8815:8808]));
  assign MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8823:8816]));
  assign MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_915_nl = (readslicef_15_8_7(MultLoop_1102_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1103_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_915_nl = nl_MultLoop_acc_915_nl[7:0];
  assign nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8863:8856]));
  assign MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8871:8864]));
  assign MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_912_nl = (readslicef_15_8_7(MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1109_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_912_nl = nl_MultLoop_acc_912_nl[7:0];
  assign nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8879:8872]));
  assign MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8887:8880]));
  assign MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_911_nl = (readslicef_15_8_7(MultLoop_1110_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1111_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_911_nl = nl_MultLoop_acc_911_nl[7:0];
  assign nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8927:8920]));
  assign MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8935:8928]));
  assign MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_908_nl = (readslicef_15_8_7(MultLoop_1116_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1117_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_908_nl = nl_MultLoop_acc_908_nl[7:0];
  assign nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8943:8936]));
  assign MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8951:8944]));
  assign MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_907_nl = (readslicef_15_8_7(MultLoop_1118_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1119_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_907_nl = nl_MultLoop_acc_907_nl[7:0];
  assign nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9183:9176]));
  assign MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9191:9184]));
  assign MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_892_nl = (readslicef_15_8_7(MultLoop_1148_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1149_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_892_nl = nl_MultLoop_acc_892_nl[7:0];
  assign nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9199:9192]));
  assign MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[9207:9200]));
  assign MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_891_nl = (readslicef_15_8_7(MultLoop_1150_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1151_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_891_nl = nl_MultLoop_acc_891_nl[7:0];
  assign nl_MultLoop_acc_1015_nl = MultLoop_acc_918_nl + MultLoop_acc_917_nl + MultLoop_acc_910_nl
      + MultLoop_acc_909_nl + MultLoop_acc_914_nl + MultLoop_acc_913_nl + MultLoop_acc_894_nl
      + MultLoop_acc_893_nl + MultLoop_acc_898_nl + MultLoop_acc_897_nl + MultLoop_acc_896_nl
      + MultLoop_acc_895_nl + MultLoop_acc_906_nl + MultLoop_acc_905_nl + MultLoop_acc_904_nl
      + MultLoop_acc_903_nl + MultLoop_acc_902_nl + MultLoop_acc_901_nl + MultLoop_acc_900_nl
      + MultLoop_acc_899_nl + MultLoop_acc_922_nl + MultLoop_acc_921_nl + MultLoop_acc_920_nl
      + MultLoop_acc_919_nl + MultLoop_acc_916_nl + MultLoop_acc_915_nl + MultLoop_acc_912_nl
      + MultLoop_acc_911_nl + MultLoop_acc_908_nl + MultLoop_acc_907_nl + MultLoop_acc_892_nl
      + MultLoop_acc_891_nl;
  assign MultLoop_acc_1015_nl = nl_MultLoop_acc_1015_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1 = MultLoop_acc_1016_nl
      + MultLoop_acc_1015_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1[7:0];
  assign nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3071:3064]));
  assign MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_128_nl = (readslicef_15_8_7(MultLoop_384_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[20:14]);
  assign MultLoop_acc_128_nl = nl_MultLoop_acc_128_nl[7:0];
  assign nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[2055:2048]));
  assign MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_192_nl = MultLoop_acc_128_nl + (readslicef_15_8_7(MultLoop_257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_192_nl = nl_MultLoop_acc_192_nl[7:0];
  assign nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2063:2056]));
  assign MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2071:2064]));
  assign MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_191_nl = (readslicef_15_8_7(MultLoop_258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_191_nl = nl_MultLoop_acc_191_nl[7:0];
  assign nl_MultLoop_acc_224_nl = MultLoop_acc_192_nl + MultLoop_acc_191_nl;
  assign MultLoop_acc_224_nl = nl_MultLoop_acc_224_nl[7:0];
  assign nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2079:2072]));
  assign MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2087:2080]));
  assign MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_190_nl = (readslicef_15_8_7(MultLoop_260_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_261_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_190_nl = nl_MultLoop_acc_190_nl[7:0];
  assign nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2095:2088]));
  assign MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2103:2096]));
  assign MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_189_nl = (readslicef_15_8_7(MultLoop_262_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_263_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_189_nl = nl_MultLoop_acc_189_nl[7:0];
  assign nl_MultLoop_acc_223_nl = MultLoop_acc_190_nl + MultLoop_acc_189_nl;
  assign MultLoop_acc_223_nl = nl_MultLoop_acc_223_nl[7:0];
  assign nl_MultLoop_acc_240_nl = MultLoop_acc_224_nl + MultLoop_acc_223_nl;
  assign MultLoop_acc_240_nl = nl_MultLoop_acc_240_nl[7:0];
  assign nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2111:2104]));
  assign MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2119:2112]));
  assign MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_188_nl = (readslicef_15_8_7(MultLoop_264_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_265_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_188_nl = nl_MultLoop_acc_188_nl[7:0];
  assign nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2127:2120]));
  assign MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2135:2128]));
  assign MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_187_nl = (readslicef_15_8_7(MultLoop_266_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_267_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_187_nl = nl_MultLoop_acc_187_nl[7:0];
  assign nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2143:2136]));
  assign MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2151:2144]));
  assign MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_186_nl = (readslicef_15_8_7(MultLoop_268_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_269_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_186_nl = nl_MultLoop_acc_186_nl[7:0];
  assign nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2159:2152]));
  assign MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2167:2160]));
  assign MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_185_nl = (readslicef_15_8_7(MultLoop_270_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_271_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_185_nl = nl_MultLoop_acc_185_nl[7:0];
  assign nl_MultLoop_acc_239_nl = MultLoop_acc_188_nl + MultLoop_acc_187_nl + MultLoop_acc_186_nl
      + MultLoop_acc_185_nl;
  assign MultLoop_acc_239_nl = nl_MultLoop_acc_239_nl[7:0];
  assign nl_MultLoop_acc_248_nl = MultLoop_acc_240_nl + MultLoop_acc_239_nl;
  assign MultLoop_acc_248_nl = nl_MultLoop_acc_248_nl[7:0];
  assign nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2239:2232]));
  assign MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2247:2240]));
  assign MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_180_nl = (readslicef_15_8_7(MultLoop_280_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_281_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_180_nl = nl_MultLoop_acc_180_nl[7:0];
  assign nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2255:2248]));
  assign MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2263:2256]));
  assign MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_179_nl = (readslicef_15_8_7(MultLoop_282_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_283_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_179_nl = nl_MultLoop_acc_179_nl[7:0];
  assign nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2175:2168]));
  assign MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2183:2176]));
  assign MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_184_nl = (readslicef_15_8_7(MultLoop_272_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_273_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_184_nl = nl_MultLoop_acc_184_nl[7:0];
  assign nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2191:2184]));
  assign MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2199:2192]));
  assign MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_183_nl = (readslicef_15_8_7(MultLoop_274_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_275_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_183_nl = nl_MultLoop_acc_183_nl[7:0];
  assign nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2207:2200]));
  assign MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2215:2208]));
  assign MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_182_nl = (readslicef_15_8_7(MultLoop_276_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_277_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_182_nl = nl_MultLoop_acc_182_nl[7:0];
  assign nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2223:2216]));
  assign MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2231:2224]));
  assign MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_181_nl = (readslicef_15_8_7(MultLoop_278_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_279_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_181_nl = nl_MultLoop_acc_181_nl[7:0];
  assign nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2271:2264]));
  assign MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2279:2272]));
  assign MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_178_nl = (readslicef_15_8_7(MultLoop_284_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_285_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_178_nl = nl_MultLoop_acc_178_nl[7:0];
  assign nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2287:2280]));
  assign MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2295:2288]));
  assign MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_177_nl = (readslicef_15_8_7(MultLoop_286_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_287_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_177_nl = nl_MultLoop_acc_177_nl[7:0];
  assign nl_MultLoop_acc_247_nl = MultLoop_acc_180_nl + MultLoop_acc_179_nl + MultLoop_acc_184_nl
      + MultLoop_acc_183_nl + MultLoop_acc_182_nl + MultLoop_acc_181_nl + MultLoop_acc_178_nl
      + MultLoop_acc_177_nl;
  assign MultLoop_acc_247_nl = nl_MultLoop_acc_247_nl[7:0];
  assign nl_MultLoop_acc_252_nl = MultLoop_acc_248_nl + MultLoop_acc_247_nl;
  assign MultLoop_acc_252_nl = nl_MultLoop_acc_252_nl[7:0];
  assign nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2303:2296]));
  assign MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2311:2304]));
  assign MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_176_nl = (readslicef_15_8_7(MultLoop_288_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_289_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_176_nl = nl_MultLoop_acc_176_nl[7:0];
  assign nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2319:2312]));
  assign MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2327:2320]));
  assign MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_175_nl = (readslicef_15_8_7(MultLoop_290_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_291_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_175_nl = nl_MultLoop_acc_175_nl[7:0];
  assign nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2335:2328]));
  assign MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2343:2336]));
  assign MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_174_nl = (readslicef_15_8_7(MultLoop_292_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_293_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_174_nl = nl_MultLoop_acc_174_nl[7:0];
  assign nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2351:2344]));
  assign MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2359:2352]));
  assign MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_173_nl = (readslicef_15_8_7(MultLoop_294_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_295_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_173_nl = nl_MultLoop_acc_173_nl[7:0];
  assign nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2367:2360]));
  assign MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2375:2368]));
  assign MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_172_nl = (readslicef_15_8_7(MultLoop_296_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_297_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_172_nl = nl_MultLoop_acc_172_nl[7:0];
  assign nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2383:2376]));
  assign MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2391:2384]));
  assign MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_171_nl = (readslicef_15_8_7(MultLoop_298_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_299_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_171_nl = nl_MultLoop_acc_171_nl[7:0];
  assign nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2399:2392]));
  assign MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2407:2400]));
  assign MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_170_nl = (readslicef_15_8_7(MultLoop_300_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_301_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_170_nl = nl_MultLoop_acc_170_nl[7:0];
  assign nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2415:2408]));
  assign MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2423:2416]));
  assign MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_169_nl = (readslicef_15_8_7(MultLoop_302_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_303_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_169_nl = nl_MultLoop_acc_169_nl[7:0];
  assign nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2495:2488]));
  assign MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2503:2496]));
  assign MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_164_nl = (readslicef_15_8_7(MultLoop_312_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_313_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_164_nl = nl_MultLoop_acc_164_nl[7:0];
  assign nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2511:2504]));
  assign MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2519:2512]));
  assign MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_163_nl = (readslicef_15_8_7(MultLoop_314_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_315_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_163_nl = nl_MultLoop_acc_163_nl[7:0];
  assign nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2527:2520]));
  assign MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2535:2528]));
  assign MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_162_nl = (readslicef_15_8_7(MultLoop_316_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_317_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_162_nl = nl_MultLoop_acc_162_nl[7:0];
  assign nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2543:2536]));
  assign MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2551:2544]));
  assign MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_161_nl = (readslicef_15_8_7(MultLoop_318_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_319_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_161_nl = nl_MultLoop_acc_161_nl[7:0];
  assign nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2431:2424]));
  assign MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2439:2432]));
  assign MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_168_nl = (readslicef_15_8_7(MultLoop_304_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_305_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_168_nl = nl_MultLoop_acc_168_nl[7:0];
  assign nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2447:2440]));
  assign MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2455:2448]));
  assign MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_167_nl = (readslicef_15_8_7(MultLoop_306_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_307_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_167_nl = nl_MultLoop_acc_167_nl[7:0];
  assign nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2463:2456]));
  assign MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2471:2464]));
  assign MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_166_nl = (readslicef_15_8_7(MultLoop_308_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_309_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_166_nl = nl_MultLoop_acc_166_nl[7:0];
  assign nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2479:2472]));
  assign MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2487:2480]));
  assign MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_165_nl = (readslicef_15_8_7(MultLoop_310_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_311_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[7:0];
  assign nl_MultLoop_acc_251_nl = MultLoop_acc_176_nl + MultLoop_acc_175_nl + MultLoop_acc_174_nl
      + MultLoop_acc_173_nl + MultLoop_acc_172_nl + MultLoop_acc_171_nl + MultLoop_acc_170_nl
      + MultLoop_acc_169_nl + MultLoop_acc_164_nl + MultLoop_acc_163_nl + MultLoop_acc_162_nl
      + MultLoop_acc_161_nl + MultLoop_acc_168_nl + MultLoop_acc_167_nl + MultLoop_acc_166_nl
      + MultLoop_acc_165_nl;
  assign MultLoop_acc_251_nl = nl_MultLoop_acc_251_nl[7:0];
  assign nl_MultLoop_acc_254_nl = MultLoop_acc_252_nl + MultLoop_acc_251_nl;
  assign MultLoop_acc_254_nl = nl_MultLoop_acc_254_nl[7:0];
  assign nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2623:2616]));
  assign MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2631:2624]));
  assign MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_156_nl = (readslicef_15_8_7(MultLoop_328_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_329_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_156_nl = nl_MultLoop_acc_156_nl[7:0];
  assign nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2639:2632]));
  assign MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2647:2640]));
  assign MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_155_nl = (readslicef_15_8_7(MultLoop_330_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_331_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_155_nl = nl_MultLoop_acc_155_nl[7:0];
  assign nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2751:2744]));
  assign MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2759:2752]));
  assign MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_148_nl = (readslicef_15_8_7(MultLoop_344_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_345_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_148_nl = nl_MultLoop_acc_148_nl[7:0];
  assign nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2767:2760]));
  assign MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2775:2768]));
  assign MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_147_nl = (readslicef_15_8_7(MultLoop_346_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_347_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_147_nl = nl_MultLoop_acc_147_nl[7:0];
  assign nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2687:2680]));
  assign MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2695:2688]));
  assign MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_152_nl = (readslicef_15_8_7(MultLoop_336_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_337_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_152_nl = nl_MultLoop_acc_152_nl[7:0];
  assign nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2703:2696]));
  assign MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2711:2704]));
  assign MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_151_nl = (readslicef_15_8_7(MultLoop_338_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_339_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_151_nl = nl_MultLoop_acc_151_nl[7:0];
  assign nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3007:3000]));
  assign MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3015:3008]));
  assign MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_132_nl = (readslicef_15_8_7(MultLoop_376_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_377_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_132_nl = nl_MultLoop_acc_132_nl[7:0];
  assign nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3023:3016]));
  assign MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3031:3024]));
  assign MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_131_nl = (readslicef_15_8_7(MultLoop_378_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_379_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_131_nl = nl_MultLoop_acc_131_nl[7:0];
  assign nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2943:2936]));
  assign MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2951:2944]));
  assign MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_136_nl = (readslicef_15_8_7(MultLoop_368_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_369_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_136_nl = nl_MultLoop_acc_136_nl[7:0];
  assign nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2959:2952]));
  assign MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2967:2960]));
  assign MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_135_nl = (readslicef_15_8_7(MultLoop_370_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_371_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_135_nl = nl_MultLoop_acc_135_nl[7:0];
  assign nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2975:2968]));
  assign MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2983:2976]));
  assign MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_134_nl = (readslicef_15_8_7(MultLoop_372_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_373_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[7:0];
  assign nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2991:2984]));
  assign MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2999:2992]));
  assign MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_133_nl = (readslicef_15_8_7(MultLoop_374_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_375_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_133_nl = nl_MultLoop_acc_133_nl[7:0];
  assign nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2815:2808]));
  assign MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2823:2816]));
  assign MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_144_nl = (readslicef_15_8_7(MultLoop_352_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_353_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_144_nl = nl_MultLoop_acc_144_nl[7:0];
  assign nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2831:2824]));
  assign MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2839:2832]));
  assign MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_143_nl = (readslicef_15_8_7(MultLoop_354_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[7:0];
  assign nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2847:2840]));
  assign MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2855:2848]));
  assign MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_142_nl = (readslicef_15_8_7(MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_357_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_142_nl = nl_MultLoop_acc_142_nl[7:0];
  assign nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2863:2856]));
  assign MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2871:2864]));
  assign MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_141_nl = (readslicef_15_8_7(MultLoop_358_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_359_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_141_nl = nl_MultLoop_acc_141_nl[7:0];
  assign nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2879:2872]));
  assign MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2887:2880]));
  assign MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_140_nl = (readslicef_15_8_7(MultLoop_360_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_361_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_140_nl = nl_MultLoop_acc_140_nl[7:0];
  assign nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2895:2888]));
  assign MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2903:2896]));
  assign MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_139_nl = (readslicef_15_8_7(MultLoop_362_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_363_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_139_nl = nl_MultLoop_acc_139_nl[7:0];
  assign nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2911:2904]));
  assign MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2919:2912]));
  assign MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_138_nl = (readslicef_15_8_7(MultLoop_364_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_365_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_138_nl = nl_MultLoop_acc_138_nl[7:0];
  assign nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2927:2920]));
  assign MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2935:2928]));
  assign MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_137_nl = (readslicef_15_8_7(MultLoop_366_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_367_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_137_nl = nl_MultLoop_acc_137_nl[7:0];
  assign nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2559:2552]));
  assign MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2567:2560]));
  assign MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_160_nl = (readslicef_15_8_7(MultLoop_320_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_160_nl = nl_MultLoop_acc_160_nl[7:0];
  assign nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2575:2568]));
  assign MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2583:2576]));
  assign MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_159_nl = (readslicef_15_8_7(MultLoop_322_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_323_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[7:0];
  assign nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2591:2584]));
  assign MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2599:2592]));
  assign MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_158_nl = (readslicef_15_8_7(MultLoop_324_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_325_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[7:0];
  assign nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2607:2600]));
  assign MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2615:2608]));
  assign MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_157_nl = (readslicef_15_8_7(MultLoop_326_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_327_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_157_nl = nl_MultLoop_acc_157_nl[7:0];
  assign nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2655:2648]));
  assign MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2663:2656]));
  assign MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_154_nl = (readslicef_15_8_7(MultLoop_332_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_333_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_154_nl = nl_MultLoop_acc_154_nl[7:0];
  assign nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2671:2664]));
  assign MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2679:2672]));
  assign MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_153_nl = (readslicef_15_8_7(MultLoop_334_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_335_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_153_nl = nl_MultLoop_acc_153_nl[7:0];
  assign nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2719:2712]));
  assign MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2727:2720]));
  assign MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_150_nl = (readslicef_15_8_7(MultLoop_340_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_341_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_150_nl = nl_MultLoop_acc_150_nl[7:0];
  assign nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2735:2728]));
  assign MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2743:2736]));
  assign MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_149_nl = (readslicef_15_8_7(MultLoop_342_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_343_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_149_nl = nl_MultLoop_acc_149_nl[7:0];
  assign nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2783:2776]));
  assign MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2791:2784]));
  assign MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_146_nl = (readslicef_15_8_7(MultLoop_348_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_349_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_146_nl = nl_MultLoop_acc_146_nl[7:0];
  assign nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2799:2792]));
  assign MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[2807:2800]));
  assign MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_145_nl = (readslicef_15_8_7(MultLoop_350_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_351_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_145_nl = nl_MultLoop_acc_145_nl[7:0];
  assign nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3039:3032]));
  assign MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3047:3040]));
  assign MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_130_nl = (readslicef_15_8_7(MultLoop_380_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_381_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_130_nl = nl_MultLoop_acc_130_nl[7:0];
  assign nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3055:3048]));
  assign MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3063:3056]));
  assign MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_129_nl = (readslicef_15_8_7(MultLoop_382_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_383_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_129_nl = nl_MultLoop_acc_129_nl[7:0];
  assign nl_MultLoop_acc_253_nl = MultLoop_acc_156_nl + MultLoop_acc_155_nl + MultLoop_acc_148_nl
      + MultLoop_acc_147_nl + MultLoop_acc_152_nl + MultLoop_acc_151_nl + MultLoop_acc_132_nl
      + MultLoop_acc_131_nl + MultLoop_acc_136_nl + MultLoop_acc_135_nl + MultLoop_acc_134_nl
      + MultLoop_acc_133_nl + MultLoop_acc_144_nl + MultLoop_acc_143_nl + MultLoop_acc_142_nl
      + MultLoop_acc_141_nl + MultLoop_acc_140_nl + MultLoop_acc_139_nl + MultLoop_acc_138_nl
      + MultLoop_acc_137_nl + MultLoop_acc_160_nl + MultLoop_acc_159_nl + MultLoop_acc_158_nl
      + MultLoop_acc_157_nl + MultLoop_acc_154_nl + MultLoop_acc_153_nl + MultLoop_acc_150_nl
      + MultLoop_acc_149_nl + MultLoop_acc_146_nl + MultLoop_acc_145_nl + MultLoop_acc_130_nl
      + MultLoop_acc_129_nl;
  assign MultLoop_acc_253_nl = nl_MultLoop_acc_253_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1 = MultLoop_acc_254_nl
      + MultLoop_acc_253_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1[7:0];
  assign nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8191:8184]));
  assign MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_763_nl = (readslicef_15_8_7(MultLoop_1024_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[55:49]);
  assign MultLoop_acc_763_nl = nl_MultLoop_acc_763_nl[7:0];
  assign nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[7175:7168]));
  assign MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_827_nl = MultLoop_acc_763_nl + (readslicef_15_8_7(MultLoop_897_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_827_nl = nl_MultLoop_acc_827_nl[7:0];
  assign nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7183:7176]));
  assign MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7191:7184]));
  assign MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_826_nl = (readslicef_15_8_7(MultLoop_898_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_899_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_826_nl = nl_MultLoop_acc_826_nl[7:0];
  assign nl_MultLoop_acc_859_nl = MultLoop_acc_827_nl + MultLoop_acc_826_nl;
  assign MultLoop_acc_859_nl = nl_MultLoop_acc_859_nl[7:0];
  assign nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7199:7192]));
  assign MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7207:7200]));
  assign MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_825_nl = (readslicef_15_8_7(MultLoop_900_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_901_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_825_nl = nl_MultLoop_acc_825_nl[7:0];
  assign nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7215:7208]));
  assign MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7223:7216]));
  assign MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_824_nl = (readslicef_15_8_7(MultLoop_902_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_903_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_824_nl = nl_MultLoop_acc_824_nl[7:0];
  assign nl_MultLoop_acc_858_nl = MultLoop_acc_825_nl + MultLoop_acc_824_nl;
  assign MultLoop_acc_858_nl = nl_MultLoop_acc_858_nl[7:0];
  assign nl_MultLoop_acc_875_nl = MultLoop_acc_859_nl + MultLoop_acc_858_nl;
  assign MultLoop_acc_875_nl = nl_MultLoop_acc_875_nl[7:0];
  assign nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7231:7224]));
  assign MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7239:7232]));
  assign MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_823_nl = (readslicef_15_8_7(MultLoop_904_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_905_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_823_nl = nl_MultLoop_acc_823_nl[7:0];
  assign nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7247:7240]));
  assign MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7255:7248]));
  assign MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_822_nl = (readslicef_15_8_7(MultLoop_906_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_907_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_822_nl = nl_MultLoop_acc_822_nl[7:0];
  assign nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7263:7256]));
  assign MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7271:7264]));
  assign MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_821_nl = (readslicef_15_8_7(MultLoop_908_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_909_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_821_nl = nl_MultLoop_acc_821_nl[7:0];
  assign nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7279:7272]));
  assign MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7287:7280]));
  assign MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_820_nl = (readslicef_15_8_7(MultLoop_910_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_911_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_820_nl = nl_MultLoop_acc_820_nl[7:0];
  assign nl_MultLoop_acc_874_nl = MultLoop_acc_823_nl + MultLoop_acc_822_nl + MultLoop_acc_821_nl
      + MultLoop_acc_820_nl;
  assign MultLoop_acc_874_nl = nl_MultLoop_acc_874_nl[7:0];
  assign nl_MultLoop_acc_883_nl = MultLoop_acc_875_nl + MultLoop_acc_874_nl;
  assign MultLoop_acc_883_nl = nl_MultLoop_acc_883_nl[7:0];
  assign nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7359:7352]));
  assign MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7367:7360]));
  assign MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_815_nl = (readslicef_15_8_7(MultLoop_920_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_921_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_815_nl = nl_MultLoop_acc_815_nl[7:0];
  assign nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7375:7368]));
  assign MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7383:7376]));
  assign MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_814_nl = (readslicef_15_8_7(MultLoop_922_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_923_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_814_nl = nl_MultLoop_acc_814_nl[7:0];
  assign nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7295:7288]));
  assign MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7303:7296]));
  assign MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_819_nl = (readslicef_15_8_7(MultLoop_912_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_913_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_819_nl = nl_MultLoop_acc_819_nl[7:0];
  assign nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7311:7304]));
  assign MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7319:7312]));
  assign MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_818_nl = (readslicef_15_8_7(MultLoop_914_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_915_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_818_nl = nl_MultLoop_acc_818_nl[7:0];
  assign nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7327:7320]));
  assign MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7335:7328]));
  assign MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_817_nl = (readslicef_15_8_7(MultLoop_916_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_917_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_817_nl = nl_MultLoop_acc_817_nl[7:0];
  assign nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7343:7336]));
  assign MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7351:7344]));
  assign MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_816_nl = (readslicef_15_8_7(MultLoop_918_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_919_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_816_nl = nl_MultLoop_acc_816_nl[7:0];
  assign nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7391:7384]));
  assign MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7399:7392]));
  assign MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_813_nl = (readslicef_15_8_7(MultLoop_924_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_925_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_813_nl = nl_MultLoop_acc_813_nl[7:0];
  assign nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7407:7400]));
  assign MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7415:7408]));
  assign MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_812_nl = (readslicef_15_8_7(MultLoop_926_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_927_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_812_nl = nl_MultLoop_acc_812_nl[7:0];
  assign nl_MultLoop_acc_882_nl = MultLoop_acc_815_nl + MultLoop_acc_814_nl + MultLoop_acc_819_nl
      + MultLoop_acc_818_nl + MultLoop_acc_817_nl + MultLoop_acc_816_nl + MultLoop_acc_813_nl
      + MultLoop_acc_812_nl;
  assign MultLoop_acc_882_nl = nl_MultLoop_acc_882_nl[7:0];
  assign nl_MultLoop_acc_887_nl = MultLoop_acc_883_nl + MultLoop_acc_882_nl;
  assign MultLoop_acc_887_nl = nl_MultLoop_acc_887_nl[7:0];
  assign nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7423:7416]));
  assign MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7431:7424]));
  assign MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_811_nl = (readslicef_15_8_7(MultLoop_928_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_929_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_811_nl = nl_MultLoop_acc_811_nl[7:0];
  assign nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7439:7432]));
  assign MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7447:7440]));
  assign MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_810_nl = (readslicef_15_8_7(MultLoop_930_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_931_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_810_nl = nl_MultLoop_acc_810_nl[7:0];
  assign nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7455:7448]));
  assign MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7463:7456]));
  assign MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_809_nl = (readslicef_15_8_7(MultLoop_932_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_933_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_809_nl = nl_MultLoop_acc_809_nl[7:0];
  assign nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7471:7464]));
  assign MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7479:7472]));
  assign MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_808_nl = (readslicef_15_8_7(MultLoop_934_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_935_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_808_nl = nl_MultLoop_acc_808_nl[7:0];
  assign nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7487:7480]));
  assign MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7495:7488]));
  assign MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_807_nl = (readslicef_15_8_7(MultLoop_936_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_937_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_807_nl = nl_MultLoop_acc_807_nl[7:0];
  assign nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7503:7496]));
  assign MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7511:7504]));
  assign MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_806_nl = (readslicef_15_8_7(MultLoop_938_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_939_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_806_nl = nl_MultLoop_acc_806_nl[7:0];
  assign nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7519:7512]));
  assign MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7527:7520]));
  assign MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_805_nl = (readslicef_15_8_7(MultLoop_940_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_941_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_805_nl = nl_MultLoop_acc_805_nl[7:0];
  assign nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7535:7528]));
  assign MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7543:7536]));
  assign MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_804_nl = (readslicef_15_8_7(MultLoop_942_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_943_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_804_nl = nl_MultLoop_acc_804_nl[7:0];
  assign nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7615:7608]));
  assign MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7623:7616]));
  assign MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_799_nl = (readslicef_15_8_7(MultLoop_952_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_953_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_799_nl = nl_MultLoop_acc_799_nl[7:0];
  assign nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7631:7624]));
  assign MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7639:7632]));
  assign MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_798_nl = (readslicef_15_8_7(MultLoop_954_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_955_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_798_nl = nl_MultLoop_acc_798_nl[7:0];
  assign nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7647:7640]));
  assign MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7655:7648]));
  assign MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_797_nl = (readslicef_15_8_7(MultLoop_956_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_957_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_797_nl = nl_MultLoop_acc_797_nl[7:0];
  assign nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7663:7656]));
  assign MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7671:7664]));
  assign MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_796_nl = (readslicef_15_8_7(MultLoop_958_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_959_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_796_nl = nl_MultLoop_acc_796_nl[7:0];
  assign nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7551:7544]));
  assign MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7559:7552]));
  assign MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_803_nl = (readslicef_15_8_7(MultLoop_944_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_945_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_803_nl = nl_MultLoop_acc_803_nl[7:0];
  assign nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7567:7560]));
  assign MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7575:7568]));
  assign MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_802_nl = (readslicef_15_8_7(MultLoop_946_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_947_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_802_nl = nl_MultLoop_acc_802_nl[7:0];
  assign nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7583:7576]));
  assign MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7591:7584]));
  assign MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_801_nl = (readslicef_15_8_7(MultLoop_948_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_949_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_801_nl = nl_MultLoop_acc_801_nl[7:0];
  assign nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7599:7592]));
  assign MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7607:7600]));
  assign MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_800_nl = (readslicef_15_8_7(MultLoop_950_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_951_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_800_nl = nl_MultLoop_acc_800_nl[7:0];
  assign nl_MultLoop_acc_886_nl = MultLoop_acc_811_nl + MultLoop_acc_810_nl + MultLoop_acc_809_nl
      + MultLoop_acc_808_nl + MultLoop_acc_807_nl + MultLoop_acc_806_nl + MultLoop_acc_805_nl
      + MultLoop_acc_804_nl + MultLoop_acc_799_nl + MultLoop_acc_798_nl + MultLoop_acc_797_nl
      + MultLoop_acc_796_nl + MultLoop_acc_803_nl + MultLoop_acc_802_nl + MultLoop_acc_801_nl
      + MultLoop_acc_800_nl;
  assign MultLoop_acc_886_nl = nl_MultLoop_acc_886_nl[7:0];
  assign nl_MultLoop_acc_889_nl = MultLoop_acc_887_nl + MultLoop_acc_886_nl;
  assign MultLoop_acc_889_nl = nl_MultLoop_acc_889_nl[7:0];
  assign nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7743:7736]));
  assign MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7751:7744]));
  assign MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_791_nl = (readslicef_15_8_7(MultLoop_968_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_969_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_791_nl = nl_MultLoop_acc_791_nl[7:0];
  assign nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7759:7752]));
  assign MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7767:7760]));
  assign MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_790_nl = (readslicef_15_8_7(MultLoop_970_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_971_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_790_nl = nl_MultLoop_acc_790_nl[7:0];
  assign nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7871:7864]));
  assign MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7879:7872]));
  assign MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_783_nl = (readslicef_15_8_7(MultLoop_984_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_985_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_783_nl = nl_MultLoop_acc_783_nl[7:0];
  assign nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7887:7880]));
  assign MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7895:7888]));
  assign MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_782_nl = (readslicef_15_8_7(MultLoop_986_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_987_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_782_nl = nl_MultLoop_acc_782_nl[7:0];
  assign nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7807:7800]));
  assign MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7815:7808]));
  assign MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_787_nl = (readslicef_15_8_7(MultLoop_976_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_977_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_787_nl = nl_MultLoop_acc_787_nl[7:0];
  assign nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7823:7816]));
  assign MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7831:7824]));
  assign MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_786_nl = (readslicef_15_8_7(MultLoop_978_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_979_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_786_nl = nl_MultLoop_acc_786_nl[7:0];
  assign nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8127:8120]));
  assign MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8135:8128]));
  assign MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_767_nl = (readslicef_15_8_7(MultLoop_1016_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1017_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_767_nl = nl_MultLoop_acc_767_nl[7:0];
  assign nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8143:8136]));
  assign MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8151:8144]));
  assign MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_766_nl = (readslicef_15_8_7(MultLoop_1018_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_766_nl = nl_MultLoop_acc_766_nl[7:0];
  assign nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8063:8056]));
  assign MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8071:8064]));
  assign MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_771_nl = (readslicef_15_8_7(MultLoop_1008_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1009_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_771_nl = nl_MultLoop_acc_771_nl[7:0];
  assign nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8079:8072]));
  assign MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8087:8080]));
  assign MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_770_nl = (readslicef_15_8_7(MultLoop_1010_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1011_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_770_nl = nl_MultLoop_acc_770_nl[7:0];
  assign nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8095:8088]));
  assign MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8103:8096]));
  assign MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_769_nl = (readslicef_15_8_7(MultLoop_1012_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1013_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_769_nl = nl_MultLoop_acc_769_nl[7:0];
  assign nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8111:8104]));
  assign MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8119:8112]));
  assign MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_768_nl = (readslicef_15_8_7(MultLoop_1014_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1015_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_768_nl = nl_MultLoop_acc_768_nl[7:0];
  assign nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7935:7928]));
  assign MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7943:7936]));
  assign MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_779_nl = (readslicef_15_8_7(MultLoop_992_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_993_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_779_nl = nl_MultLoop_acc_779_nl[7:0];
  assign nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7951:7944]));
  assign MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7959:7952]));
  assign MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_778_nl = (readslicef_15_8_7(MultLoop_994_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_778_nl = nl_MultLoop_acc_778_nl[7:0];
  assign nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7967:7960]));
  assign MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7975:7968]));
  assign MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_777_nl = (readslicef_15_8_7(MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_997_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_777_nl = nl_MultLoop_acc_777_nl[7:0];
  assign nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7983:7976]));
  assign MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7991:7984]));
  assign MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_776_nl = (readslicef_15_8_7(MultLoop_998_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_999_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_776_nl = nl_MultLoop_acc_776_nl[7:0];
  assign nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7999:7992]));
  assign MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8007:8000]));
  assign MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_775_nl = (readslicef_15_8_7(MultLoop_1000_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1001_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_775_nl = nl_MultLoop_acc_775_nl[7:0];
  assign nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8015:8008]));
  assign MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8023:8016]));
  assign MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_774_nl = (readslicef_15_8_7(MultLoop_1002_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1003_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_774_nl = nl_MultLoop_acc_774_nl[7:0];
  assign nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8031:8024]));
  assign MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8039:8032]));
  assign MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_773_nl = (readslicef_15_8_7(MultLoop_1004_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1005_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_773_nl = nl_MultLoop_acc_773_nl[7:0];
  assign nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8047:8040]));
  assign MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8055:8048]));
  assign MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_772_nl = (readslicef_15_8_7(MultLoop_1006_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1007_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_772_nl = nl_MultLoop_acc_772_nl[7:0];
  assign nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7679:7672]));
  assign MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7687:7680]));
  assign MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_795_nl = (readslicef_15_8_7(MultLoop_960_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_795_nl = nl_MultLoop_acc_795_nl[7:0];
  assign nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7695:7688]));
  assign MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7703:7696]));
  assign MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_794_nl = (readslicef_15_8_7(MultLoop_962_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_963_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_794_nl = nl_MultLoop_acc_794_nl[7:0];
  assign nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7711:7704]));
  assign MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7719:7712]));
  assign MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_793_nl = (readslicef_15_8_7(MultLoop_964_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_965_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_793_nl = nl_MultLoop_acc_793_nl[7:0];
  assign nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7727:7720]));
  assign MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7735:7728]));
  assign MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_792_nl = (readslicef_15_8_7(MultLoop_966_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_967_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_792_nl = nl_MultLoop_acc_792_nl[7:0];
  assign nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7775:7768]));
  assign MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7783:7776]));
  assign MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_789_nl = (readslicef_15_8_7(MultLoop_972_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_973_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_789_nl = nl_MultLoop_acc_789_nl[7:0];
  assign nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7791:7784]));
  assign MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7799:7792]));
  assign MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_788_nl = (readslicef_15_8_7(MultLoop_974_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_975_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_788_nl = nl_MultLoop_acc_788_nl[7:0];
  assign nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7839:7832]));
  assign MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7847:7840]));
  assign MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_785_nl = (readslicef_15_8_7(MultLoop_980_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_981_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_785_nl = nl_MultLoop_acc_785_nl[7:0];
  assign nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7855:7848]));
  assign MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7863:7856]));
  assign MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_784_nl = (readslicef_15_8_7(MultLoop_982_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_983_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_784_nl = nl_MultLoop_acc_784_nl[7:0];
  assign nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7903:7896]));
  assign MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7911:7904]));
  assign MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_781_nl = (readslicef_15_8_7(MultLoop_988_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_989_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_781_nl = nl_MultLoop_acc_781_nl[7:0];
  assign nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7919:7912]));
  assign MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7927:7920]));
  assign MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_780_nl = (readslicef_15_8_7(MultLoop_990_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_991_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_780_nl = nl_MultLoop_acc_780_nl[7:0];
  assign nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8159:8152]));
  assign MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8167:8160]));
  assign MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_765_nl = (readslicef_15_8_7(MultLoop_1020_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1021_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_765_nl = nl_MultLoop_acc_765_nl[7:0];
  assign nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8175:8168]));
  assign MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[8183:8176]));
  assign MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_764_nl = (readslicef_15_8_7(MultLoop_1022_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_1023_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_764_nl = nl_MultLoop_acc_764_nl[7:0];
  assign nl_MultLoop_acc_888_nl = MultLoop_acc_791_nl + MultLoop_acc_790_nl + MultLoop_acc_783_nl
      + MultLoop_acc_782_nl + MultLoop_acc_787_nl + MultLoop_acc_786_nl + MultLoop_acc_767_nl
      + MultLoop_acc_766_nl + MultLoop_acc_771_nl + MultLoop_acc_770_nl + MultLoop_acc_769_nl
      + MultLoop_acc_768_nl + MultLoop_acc_779_nl + MultLoop_acc_778_nl + MultLoop_acc_777_nl
      + MultLoop_acc_776_nl + MultLoop_acc_775_nl + MultLoop_acc_774_nl + MultLoop_acc_773_nl
      + MultLoop_acc_772_nl + MultLoop_acc_795_nl + MultLoop_acc_794_nl + MultLoop_acc_793_nl
      + MultLoop_acc_792_nl + MultLoop_acc_789_nl + MultLoop_acc_788_nl + MultLoop_acc_785_nl
      + MultLoop_acc_784_nl + MultLoop_acc_781_nl + MultLoop_acc_780_nl + MultLoop_acc_765_nl
      + MultLoop_acc_764_nl;
  assign MultLoop_acc_888_nl = nl_MultLoop_acc_888_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1 = MultLoop_acc_889_nl
      + MultLoop_acc_888_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1[7:0];
  assign nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4095:4088]));
  assign MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_255_nl = (readslicef_15_8_7(MultLoop_512_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[27:21]);
  assign MultLoop_acc_255_nl = nl_MultLoop_acc_255_nl[7:0];
  assign nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[3079:3072]));
  assign MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_319_nl = MultLoop_acc_255_nl + (readslicef_15_8_7(MultLoop_385_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_319_nl = nl_MultLoop_acc_319_nl[7:0];
  assign nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3087:3080]));
  assign MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3095:3088]));
  assign MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_318_nl = (readslicef_15_8_7(MultLoop_386_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_387_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_318_nl = nl_MultLoop_acc_318_nl[7:0];
  assign nl_MultLoop_acc_351_nl = MultLoop_acc_319_nl + MultLoop_acc_318_nl;
  assign MultLoop_acc_351_nl = nl_MultLoop_acc_351_nl[7:0];
  assign nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3103:3096]));
  assign MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3111:3104]));
  assign MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_317_nl = (readslicef_15_8_7(MultLoop_388_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_389_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_317_nl = nl_MultLoop_acc_317_nl[7:0];
  assign nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3119:3112]));
  assign MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3127:3120]));
  assign MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_316_nl = (readslicef_15_8_7(MultLoop_390_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_316_nl = nl_MultLoop_acc_316_nl[7:0];
  assign nl_MultLoop_acc_350_nl = MultLoop_acc_317_nl + MultLoop_acc_316_nl;
  assign MultLoop_acc_350_nl = nl_MultLoop_acc_350_nl[7:0];
  assign nl_MultLoop_acc_367_nl = MultLoop_acc_351_nl + MultLoop_acc_350_nl;
  assign MultLoop_acc_367_nl = nl_MultLoop_acc_367_nl[7:0];
  assign nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3135:3128]));
  assign MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3143:3136]));
  assign MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_315_nl = (readslicef_15_8_7(MultLoop_392_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_393_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_315_nl = nl_MultLoop_acc_315_nl[7:0];
  assign nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3151:3144]));
  assign MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3159:3152]));
  assign MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_314_nl = (readslicef_15_8_7(MultLoop_394_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_395_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_314_nl = nl_MultLoop_acc_314_nl[7:0];
  assign nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3167:3160]));
  assign MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3175:3168]));
  assign MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_313_nl = (readslicef_15_8_7(MultLoop_396_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_397_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_313_nl = nl_MultLoop_acc_313_nl[7:0];
  assign nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3183:3176]));
  assign MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3191:3184]));
  assign MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_312_nl = (readslicef_15_8_7(MultLoop_398_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_399_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_312_nl = nl_MultLoop_acc_312_nl[7:0];
  assign nl_MultLoop_acc_366_nl = MultLoop_acc_315_nl + MultLoop_acc_314_nl + MultLoop_acc_313_nl
      + MultLoop_acc_312_nl;
  assign MultLoop_acc_366_nl = nl_MultLoop_acc_366_nl[7:0];
  assign nl_MultLoop_acc_375_nl = MultLoop_acc_367_nl + MultLoop_acc_366_nl;
  assign MultLoop_acc_375_nl = nl_MultLoop_acc_375_nl[7:0];
  assign nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3263:3256]));
  assign MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3271:3264]));
  assign MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_307_nl = (readslicef_15_8_7(MultLoop_408_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_409_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[7:0];
  assign nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3279:3272]));
  assign MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3287:3280]));
  assign MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_306_nl = (readslicef_15_8_7(MultLoop_410_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_411_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_306_nl = nl_MultLoop_acc_306_nl[7:0];
  assign nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3199:3192]));
  assign MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3207:3200]));
  assign MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_311_nl = (readslicef_15_8_7(MultLoop_400_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_401_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_311_nl = nl_MultLoop_acc_311_nl[7:0];
  assign nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3215:3208]));
  assign MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3223:3216]));
  assign MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_310_nl = (readslicef_15_8_7(MultLoop_402_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_403_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[7:0];
  assign nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3231:3224]));
  assign MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3239:3232]));
  assign MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_309_nl = (readslicef_15_8_7(MultLoop_404_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_405_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_309_nl = nl_MultLoop_acc_309_nl[7:0];
  assign nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3247:3240]));
  assign MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3255:3248]));
  assign MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_308_nl = (readslicef_15_8_7(MultLoop_406_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_407_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_308_nl = nl_MultLoop_acc_308_nl[7:0];
  assign nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3295:3288]));
  assign MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3303:3296]));
  assign MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_305_nl = (readslicef_15_8_7(MultLoop_412_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_413_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_305_nl = nl_MultLoop_acc_305_nl[7:0];
  assign nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3311:3304]));
  assign MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3319:3312]));
  assign MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_304_nl = (readslicef_15_8_7(MultLoop_414_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_415_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[7:0];
  assign nl_MultLoop_acc_374_nl = MultLoop_acc_307_nl + MultLoop_acc_306_nl + MultLoop_acc_311_nl
      + MultLoop_acc_310_nl + MultLoop_acc_309_nl + MultLoop_acc_308_nl + MultLoop_acc_305_nl
      + MultLoop_acc_304_nl;
  assign MultLoop_acc_374_nl = nl_MultLoop_acc_374_nl[7:0];
  assign nl_MultLoop_acc_379_nl = MultLoop_acc_375_nl + MultLoop_acc_374_nl;
  assign MultLoop_acc_379_nl = nl_MultLoop_acc_379_nl[7:0];
  assign nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3327:3320]));
  assign MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3335:3328]));
  assign MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_303_nl = (readslicef_15_8_7(MultLoop_416_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_417_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_303_nl = nl_MultLoop_acc_303_nl[7:0];
  assign nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3343:3336]));
  assign MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3351:3344]));
  assign MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_302_nl = (readslicef_15_8_7(MultLoop_418_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_419_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_302_nl = nl_MultLoop_acc_302_nl[7:0];
  assign nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3359:3352]));
  assign MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3367:3360]));
  assign MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_301_nl = (readslicef_15_8_7(MultLoop_420_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_421_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_301_nl = nl_MultLoop_acc_301_nl[7:0];
  assign nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3375:3368]));
  assign MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3383:3376]));
  assign MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_300_nl = (readslicef_15_8_7(MultLoop_422_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_423_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_300_nl = nl_MultLoop_acc_300_nl[7:0];
  assign nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3391:3384]));
  assign MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3399:3392]));
  assign MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_299_nl = (readslicef_15_8_7(MultLoop_424_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_425_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_299_nl = nl_MultLoop_acc_299_nl[7:0];
  assign nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3407:3400]));
  assign MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3415:3408]));
  assign MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_298_nl = (readslicef_15_8_7(MultLoop_426_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_427_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_298_nl = nl_MultLoop_acc_298_nl[7:0];
  assign nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3423:3416]));
  assign MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3431:3424]));
  assign MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_297_nl = (readslicef_15_8_7(MultLoop_428_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_429_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_297_nl = nl_MultLoop_acc_297_nl[7:0];
  assign nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3439:3432]));
  assign MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3447:3440]));
  assign MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_296_nl = (readslicef_15_8_7(MultLoop_430_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_431_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_296_nl = nl_MultLoop_acc_296_nl[7:0];
  assign nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3519:3512]));
  assign MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3527:3520]));
  assign MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_291_nl = (readslicef_15_8_7(MultLoop_440_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_441_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_291_nl = nl_MultLoop_acc_291_nl[7:0];
  assign nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3535:3528]));
  assign MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3543:3536]));
  assign MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_290_nl = (readslicef_15_8_7(MultLoop_442_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_443_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_290_nl = nl_MultLoop_acc_290_nl[7:0];
  assign nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3551:3544]));
  assign MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3559:3552]));
  assign MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_289_nl = (readslicef_15_8_7(MultLoop_444_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_445_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_289_nl = nl_MultLoop_acc_289_nl[7:0];
  assign nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3567:3560]));
  assign MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3575:3568]));
  assign MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_288_nl = (readslicef_15_8_7(MultLoop_446_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_447_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_288_nl = nl_MultLoop_acc_288_nl[7:0];
  assign nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3455:3448]));
  assign MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3463:3456]));
  assign MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_295_nl = (readslicef_15_8_7(MultLoop_432_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_433_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_295_nl = nl_MultLoop_acc_295_nl[7:0];
  assign nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3471:3464]));
  assign MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3479:3472]));
  assign MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_294_nl = (readslicef_15_8_7(MultLoop_434_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_435_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_294_nl = nl_MultLoop_acc_294_nl[7:0];
  assign nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3487:3480]));
  assign MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3495:3488]));
  assign MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_293_nl = (readslicef_15_8_7(MultLoop_436_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_437_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_293_nl = nl_MultLoop_acc_293_nl[7:0];
  assign nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3503:3496]));
  assign MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3511:3504]));
  assign MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_292_nl = (readslicef_15_8_7(MultLoop_438_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_439_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_292_nl = nl_MultLoop_acc_292_nl[7:0];
  assign nl_MultLoop_acc_378_nl = MultLoop_acc_303_nl + MultLoop_acc_302_nl + MultLoop_acc_301_nl
      + MultLoop_acc_300_nl + MultLoop_acc_299_nl + MultLoop_acc_298_nl + MultLoop_acc_297_nl
      + MultLoop_acc_296_nl + MultLoop_acc_291_nl + MultLoop_acc_290_nl + MultLoop_acc_289_nl
      + MultLoop_acc_288_nl + MultLoop_acc_295_nl + MultLoop_acc_294_nl + MultLoop_acc_293_nl
      + MultLoop_acc_292_nl;
  assign MultLoop_acc_378_nl = nl_MultLoop_acc_378_nl[7:0];
  assign nl_MultLoop_acc_381_nl = MultLoop_acc_379_nl + MultLoop_acc_378_nl;
  assign MultLoop_acc_381_nl = nl_MultLoop_acc_381_nl[7:0];
  assign nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3647:3640]));
  assign MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3655:3648]));
  assign MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_283_nl = (readslicef_15_8_7(MultLoop_456_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_457_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_283_nl = nl_MultLoop_acc_283_nl[7:0];
  assign nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3663:3656]));
  assign MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3671:3664]));
  assign MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_282_nl = (readslicef_15_8_7(MultLoop_458_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_459_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_282_nl = nl_MultLoop_acc_282_nl[7:0];
  assign nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3775:3768]));
  assign MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3783:3776]));
  assign MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_275_nl = (readslicef_15_8_7(MultLoop_472_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_473_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_275_nl = nl_MultLoop_acc_275_nl[7:0];
  assign nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3791:3784]));
  assign MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3799:3792]));
  assign MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_274_nl = (readslicef_15_8_7(MultLoop_474_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_475_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_274_nl = nl_MultLoop_acc_274_nl[7:0];
  assign nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3711:3704]));
  assign MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3719:3712]));
  assign MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_279_nl = (readslicef_15_8_7(MultLoop_464_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_465_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_279_nl = nl_MultLoop_acc_279_nl[7:0];
  assign nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3727:3720]));
  assign MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3735:3728]));
  assign MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_278_nl = (readslicef_15_8_7(MultLoop_466_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_467_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_278_nl = nl_MultLoop_acc_278_nl[7:0];
  assign nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4031:4024]));
  assign MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4039:4032]));
  assign MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_259_nl = (readslicef_15_8_7(MultLoop_504_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_505_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_259_nl = nl_MultLoop_acc_259_nl[7:0];
  assign nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4047:4040]));
  assign MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4055:4048]));
  assign MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_258_nl = (readslicef_15_8_7(MultLoop_506_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_258_nl = nl_MultLoop_acc_258_nl[7:0];
  assign nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3967:3960]));
  assign MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3975:3968]));
  assign MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_263_nl = (readslicef_15_8_7(MultLoop_496_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_497_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_263_nl = nl_MultLoop_acc_263_nl[7:0];
  assign nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3983:3976]));
  assign MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3991:3984]));
  assign MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_262_nl = (readslicef_15_8_7(MultLoop_498_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_499_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_262_nl = nl_MultLoop_acc_262_nl[7:0];
  assign nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3999:3992]));
  assign MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4007:4000]));
  assign MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_261_nl = (readslicef_15_8_7(MultLoop_500_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_501_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_261_nl = nl_MultLoop_acc_261_nl[7:0];
  assign nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4015:4008]));
  assign MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4023:4016]));
  assign MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_260_nl = (readslicef_15_8_7(MultLoop_502_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_503_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_260_nl = nl_MultLoop_acc_260_nl[7:0];
  assign nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3839:3832]));
  assign MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3847:3840]));
  assign MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_271_nl = (readslicef_15_8_7(MultLoop_480_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_481_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[7:0];
  assign nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3855:3848]));
  assign MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3863:3856]));
  assign MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_270_nl = (readslicef_15_8_7(MultLoop_482_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[7:0];
  assign nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3871:3864]));
  assign MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3879:3872]));
  assign MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_269_nl = (readslicef_15_8_7(MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_485_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_269_nl = nl_MultLoop_acc_269_nl[7:0];
  assign nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3887:3880]));
  assign MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3895:3888]));
  assign MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_268_nl = (readslicef_15_8_7(MultLoop_486_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_487_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_268_nl = nl_MultLoop_acc_268_nl[7:0];
  assign nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3903:3896]));
  assign MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3911:3904]));
  assign MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_267_nl = (readslicef_15_8_7(MultLoop_488_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_489_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_267_nl = nl_MultLoop_acc_267_nl[7:0];
  assign nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3919:3912]));
  assign MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3927:3920]));
  assign MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_266_nl = (readslicef_15_8_7(MultLoop_490_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_491_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_266_nl = nl_MultLoop_acc_266_nl[7:0];
  assign nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3935:3928]));
  assign MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3943:3936]));
  assign MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_265_nl = (readslicef_15_8_7(MultLoop_492_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_493_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_265_nl = nl_MultLoop_acc_265_nl[7:0];
  assign nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3951:3944]));
  assign MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3959:3952]));
  assign MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_264_nl = (readslicef_15_8_7(MultLoop_494_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_495_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_264_nl = nl_MultLoop_acc_264_nl[7:0];
  assign nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3583:3576]));
  assign MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3591:3584]));
  assign MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_287_nl = (readslicef_15_8_7(MultLoop_448_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_287_nl = nl_MultLoop_acc_287_nl[7:0];
  assign nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3599:3592]));
  assign MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3607:3600]));
  assign MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_286_nl = (readslicef_15_8_7(MultLoop_450_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_451_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_286_nl = nl_MultLoop_acc_286_nl[7:0];
  assign nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3615:3608]));
  assign MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3623:3616]));
  assign MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_285_nl = (readslicef_15_8_7(MultLoop_452_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_453_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_285_nl = nl_MultLoop_acc_285_nl[7:0];
  assign nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3631:3624]));
  assign MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3639:3632]));
  assign MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_284_nl = (readslicef_15_8_7(MultLoop_454_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_455_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_284_nl = nl_MultLoop_acc_284_nl[7:0];
  assign nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3679:3672]));
  assign MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3687:3680]));
  assign MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_281_nl = (readslicef_15_8_7(MultLoop_460_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_461_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_281_nl = nl_MultLoop_acc_281_nl[7:0];
  assign nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3695:3688]));
  assign MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3703:3696]));
  assign MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_280_nl = (readslicef_15_8_7(MultLoop_462_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_463_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_280_nl = nl_MultLoop_acc_280_nl[7:0];
  assign nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3743:3736]));
  assign MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3751:3744]));
  assign MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_277_nl = (readslicef_15_8_7(MultLoop_468_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_469_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_277_nl = nl_MultLoop_acc_277_nl[7:0];
  assign nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3759:3752]));
  assign MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3767:3760]));
  assign MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_276_nl = (readslicef_15_8_7(MultLoop_470_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_471_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_276_nl = nl_MultLoop_acc_276_nl[7:0];
  assign nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3807:3800]));
  assign MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3815:3808]));
  assign MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_273_nl = (readslicef_15_8_7(MultLoop_476_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_477_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_273_nl = nl_MultLoop_acc_273_nl[7:0];
  assign nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3823:3816]));
  assign MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[3831:3824]));
  assign MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_272_nl = (readslicef_15_8_7(MultLoop_478_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_479_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_272_nl = nl_MultLoop_acc_272_nl[7:0];
  assign nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4063:4056]));
  assign MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4071:4064]));
  assign MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_257_nl = (readslicef_15_8_7(MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_509_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_257_nl = nl_MultLoop_acc_257_nl[7:0];
  assign nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4079:4072]));
  assign MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4087:4080]));
  assign MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_256_nl = (readslicef_15_8_7(MultLoop_510_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_511_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_256_nl = nl_MultLoop_acc_256_nl[7:0];
  assign nl_MultLoop_acc_380_nl = MultLoop_acc_283_nl + MultLoop_acc_282_nl + MultLoop_acc_275_nl
      + MultLoop_acc_274_nl + MultLoop_acc_279_nl + MultLoop_acc_278_nl + MultLoop_acc_259_nl
      + MultLoop_acc_258_nl + MultLoop_acc_263_nl + MultLoop_acc_262_nl + MultLoop_acc_261_nl
      + MultLoop_acc_260_nl + MultLoop_acc_271_nl + MultLoop_acc_270_nl + MultLoop_acc_269_nl
      + MultLoop_acc_268_nl + MultLoop_acc_267_nl + MultLoop_acc_266_nl + MultLoop_acc_265_nl
      + MultLoop_acc_264_nl + MultLoop_acc_287_nl + MultLoop_acc_286_nl + MultLoop_acc_285_nl
      + MultLoop_acc_284_nl + MultLoop_acc_281_nl + MultLoop_acc_280_nl + MultLoop_acc_277_nl
      + MultLoop_acc_276_nl + MultLoop_acc_273_nl + MultLoop_acc_272_nl + MultLoop_acc_257_nl
      + MultLoop_acc_256_nl;
  assign MultLoop_acc_380_nl = nl_MultLoop_acc_380_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1 = MultLoop_acc_381_nl
      + MultLoop_acc_380_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1[7:0];
  assign nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7167:7160]));
  assign MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_636_nl = (readslicef_15_8_7(MultLoop_896_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[48:42]);
  assign MultLoop_acc_636_nl = nl_MultLoop_acc_636_nl[7:0];
  assign nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[6151:6144]));
  assign MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_700_nl = MultLoop_acc_636_nl + (readslicef_15_8_7(MultLoop_769_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_700_nl = nl_MultLoop_acc_700_nl[7:0];
  assign nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6159:6152]));
  assign MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6167:6160]));
  assign MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_699_nl = (readslicef_15_8_7(MultLoop_770_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_771_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_699_nl = nl_MultLoop_acc_699_nl[7:0];
  assign nl_MultLoop_acc_732_nl = MultLoop_acc_700_nl + MultLoop_acc_699_nl;
  assign MultLoop_acc_732_nl = nl_MultLoop_acc_732_nl[7:0];
  assign nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6175:6168]));
  assign MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6183:6176]));
  assign MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_698_nl = (readslicef_15_8_7(MultLoop_772_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_773_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_698_nl = nl_MultLoop_acc_698_nl[7:0];
  assign nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6191:6184]));
  assign MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6199:6192]));
  assign MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_697_nl = (readslicef_15_8_7(MultLoop_774_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_697_nl = nl_MultLoop_acc_697_nl[7:0];
  assign nl_MultLoop_acc_731_nl = MultLoop_acc_698_nl + MultLoop_acc_697_nl;
  assign MultLoop_acc_731_nl = nl_MultLoop_acc_731_nl[7:0];
  assign nl_MultLoop_acc_748_nl = MultLoop_acc_732_nl + MultLoop_acc_731_nl;
  assign MultLoop_acc_748_nl = nl_MultLoop_acc_748_nl[7:0];
  assign nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6207:6200]));
  assign MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6215:6208]));
  assign MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_696_nl = (readslicef_15_8_7(MultLoop_776_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_777_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_696_nl = nl_MultLoop_acc_696_nl[7:0];
  assign nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6223:6216]));
  assign MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6231:6224]));
  assign MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_695_nl = (readslicef_15_8_7(MultLoop_778_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_779_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_695_nl = nl_MultLoop_acc_695_nl[7:0];
  assign nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6239:6232]));
  assign MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6247:6240]));
  assign MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_694_nl = (readslicef_15_8_7(MultLoop_780_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_781_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_694_nl = nl_MultLoop_acc_694_nl[7:0];
  assign nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6255:6248]));
  assign MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6263:6256]));
  assign MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_693_nl = (readslicef_15_8_7(MultLoop_782_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_783_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_693_nl = nl_MultLoop_acc_693_nl[7:0];
  assign nl_MultLoop_acc_747_nl = MultLoop_acc_696_nl + MultLoop_acc_695_nl + MultLoop_acc_694_nl
      + MultLoop_acc_693_nl;
  assign MultLoop_acc_747_nl = nl_MultLoop_acc_747_nl[7:0];
  assign nl_MultLoop_acc_756_nl = MultLoop_acc_748_nl + MultLoop_acc_747_nl;
  assign MultLoop_acc_756_nl = nl_MultLoop_acc_756_nl[7:0];
  assign nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6335:6328]));
  assign MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6343:6336]));
  assign MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_688_nl = (readslicef_15_8_7(MultLoop_792_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_793_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_688_nl = nl_MultLoop_acc_688_nl[7:0];
  assign nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6351:6344]));
  assign MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6359:6352]));
  assign MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_687_nl = (readslicef_15_8_7(MultLoop_794_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_795_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_687_nl = nl_MultLoop_acc_687_nl[7:0];
  assign nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6271:6264]));
  assign MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6279:6272]));
  assign MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_692_nl = (readslicef_15_8_7(MultLoop_784_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_785_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_692_nl = nl_MultLoop_acc_692_nl[7:0];
  assign nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6287:6280]));
  assign MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6295:6288]));
  assign MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_691_nl = (readslicef_15_8_7(MultLoop_786_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_787_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_691_nl = nl_MultLoop_acc_691_nl[7:0];
  assign nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6303:6296]));
  assign MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6311:6304]));
  assign MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_690_nl = (readslicef_15_8_7(MultLoop_788_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_789_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_690_nl = nl_MultLoop_acc_690_nl[7:0];
  assign nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6319:6312]));
  assign MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6327:6320]));
  assign MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_689_nl = (readslicef_15_8_7(MultLoop_790_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_791_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_689_nl = nl_MultLoop_acc_689_nl[7:0];
  assign nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6367:6360]));
  assign MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6375:6368]));
  assign MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_686_nl = (readslicef_15_8_7(MultLoop_796_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_797_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_686_nl = nl_MultLoop_acc_686_nl[7:0];
  assign nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6383:6376]));
  assign MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6391:6384]));
  assign MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_685_nl = (readslicef_15_8_7(MultLoop_798_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_799_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_685_nl = nl_MultLoop_acc_685_nl[7:0];
  assign nl_MultLoop_acc_755_nl = MultLoop_acc_688_nl + MultLoop_acc_687_nl + MultLoop_acc_692_nl
      + MultLoop_acc_691_nl + MultLoop_acc_690_nl + MultLoop_acc_689_nl + MultLoop_acc_686_nl
      + MultLoop_acc_685_nl;
  assign MultLoop_acc_755_nl = nl_MultLoop_acc_755_nl[7:0];
  assign nl_MultLoop_acc_760_nl = MultLoop_acc_756_nl + MultLoop_acc_755_nl;
  assign MultLoop_acc_760_nl = nl_MultLoop_acc_760_nl[7:0];
  assign nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6399:6392]));
  assign MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6407:6400]));
  assign MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_684_nl = (readslicef_15_8_7(MultLoop_800_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_801_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_684_nl = nl_MultLoop_acc_684_nl[7:0];
  assign nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6415:6408]));
  assign MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6423:6416]));
  assign MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_683_nl = (readslicef_15_8_7(MultLoop_802_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_803_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_683_nl = nl_MultLoop_acc_683_nl[7:0];
  assign nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6431:6424]));
  assign MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6439:6432]));
  assign MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_682_nl = (readslicef_15_8_7(MultLoop_804_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_805_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_682_nl = nl_MultLoop_acc_682_nl[7:0];
  assign nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6447:6440]));
  assign MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6455:6448]));
  assign MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_681_nl = (readslicef_15_8_7(MultLoop_806_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_807_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_681_nl = nl_MultLoop_acc_681_nl[7:0];
  assign nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6463:6456]));
  assign MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6471:6464]));
  assign MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_680_nl = (readslicef_15_8_7(MultLoop_808_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_809_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_680_nl = nl_MultLoop_acc_680_nl[7:0];
  assign nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6479:6472]));
  assign MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6487:6480]));
  assign MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_679_nl = (readslicef_15_8_7(MultLoop_810_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_811_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_679_nl = nl_MultLoop_acc_679_nl[7:0];
  assign nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6495:6488]));
  assign MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6503:6496]));
  assign MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_678_nl = (readslicef_15_8_7(MultLoop_812_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_813_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_678_nl = nl_MultLoop_acc_678_nl[7:0];
  assign nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6511:6504]));
  assign MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6519:6512]));
  assign MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_677_nl = (readslicef_15_8_7(MultLoop_814_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_815_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_677_nl = nl_MultLoop_acc_677_nl[7:0];
  assign nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6591:6584]));
  assign MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6599:6592]));
  assign MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_672_nl = (readslicef_15_8_7(MultLoop_824_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_825_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_672_nl = nl_MultLoop_acc_672_nl[7:0];
  assign nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6607:6600]));
  assign MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6615:6608]));
  assign MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_671_nl = (readslicef_15_8_7(MultLoop_826_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_827_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_671_nl = nl_MultLoop_acc_671_nl[7:0];
  assign nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6623:6616]));
  assign MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6631:6624]));
  assign MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_670_nl = (readslicef_15_8_7(MultLoop_828_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_829_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_670_nl = nl_MultLoop_acc_670_nl[7:0];
  assign nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6639:6632]));
  assign MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6647:6640]));
  assign MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_669_nl = (readslicef_15_8_7(MultLoop_830_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_831_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_669_nl = nl_MultLoop_acc_669_nl[7:0];
  assign nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6527:6520]));
  assign MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6535:6528]));
  assign MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_676_nl = (readslicef_15_8_7(MultLoop_816_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_817_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_676_nl = nl_MultLoop_acc_676_nl[7:0];
  assign nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6543:6536]));
  assign MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6551:6544]));
  assign MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_675_nl = (readslicef_15_8_7(MultLoop_818_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_819_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_675_nl = nl_MultLoop_acc_675_nl[7:0];
  assign nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6559:6552]));
  assign MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6567:6560]));
  assign MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_674_nl = (readslicef_15_8_7(MultLoop_820_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_821_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_674_nl = nl_MultLoop_acc_674_nl[7:0];
  assign nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6575:6568]));
  assign MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6583:6576]));
  assign MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_673_nl = (readslicef_15_8_7(MultLoop_822_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_823_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_673_nl = nl_MultLoop_acc_673_nl[7:0];
  assign nl_MultLoop_acc_759_nl = MultLoop_acc_684_nl + MultLoop_acc_683_nl + MultLoop_acc_682_nl
      + MultLoop_acc_681_nl + MultLoop_acc_680_nl + MultLoop_acc_679_nl + MultLoop_acc_678_nl
      + MultLoop_acc_677_nl + MultLoop_acc_672_nl + MultLoop_acc_671_nl + MultLoop_acc_670_nl
      + MultLoop_acc_669_nl + MultLoop_acc_676_nl + MultLoop_acc_675_nl + MultLoop_acc_674_nl
      + MultLoop_acc_673_nl;
  assign MultLoop_acc_759_nl = nl_MultLoop_acc_759_nl[7:0];
  assign nl_MultLoop_acc_762_nl = MultLoop_acc_760_nl + MultLoop_acc_759_nl;
  assign MultLoop_acc_762_nl = nl_MultLoop_acc_762_nl[7:0];
  assign nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6719:6712]));
  assign MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6727:6720]));
  assign MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_664_nl = (readslicef_15_8_7(MultLoop_840_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_841_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_664_nl = nl_MultLoop_acc_664_nl[7:0];
  assign nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6735:6728]));
  assign MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6743:6736]));
  assign MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_663_nl = (readslicef_15_8_7(MultLoop_842_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_843_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_663_nl = nl_MultLoop_acc_663_nl[7:0];
  assign nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6847:6840]));
  assign MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6855:6848]));
  assign MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_656_nl = (readslicef_15_8_7(MultLoop_856_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_857_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_656_nl = nl_MultLoop_acc_656_nl[7:0];
  assign nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6863:6856]));
  assign MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6871:6864]));
  assign MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_655_nl = (readslicef_15_8_7(MultLoop_858_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_859_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_655_nl = nl_MultLoop_acc_655_nl[7:0];
  assign nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6783:6776]));
  assign MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6791:6784]));
  assign MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_660_nl = (readslicef_15_8_7(MultLoop_848_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_849_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_660_nl = nl_MultLoop_acc_660_nl[7:0];
  assign nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6799:6792]));
  assign MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6807:6800]));
  assign MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_659_nl = (readslicef_15_8_7(MultLoop_850_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_851_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_659_nl = nl_MultLoop_acc_659_nl[7:0];
  assign nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7103:7096]));
  assign MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7111:7104]));
  assign MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_640_nl = (readslicef_15_8_7(MultLoop_888_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_889_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_640_nl = nl_MultLoop_acc_640_nl[7:0];
  assign nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7119:7112]));
  assign MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7127:7120]));
  assign MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_639_nl = (readslicef_15_8_7(MultLoop_890_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_891_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_639_nl = nl_MultLoop_acc_639_nl[7:0];
  assign nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7039:7032]));
  assign MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7047:7040]));
  assign MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_644_nl = (readslicef_15_8_7(MultLoop_880_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_881_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_644_nl = nl_MultLoop_acc_644_nl[7:0];
  assign nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7055:7048]));
  assign MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7063:7056]));
  assign MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_643_nl = (readslicef_15_8_7(MultLoop_882_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_883_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_643_nl = nl_MultLoop_acc_643_nl[7:0];
  assign nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7071:7064]));
  assign MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7079:7072]));
  assign MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_642_nl = (readslicef_15_8_7(MultLoop_884_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_885_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_642_nl = nl_MultLoop_acc_642_nl[7:0];
  assign nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7087:7080]));
  assign MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7095:7088]));
  assign MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_641_nl = (readslicef_15_8_7(MultLoop_886_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_887_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_641_nl = nl_MultLoop_acc_641_nl[7:0];
  assign nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6911:6904]));
  assign MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6919:6912]));
  assign MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_652_nl = (readslicef_15_8_7(MultLoop_864_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_865_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_652_nl = nl_MultLoop_acc_652_nl[7:0];
  assign nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6927:6920]));
  assign MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6935:6928]));
  assign MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_651_nl = (readslicef_15_8_7(MultLoop_866_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_651_nl = nl_MultLoop_acc_651_nl[7:0];
  assign nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6943:6936]));
  assign MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6951:6944]));
  assign MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_650_nl = (readslicef_15_8_7(MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_869_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_650_nl = nl_MultLoop_acc_650_nl[7:0];
  assign nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6959:6952]));
  assign MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6967:6960]));
  assign MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_649_nl = (readslicef_15_8_7(MultLoop_870_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_871_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_649_nl = nl_MultLoop_acc_649_nl[7:0];
  assign nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6975:6968]));
  assign MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6983:6976]));
  assign MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_648_nl = (readslicef_15_8_7(MultLoop_872_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_873_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_648_nl = nl_MultLoop_acc_648_nl[7:0];
  assign nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6991:6984]));
  assign MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6999:6992]));
  assign MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_647_nl = (readslicef_15_8_7(MultLoop_874_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_875_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_647_nl = nl_MultLoop_acc_647_nl[7:0];
  assign nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7007:7000]));
  assign MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7015:7008]));
  assign MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_646_nl = (readslicef_15_8_7(MultLoop_876_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_877_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_646_nl = nl_MultLoop_acc_646_nl[7:0];
  assign nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7023:7016]));
  assign MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7031:7024]));
  assign MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_645_nl = (readslicef_15_8_7(MultLoop_878_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_879_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_645_nl = nl_MultLoop_acc_645_nl[7:0];
  assign nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6655:6648]));
  assign MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6663:6656]));
  assign MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_668_nl = (readslicef_15_8_7(MultLoop_832_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_668_nl = nl_MultLoop_acc_668_nl[7:0];
  assign nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6671:6664]));
  assign MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6679:6672]));
  assign MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_667_nl = (readslicef_15_8_7(MultLoop_834_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_835_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_667_nl = nl_MultLoop_acc_667_nl[7:0];
  assign nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6687:6680]));
  assign MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6695:6688]));
  assign MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_666_nl = (readslicef_15_8_7(MultLoop_836_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_837_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_666_nl = nl_MultLoop_acc_666_nl[7:0];
  assign nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6703:6696]));
  assign MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6711:6704]));
  assign MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_665_nl = (readslicef_15_8_7(MultLoop_838_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_839_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_665_nl = nl_MultLoop_acc_665_nl[7:0];
  assign nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6751:6744]));
  assign MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6759:6752]));
  assign MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_662_nl = (readslicef_15_8_7(MultLoop_844_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_845_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_662_nl = nl_MultLoop_acc_662_nl[7:0];
  assign nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6767:6760]));
  assign MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6775:6768]));
  assign MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_661_nl = (readslicef_15_8_7(MultLoop_846_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_847_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_661_nl = nl_MultLoop_acc_661_nl[7:0];
  assign nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6815:6808]));
  assign MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6823:6816]));
  assign MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_658_nl = (readslicef_15_8_7(MultLoop_852_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_853_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_658_nl = nl_MultLoop_acc_658_nl[7:0];
  assign nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6831:6824]));
  assign MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6839:6832]));
  assign MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_657_nl = (readslicef_15_8_7(MultLoop_854_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_855_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_657_nl = nl_MultLoop_acc_657_nl[7:0];
  assign nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6879:6872]));
  assign MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6887:6880]));
  assign MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_654_nl = (readslicef_15_8_7(MultLoop_860_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_861_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_654_nl = nl_MultLoop_acc_654_nl[7:0];
  assign nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6895:6888]));
  assign MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6903:6896]));
  assign MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_653_nl = (readslicef_15_8_7(MultLoop_862_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_863_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_653_nl = nl_MultLoop_acc_653_nl[7:0];
  assign nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7135:7128]));
  assign MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7143:7136]));
  assign MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_638_nl = (readslicef_15_8_7(MultLoop_892_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_893_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_638_nl = nl_MultLoop_acc_638_nl[7:0];
  assign nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7151:7144]));
  assign MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[7159:7152]));
  assign MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_637_nl = (readslicef_15_8_7(MultLoop_894_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_895_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_637_nl = nl_MultLoop_acc_637_nl[7:0];
  assign nl_MultLoop_acc_761_nl = MultLoop_acc_664_nl + MultLoop_acc_663_nl + MultLoop_acc_656_nl
      + MultLoop_acc_655_nl + MultLoop_acc_660_nl + MultLoop_acc_659_nl + MultLoop_acc_640_nl
      + MultLoop_acc_639_nl + MultLoop_acc_644_nl + MultLoop_acc_643_nl + MultLoop_acc_642_nl
      + MultLoop_acc_641_nl + MultLoop_acc_652_nl + MultLoop_acc_651_nl + MultLoop_acc_650_nl
      + MultLoop_acc_649_nl + MultLoop_acc_648_nl + MultLoop_acc_647_nl + MultLoop_acc_646_nl
      + MultLoop_acc_645_nl + MultLoop_acc_668_nl + MultLoop_acc_667_nl + MultLoop_acc_666_nl
      + MultLoop_acc_665_nl + MultLoop_acc_662_nl + MultLoop_acc_661_nl + MultLoop_acc_658_nl
      + MultLoop_acc_657_nl + MultLoop_acc_654_nl + MultLoop_acc_653_nl + MultLoop_acc_638_nl
      + MultLoop_acc_637_nl;
  assign MultLoop_acc_761_nl = nl_MultLoop_acc_761_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1 = MultLoop_acc_762_nl
      + MultLoop_acc_761_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1[7:0];
  assign nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5119:5112]));
  assign MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_382_nl = (readslicef_15_8_7(MultLoop_640_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[34:28]);
  assign MultLoop_acc_382_nl = nl_MultLoop_acc_382_nl[7:0];
  assign nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[4103:4096]));
  assign MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_446_nl = MultLoop_acc_382_nl + (readslicef_15_8_7(MultLoop_513_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_446_nl = nl_MultLoop_acc_446_nl[7:0];
  assign nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4111:4104]));
  assign MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4119:4112]));
  assign MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_445_nl = (readslicef_15_8_7(MultLoop_514_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_515_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_445_nl = nl_MultLoop_acc_445_nl[7:0];
  assign nl_MultLoop_acc_478_nl = MultLoop_acc_446_nl + MultLoop_acc_445_nl;
  assign MultLoop_acc_478_nl = nl_MultLoop_acc_478_nl[7:0];
  assign nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4127:4120]));
  assign MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4135:4128]));
  assign MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_444_nl = (readslicef_15_8_7(MultLoop_516_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_517_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_444_nl = nl_MultLoop_acc_444_nl[7:0];
  assign nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4143:4136]));
  assign MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4151:4144]));
  assign MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_443_nl = (readslicef_15_8_7(MultLoop_518_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_443_nl = nl_MultLoop_acc_443_nl[7:0];
  assign nl_MultLoop_acc_477_nl = MultLoop_acc_444_nl + MultLoop_acc_443_nl;
  assign MultLoop_acc_477_nl = nl_MultLoop_acc_477_nl[7:0];
  assign nl_MultLoop_acc_494_nl = MultLoop_acc_478_nl + MultLoop_acc_477_nl;
  assign MultLoop_acc_494_nl = nl_MultLoop_acc_494_nl[7:0];
  assign nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4159:4152]));
  assign MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4167:4160]));
  assign MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_442_nl = (readslicef_15_8_7(MultLoop_520_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_521_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_442_nl = nl_MultLoop_acc_442_nl[7:0];
  assign nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4175:4168]));
  assign MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4183:4176]));
  assign MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_441_nl = (readslicef_15_8_7(MultLoop_522_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_523_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_441_nl = nl_MultLoop_acc_441_nl[7:0];
  assign nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4191:4184]));
  assign MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4199:4192]));
  assign MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_440_nl = (readslicef_15_8_7(MultLoop_524_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_525_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_440_nl = nl_MultLoop_acc_440_nl[7:0];
  assign nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4207:4200]));
  assign MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4215:4208]));
  assign MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_439_nl = (readslicef_15_8_7(MultLoop_526_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_527_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_439_nl = nl_MultLoop_acc_439_nl[7:0];
  assign nl_MultLoop_acc_493_nl = MultLoop_acc_442_nl + MultLoop_acc_441_nl + MultLoop_acc_440_nl
      + MultLoop_acc_439_nl;
  assign MultLoop_acc_493_nl = nl_MultLoop_acc_493_nl[7:0];
  assign nl_MultLoop_acc_502_nl = MultLoop_acc_494_nl + MultLoop_acc_493_nl;
  assign MultLoop_acc_502_nl = nl_MultLoop_acc_502_nl[7:0];
  assign nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4287:4280]));
  assign MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4295:4288]));
  assign MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_434_nl = (readslicef_15_8_7(MultLoop_536_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_537_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_434_nl = nl_MultLoop_acc_434_nl[7:0];
  assign nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4303:4296]));
  assign MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4311:4304]));
  assign MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_433_nl = (readslicef_15_8_7(MultLoop_538_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_539_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_433_nl = nl_MultLoop_acc_433_nl[7:0];
  assign nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4223:4216]));
  assign MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4231:4224]));
  assign MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_438_nl = (readslicef_15_8_7(MultLoop_528_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_529_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_438_nl = nl_MultLoop_acc_438_nl[7:0];
  assign nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4239:4232]));
  assign MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4247:4240]));
  assign MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_437_nl = (readslicef_15_8_7(MultLoop_530_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_531_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_437_nl = nl_MultLoop_acc_437_nl[7:0];
  assign nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4255:4248]));
  assign MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4263:4256]));
  assign MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_436_nl = (readslicef_15_8_7(MultLoop_532_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_533_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_436_nl = nl_MultLoop_acc_436_nl[7:0];
  assign nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4271:4264]));
  assign MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4279:4272]));
  assign MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_435_nl = (readslicef_15_8_7(MultLoop_534_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_535_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_435_nl = nl_MultLoop_acc_435_nl[7:0];
  assign nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4319:4312]));
  assign MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4327:4320]));
  assign MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_432_nl = (readslicef_15_8_7(MultLoop_540_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_541_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_432_nl = nl_MultLoop_acc_432_nl[7:0];
  assign nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4335:4328]));
  assign MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4343:4336]));
  assign MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_431_nl = (readslicef_15_8_7(MultLoop_542_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_543_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_431_nl = nl_MultLoop_acc_431_nl[7:0];
  assign nl_MultLoop_acc_501_nl = MultLoop_acc_434_nl + MultLoop_acc_433_nl + MultLoop_acc_438_nl
      + MultLoop_acc_437_nl + MultLoop_acc_436_nl + MultLoop_acc_435_nl + MultLoop_acc_432_nl
      + MultLoop_acc_431_nl;
  assign MultLoop_acc_501_nl = nl_MultLoop_acc_501_nl[7:0];
  assign nl_MultLoop_acc_506_nl = MultLoop_acc_502_nl + MultLoop_acc_501_nl;
  assign MultLoop_acc_506_nl = nl_MultLoop_acc_506_nl[7:0];
  assign nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4351:4344]));
  assign MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4359:4352]));
  assign MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_430_nl = (readslicef_15_8_7(MultLoop_544_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_545_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_430_nl = nl_MultLoop_acc_430_nl[7:0];
  assign nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4367:4360]));
  assign MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4375:4368]));
  assign MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_429_nl = (readslicef_15_8_7(MultLoop_546_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_547_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_429_nl = nl_MultLoop_acc_429_nl[7:0];
  assign nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4383:4376]));
  assign MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4391:4384]));
  assign MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_428_nl = (readslicef_15_8_7(MultLoop_548_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_549_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_428_nl = nl_MultLoop_acc_428_nl[7:0];
  assign nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4399:4392]));
  assign MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4407:4400]));
  assign MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_427_nl = (readslicef_15_8_7(MultLoop_550_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_551_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_427_nl = nl_MultLoop_acc_427_nl[7:0];
  assign nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4415:4408]));
  assign MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4423:4416]));
  assign MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_426_nl = (readslicef_15_8_7(MultLoop_552_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_553_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_426_nl = nl_MultLoop_acc_426_nl[7:0];
  assign nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4431:4424]));
  assign MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4439:4432]));
  assign MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_425_nl = (readslicef_15_8_7(MultLoop_554_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_555_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_425_nl = nl_MultLoop_acc_425_nl[7:0];
  assign nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4447:4440]));
  assign MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4455:4448]));
  assign MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_424_nl = (readslicef_15_8_7(MultLoop_556_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_557_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_424_nl = nl_MultLoop_acc_424_nl[7:0];
  assign nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4463:4456]));
  assign MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4471:4464]));
  assign MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_423_nl = (readslicef_15_8_7(MultLoop_558_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_559_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_423_nl = nl_MultLoop_acc_423_nl[7:0];
  assign nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4543:4536]));
  assign MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4551:4544]));
  assign MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_418_nl = (readslicef_15_8_7(MultLoop_568_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_569_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_418_nl = nl_MultLoop_acc_418_nl[7:0];
  assign nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4559:4552]));
  assign MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4567:4560]));
  assign MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_417_nl = (readslicef_15_8_7(MultLoop_570_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_571_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_417_nl = nl_MultLoop_acc_417_nl[7:0];
  assign nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4575:4568]));
  assign MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4583:4576]));
  assign MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_416_nl = (readslicef_15_8_7(MultLoop_572_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_573_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_416_nl = nl_MultLoop_acc_416_nl[7:0];
  assign nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4591:4584]));
  assign MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4599:4592]));
  assign MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_415_nl = (readslicef_15_8_7(MultLoop_574_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_575_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_415_nl = nl_MultLoop_acc_415_nl[7:0];
  assign nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4479:4472]));
  assign MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4487:4480]));
  assign MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_422_nl = (readslicef_15_8_7(MultLoop_560_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_561_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_422_nl = nl_MultLoop_acc_422_nl[7:0];
  assign nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4495:4488]));
  assign MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4503:4496]));
  assign MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_421_nl = (readslicef_15_8_7(MultLoop_562_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_563_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_421_nl = nl_MultLoop_acc_421_nl[7:0];
  assign nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4511:4504]));
  assign MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4519:4512]));
  assign MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_420_nl = (readslicef_15_8_7(MultLoop_564_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_565_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_420_nl = nl_MultLoop_acc_420_nl[7:0];
  assign nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4527:4520]));
  assign MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4535:4528]));
  assign MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_419_nl = (readslicef_15_8_7(MultLoop_566_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_567_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_419_nl = nl_MultLoop_acc_419_nl[7:0];
  assign nl_MultLoop_acc_505_nl = MultLoop_acc_430_nl + MultLoop_acc_429_nl + MultLoop_acc_428_nl
      + MultLoop_acc_427_nl + MultLoop_acc_426_nl + MultLoop_acc_425_nl + MultLoop_acc_424_nl
      + MultLoop_acc_423_nl + MultLoop_acc_418_nl + MultLoop_acc_417_nl + MultLoop_acc_416_nl
      + MultLoop_acc_415_nl + MultLoop_acc_422_nl + MultLoop_acc_421_nl + MultLoop_acc_420_nl
      + MultLoop_acc_419_nl;
  assign MultLoop_acc_505_nl = nl_MultLoop_acc_505_nl[7:0];
  assign nl_MultLoop_acc_508_nl = MultLoop_acc_506_nl + MultLoop_acc_505_nl;
  assign MultLoop_acc_508_nl = nl_MultLoop_acc_508_nl[7:0];
  assign nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4671:4664]));
  assign MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4679:4672]));
  assign MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_410_nl = (readslicef_15_8_7(MultLoop_584_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_585_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_410_nl = nl_MultLoop_acc_410_nl[7:0];
  assign nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4687:4680]));
  assign MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4695:4688]));
  assign MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_409_nl = (readslicef_15_8_7(MultLoop_586_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_587_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_409_nl = nl_MultLoop_acc_409_nl[7:0];
  assign nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4799:4792]));
  assign MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4807:4800]));
  assign MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_402_nl = (readslicef_15_8_7(MultLoop_600_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_601_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_402_nl = nl_MultLoop_acc_402_nl[7:0];
  assign nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4815:4808]));
  assign MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4823:4816]));
  assign MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_401_nl = (readslicef_15_8_7(MultLoop_602_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_603_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_401_nl = nl_MultLoop_acc_401_nl[7:0];
  assign nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4735:4728]));
  assign MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4743:4736]));
  assign MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_406_nl = (readslicef_15_8_7(MultLoop_592_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_593_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_406_nl = nl_MultLoop_acc_406_nl[7:0];
  assign nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4751:4744]));
  assign MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4759:4752]));
  assign MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_405_nl = (readslicef_15_8_7(MultLoop_594_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_595_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_405_nl = nl_MultLoop_acc_405_nl[7:0];
  assign nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5055:5048]));
  assign MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5063:5056]));
  assign MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_386_nl = (readslicef_15_8_7(MultLoop_632_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_633_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_386_nl = nl_MultLoop_acc_386_nl[7:0];
  assign nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5071:5064]));
  assign MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5079:5072]));
  assign MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_385_nl = (readslicef_15_8_7(MultLoop_634_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_635_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_385_nl = nl_MultLoop_acc_385_nl[7:0];
  assign nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4991:4984]));
  assign MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4999:4992]));
  assign MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_390_nl = (readslicef_15_8_7(MultLoop_624_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_625_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_390_nl = nl_MultLoop_acc_390_nl[7:0];
  assign nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5007:5000]));
  assign MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5015:5008]));
  assign MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_389_nl = (readslicef_15_8_7(MultLoop_626_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_627_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_389_nl = nl_MultLoop_acc_389_nl[7:0];
  assign nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5023:5016]));
  assign MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5031:5024]));
  assign MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_388_nl = (readslicef_15_8_7(MultLoop_628_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_629_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_388_nl = nl_MultLoop_acc_388_nl[7:0];
  assign nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5039:5032]));
  assign MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5047:5040]));
  assign MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_387_nl = (readslicef_15_8_7(MultLoop_630_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_631_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_387_nl = nl_MultLoop_acc_387_nl[7:0];
  assign nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4863:4856]));
  assign MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4871:4864]));
  assign MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_398_nl = (readslicef_15_8_7(MultLoop_608_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_609_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_398_nl = nl_MultLoop_acc_398_nl[7:0];
  assign nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4879:4872]));
  assign MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4887:4880]));
  assign MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_397_nl = (readslicef_15_8_7(MultLoop_610_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_397_nl = nl_MultLoop_acc_397_nl[7:0];
  assign nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4895:4888]));
  assign MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4903:4896]));
  assign MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_396_nl = (readslicef_15_8_7(MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_613_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_396_nl = nl_MultLoop_acc_396_nl[7:0];
  assign nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4911:4904]));
  assign MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4919:4912]));
  assign MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_395_nl = (readslicef_15_8_7(MultLoop_614_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_615_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_395_nl = nl_MultLoop_acc_395_nl[7:0];
  assign nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4927:4920]));
  assign MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4935:4928]));
  assign MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_394_nl = (readslicef_15_8_7(MultLoop_616_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_617_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_394_nl = nl_MultLoop_acc_394_nl[7:0];
  assign nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4943:4936]));
  assign MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4951:4944]));
  assign MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_393_nl = (readslicef_15_8_7(MultLoop_618_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_619_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_393_nl = nl_MultLoop_acc_393_nl[7:0];
  assign nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4959:4952]));
  assign MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4967:4960]));
  assign MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_392_nl = (readslicef_15_8_7(MultLoop_620_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_621_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_392_nl = nl_MultLoop_acc_392_nl[7:0];
  assign nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4975:4968]));
  assign MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4983:4976]));
  assign MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_391_nl = (readslicef_15_8_7(MultLoop_622_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_623_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_391_nl = nl_MultLoop_acc_391_nl[7:0];
  assign nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4607:4600]));
  assign MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4615:4608]));
  assign MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_414_nl = (readslicef_15_8_7(MultLoop_576_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_414_nl = nl_MultLoop_acc_414_nl[7:0];
  assign nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4623:4616]));
  assign MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4631:4624]));
  assign MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_413_nl = (readslicef_15_8_7(MultLoop_578_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_579_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_413_nl = nl_MultLoop_acc_413_nl[7:0];
  assign nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4639:4632]));
  assign MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4647:4640]));
  assign MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_412_nl = (readslicef_15_8_7(MultLoop_580_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_581_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_412_nl = nl_MultLoop_acc_412_nl[7:0];
  assign nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4655:4648]));
  assign MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4663:4656]));
  assign MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_411_nl = (readslicef_15_8_7(MultLoop_582_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_583_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_411_nl = nl_MultLoop_acc_411_nl[7:0];
  assign nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4703:4696]));
  assign MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4711:4704]));
  assign MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_408_nl = (readslicef_15_8_7(MultLoop_588_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_589_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_408_nl = nl_MultLoop_acc_408_nl[7:0];
  assign nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4719:4712]));
  assign MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4727:4720]));
  assign MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_407_nl = (readslicef_15_8_7(MultLoop_590_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_591_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_407_nl = nl_MultLoop_acc_407_nl[7:0];
  assign nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4767:4760]));
  assign MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4775:4768]));
  assign MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_404_nl = (readslicef_15_8_7(MultLoop_596_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_597_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_404_nl = nl_MultLoop_acc_404_nl[7:0];
  assign nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4783:4776]));
  assign MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4791:4784]));
  assign MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_403_nl = (readslicef_15_8_7(MultLoop_598_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_599_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_403_nl = nl_MultLoop_acc_403_nl[7:0];
  assign nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4831:4824]));
  assign MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4839:4832]));
  assign MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_400_nl = (readslicef_15_8_7(MultLoop_604_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_605_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_400_nl = nl_MultLoop_acc_400_nl[7:0];
  assign nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4847:4840]));
  assign MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[4855:4848]));
  assign MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_399_nl = (readslicef_15_8_7(MultLoop_606_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_607_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_399_nl = nl_MultLoop_acc_399_nl[7:0];
  assign nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5087:5080]));
  assign MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5095:5088]));
  assign MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_384_nl = (readslicef_15_8_7(MultLoop_636_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_637_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_384_nl = nl_MultLoop_acc_384_nl[7:0];
  assign nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5103:5096]));
  assign MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5111:5104]));
  assign MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_383_nl = (readslicef_15_8_7(MultLoop_638_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_639_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_383_nl = nl_MultLoop_acc_383_nl[7:0];
  assign nl_MultLoop_acc_507_nl = MultLoop_acc_410_nl + MultLoop_acc_409_nl + MultLoop_acc_402_nl
      + MultLoop_acc_401_nl + MultLoop_acc_406_nl + MultLoop_acc_405_nl + MultLoop_acc_386_nl
      + MultLoop_acc_385_nl + MultLoop_acc_390_nl + MultLoop_acc_389_nl + MultLoop_acc_388_nl
      + MultLoop_acc_387_nl + MultLoop_acc_398_nl + MultLoop_acc_397_nl + MultLoop_acc_396_nl
      + MultLoop_acc_395_nl + MultLoop_acc_394_nl + MultLoop_acc_393_nl + MultLoop_acc_392_nl
      + MultLoop_acc_391_nl + MultLoop_acc_414_nl + MultLoop_acc_413_nl + MultLoop_acc_412_nl
      + MultLoop_acc_411_nl + MultLoop_acc_408_nl + MultLoop_acc_407_nl + MultLoop_acc_404_nl
      + MultLoop_acc_403_nl + MultLoop_acc_400_nl + MultLoop_acc_399_nl + MultLoop_acc_384_nl
      + MultLoop_acc_383_nl;
  assign MultLoop_acc_507_nl = nl_MultLoop_acc_507_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1 = MultLoop_acc_508_nl
      + MultLoop_acc_507_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1[7:0];
  assign nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6143:6136]));
  assign MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_509_nl = (readslicef_15_8_7(MultLoop_768_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + conv_s2s_7_8(b4_rsci_idat_mxwt[41:35]);
  assign MultLoop_acc_509_nl = nl_MultLoop_acc_509_nl[7:0];
  assign nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289))
      * $signed((w4_rsci_idat_mxwt[5127:5120]));
  assign MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_573_nl = MultLoop_acc_509_nl + (readslicef_15_8_7(MultLoop_641_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_573_nl = nl_MultLoop_acc_573_nl[7:0];
  assign nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5135:5128]));
  assign MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5143:5136]));
  assign MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_572_nl = (readslicef_15_8_7(MultLoop_642_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_643_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_572_nl = nl_MultLoop_acc_572_nl[7:0];
  assign nl_MultLoop_acc_605_nl = MultLoop_acc_573_nl + MultLoop_acc_572_nl;
  assign MultLoop_acc_605_nl = nl_MultLoop_acc_605_nl[7:0];
  assign nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5151:5144]));
  assign MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5159:5152]));
  assign MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_571_nl = (readslicef_15_8_7(MultLoop_644_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_645_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_571_nl = nl_MultLoop_acc_571_nl[7:0];
  assign nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5167:5160]));
  assign MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5175:5168]));
  assign MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_570_nl = (readslicef_15_8_7(MultLoop_646_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_570_nl = nl_MultLoop_acc_570_nl[7:0];
  assign nl_MultLoop_acc_604_nl = MultLoop_acc_571_nl + MultLoop_acc_570_nl;
  assign MultLoop_acc_604_nl = nl_MultLoop_acc_604_nl[7:0];
  assign nl_MultLoop_acc_621_nl = MultLoop_acc_605_nl + MultLoop_acc_604_nl;
  assign MultLoop_acc_621_nl = nl_MultLoop_acc_621_nl[7:0];
  assign nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5183:5176]));
  assign MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5191:5184]));
  assign MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_569_nl = (readslicef_15_8_7(MultLoop_648_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_649_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_569_nl = nl_MultLoop_acc_569_nl[7:0];
  assign nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5199:5192]));
  assign MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5207:5200]));
  assign MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_568_nl = (readslicef_15_8_7(MultLoop_650_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_651_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_568_nl = nl_MultLoop_acc_568_nl[7:0];
  assign nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5215:5208]));
  assign MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5223:5216]));
  assign MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_567_nl = (readslicef_15_8_7(MultLoop_652_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_653_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_567_nl = nl_MultLoop_acc_567_nl[7:0];
  assign nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5231:5224]));
  assign MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5239:5232]));
  assign MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_566_nl = (readslicef_15_8_7(MultLoop_654_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_655_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_566_nl = nl_MultLoop_acc_566_nl[7:0];
  assign nl_MultLoop_acc_620_nl = MultLoop_acc_569_nl + MultLoop_acc_568_nl + MultLoop_acc_567_nl
      + MultLoop_acc_566_nl;
  assign MultLoop_acc_620_nl = nl_MultLoop_acc_620_nl[7:0];
  assign nl_MultLoop_acc_629_nl = MultLoop_acc_621_nl + MultLoop_acc_620_nl;
  assign MultLoop_acc_629_nl = nl_MultLoop_acc_629_nl[7:0];
  assign nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5311:5304]));
  assign MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5319:5312]));
  assign MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_561_nl = (readslicef_15_8_7(MultLoop_664_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_665_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_561_nl = nl_MultLoop_acc_561_nl[7:0];
  assign nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5327:5320]));
  assign MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5335:5328]));
  assign MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_560_nl = (readslicef_15_8_7(MultLoop_666_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_667_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_560_nl = nl_MultLoop_acc_560_nl[7:0];
  assign nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5247:5240]));
  assign MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5255:5248]));
  assign MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_565_nl = (readslicef_15_8_7(MultLoop_656_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_657_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_565_nl = nl_MultLoop_acc_565_nl[7:0];
  assign nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5263:5256]));
  assign MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5271:5264]));
  assign MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_564_nl = (readslicef_15_8_7(MultLoop_658_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_659_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_564_nl = nl_MultLoop_acc_564_nl[7:0];
  assign nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5279:5272]));
  assign MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5287:5280]));
  assign MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_563_nl = (readslicef_15_8_7(MultLoop_660_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_661_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_563_nl = nl_MultLoop_acc_563_nl[7:0];
  assign nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5295:5288]));
  assign MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5303:5296]));
  assign MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_562_nl = (readslicef_15_8_7(MultLoop_662_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_663_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_562_nl = nl_MultLoop_acc_562_nl[7:0];
  assign nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5343:5336]));
  assign MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5351:5344]));
  assign MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_559_nl = (readslicef_15_8_7(MultLoop_668_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_669_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_559_nl = nl_MultLoop_acc_559_nl[7:0];
  assign nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5359:5352]));
  assign MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5367:5360]));
  assign MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_558_nl = (readslicef_15_8_7(MultLoop_670_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_671_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_558_nl = nl_MultLoop_acc_558_nl[7:0];
  assign nl_MultLoop_acc_628_nl = MultLoop_acc_561_nl + MultLoop_acc_560_nl + MultLoop_acc_565_nl
      + MultLoop_acc_564_nl + MultLoop_acc_563_nl + MultLoop_acc_562_nl + MultLoop_acc_559_nl
      + MultLoop_acc_558_nl;
  assign MultLoop_acc_628_nl = nl_MultLoop_acc_628_nl[7:0];
  assign nl_MultLoop_acc_633_nl = MultLoop_acc_629_nl + MultLoop_acc_628_nl;
  assign MultLoop_acc_633_nl = nl_MultLoop_acc_633_nl[7:0];
  assign nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5375:5368]));
  assign MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5383:5376]));
  assign MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_557_nl = (readslicef_15_8_7(MultLoop_672_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_673_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_557_nl = nl_MultLoop_acc_557_nl[7:0];
  assign nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5391:5384]));
  assign MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5399:5392]));
  assign MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_556_nl = (readslicef_15_8_7(MultLoop_674_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_675_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_556_nl = nl_MultLoop_acc_556_nl[7:0];
  assign nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5407:5400]));
  assign MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5415:5408]));
  assign MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_555_nl = (readslicef_15_8_7(MultLoop_676_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_677_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_555_nl = nl_MultLoop_acc_555_nl[7:0];
  assign nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5423:5416]));
  assign MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5431:5424]));
  assign MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_554_nl = (readslicef_15_8_7(MultLoop_678_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_679_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_554_nl = nl_MultLoop_acc_554_nl[7:0];
  assign nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5439:5432]));
  assign MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5447:5440]));
  assign MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_553_nl = (readslicef_15_8_7(MultLoop_680_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_681_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_553_nl = nl_MultLoop_acc_553_nl[7:0];
  assign nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5455:5448]));
  assign MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5463:5456]));
  assign MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_552_nl = (readslicef_15_8_7(MultLoop_682_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_683_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_552_nl = nl_MultLoop_acc_552_nl[7:0];
  assign nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5471:5464]));
  assign MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5479:5472]));
  assign MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_551_nl = (readslicef_15_8_7(MultLoop_684_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_685_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_551_nl = nl_MultLoop_acc_551_nl[7:0];
  assign nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5487:5480]));
  assign MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5495:5488]));
  assign MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_550_nl = (readslicef_15_8_7(MultLoop_686_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_687_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_550_nl = nl_MultLoop_acc_550_nl[7:0];
  assign nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5567:5560]));
  assign MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5575:5568]));
  assign MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_545_nl = (readslicef_15_8_7(MultLoop_696_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_697_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_545_nl = nl_MultLoop_acc_545_nl[7:0];
  assign nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5583:5576]));
  assign MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5591:5584]));
  assign MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_544_nl = (readslicef_15_8_7(MultLoop_698_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_699_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_544_nl = nl_MultLoop_acc_544_nl[7:0];
  assign nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5599:5592]));
  assign MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5607:5600]));
  assign MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_543_nl = (readslicef_15_8_7(MultLoop_700_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_701_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_543_nl = nl_MultLoop_acc_543_nl[7:0];
  assign nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5615:5608]));
  assign MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5623:5616]));
  assign MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_542_nl = (readslicef_15_8_7(MultLoop_702_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_703_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_542_nl = nl_MultLoop_acc_542_nl[7:0];
  assign nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5503:5496]));
  assign MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5511:5504]));
  assign MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_549_nl = (readslicef_15_8_7(MultLoop_688_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_689_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_549_nl = nl_MultLoop_acc_549_nl[7:0];
  assign nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5519:5512]));
  assign MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5527:5520]));
  assign MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_548_nl = (readslicef_15_8_7(MultLoop_690_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_691_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_548_nl = nl_MultLoop_acc_548_nl[7:0];
  assign nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5535:5528]));
  assign MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5543:5536]));
  assign MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_547_nl = (readslicef_15_8_7(MultLoop_692_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_693_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_547_nl = nl_MultLoop_acc_547_nl[7:0];
  assign nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5551:5544]));
  assign MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5559:5552]));
  assign MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_546_nl = (readslicef_15_8_7(MultLoop_694_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_695_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_546_nl = nl_MultLoop_acc_546_nl[7:0];
  assign nl_MultLoop_acc_632_nl = MultLoop_acc_557_nl + MultLoop_acc_556_nl + MultLoop_acc_555_nl
      + MultLoop_acc_554_nl + MultLoop_acc_553_nl + MultLoop_acc_552_nl + MultLoop_acc_551_nl
      + MultLoop_acc_550_nl + MultLoop_acc_545_nl + MultLoop_acc_544_nl + MultLoop_acc_543_nl
      + MultLoop_acc_542_nl + MultLoop_acc_549_nl + MultLoop_acc_548_nl + MultLoop_acc_547_nl
      + MultLoop_acc_546_nl;
  assign MultLoop_acc_632_nl = nl_MultLoop_acc_632_nl[7:0];
  assign nl_MultLoop_acc_635_nl = MultLoop_acc_633_nl + MultLoop_acc_632_nl;
  assign MultLoop_acc_635_nl = nl_MultLoop_acc_635_nl[7:0];
  assign nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5695:5688]));
  assign MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5703:5696]));
  assign MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_537_nl = (readslicef_15_8_7(MultLoop_712_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_713_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_537_nl = nl_MultLoop_acc_537_nl[7:0];
  assign nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5711:5704]));
  assign MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5719:5712]));
  assign MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_536_nl = (readslicef_15_8_7(MultLoop_714_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_715_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_536_nl = nl_MultLoop_acc_536_nl[7:0];
  assign nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5823:5816]));
  assign MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5831:5824]));
  assign MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_529_nl = (readslicef_15_8_7(MultLoop_728_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_729_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_529_nl = nl_MultLoop_acc_529_nl[7:0];
  assign nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5839:5832]));
  assign MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5847:5840]));
  assign MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_528_nl = (readslicef_15_8_7(MultLoop_730_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_731_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_528_nl = nl_MultLoop_acc_528_nl[7:0];
  assign nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5759:5752]));
  assign MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5767:5760]));
  assign MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_533_nl = (readslicef_15_8_7(MultLoop_720_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_721_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_533_nl = nl_MultLoop_acc_533_nl[7:0];
  assign nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5775:5768]));
  assign MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5783:5776]));
  assign MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_532_nl = (readslicef_15_8_7(MultLoop_722_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_723_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_532_nl = nl_MultLoop_acc_532_nl[7:0];
  assign nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6079:6072]));
  assign MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6087:6080]));
  assign MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_513_nl = (readslicef_15_8_7(MultLoop_760_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_761_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_513_nl = nl_MultLoop_acc_513_nl[7:0];
  assign nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6095:6088]));
  assign MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6103:6096]));
  assign MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_512_nl = (readslicef_15_8_7(MultLoop_762_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_763_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_512_nl = nl_MultLoop_acc_512_nl[7:0];
  assign nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6015:6008]));
  assign MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6023:6016]));
  assign MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_517_nl = (readslicef_15_8_7(MultLoop_752_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_753_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_517_nl = nl_MultLoop_acc_517_nl[7:0];
  assign nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6031:6024]));
  assign MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6039:6032]));
  assign MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_516_nl = (readslicef_15_8_7(MultLoop_754_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_755_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_516_nl = nl_MultLoop_acc_516_nl[7:0];
  assign nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6047:6040]));
  assign MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6055:6048]));
  assign MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_515_nl = (readslicef_15_8_7(MultLoop_756_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_757_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_515_nl = nl_MultLoop_acc_515_nl[7:0];
  assign nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6063:6056]));
  assign MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6071:6064]));
  assign MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_514_nl = (readslicef_15_8_7(MultLoop_758_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_759_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_514_nl = nl_MultLoop_acc_514_nl[7:0];
  assign nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5887:5880]));
  assign MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5895:5888]));
  assign MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_525_nl = (readslicef_15_8_7(MultLoop_736_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_737_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_525_nl = nl_MultLoop_acc_525_nl[7:0];
  assign nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5903:5896]));
  assign MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5911:5904]));
  assign MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_524_nl = (readslicef_15_8_7(MultLoop_738_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_524_nl = nl_MultLoop_acc_524_nl[7:0];
  assign nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5919:5912]));
  assign MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5927:5920]));
  assign MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_523_nl = (readslicef_15_8_7(MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_741_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_523_nl = nl_MultLoop_acc_523_nl[7:0];
  assign nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5935:5928]));
  assign MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5943:5936]));
  assign MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_522_nl = (readslicef_15_8_7(MultLoop_742_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_743_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_522_nl = nl_MultLoop_acc_522_nl[7:0];
  assign nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5951:5944]));
  assign MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5959:5952]));
  assign MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_521_nl = (readslicef_15_8_7(MultLoop_744_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_745_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_521_nl = nl_MultLoop_acc_521_nl[7:0];
  assign nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5967:5960]));
  assign MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5975:5968]));
  assign MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_520_nl = (readslicef_15_8_7(MultLoop_746_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_747_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_520_nl = nl_MultLoop_acc_520_nl[7:0];
  assign nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5983:5976]));
  assign MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5991:5984]));
  assign MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_519_nl = (readslicef_15_8_7(MultLoop_748_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_749_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_519_nl = nl_MultLoop_acc_519_nl[7:0];
  assign nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5999:5992]));
  assign MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6007:6000]));
  assign MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_518_nl = (readslicef_15_8_7(MultLoop_750_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_751_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_518_nl = nl_MultLoop_acc_518_nl[7:0];
  assign nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5631:5624]));
  assign MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5639:5632]));
  assign MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_541_nl = (readslicef_15_8_7(MultLoop_704_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_541_nl = nl_MultLoop_acc_541_nl[7:0];
  assign nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5647:5640]));
  assign MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5655:5648]));
  assign MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_540_nl = (readslicef_15_8_7(MultLoop_706_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_707_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_540_nl = nl_MultLoop_acc_540_nl[7:0];
  assign nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5663:5656]));
  assign MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5671:5664]));
  assign MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_539_nl = (readslicef_15_8_7(MultLoop_708_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_709_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_539_nl = nl_MultLoop_acc_539_nl[7:0];
  assign nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5679:5672]));
  assign MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5687:5680]));
  assign MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_538_nl = (readslicef_15_8_7(MultLoop_710_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_711_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_538_nl = nl_MultLoop_acc_538_nl[7:0];
  assign nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5727:5720]));
  assign MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5735:5728]));
  assign MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_535_nl = (readslicef_15_8_7(MultLoop_716_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_717_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_535_nl = nl_MultLoop_acc_535_nl[7:0];
  assign nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5743:5736]));
  assign MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5751:5744]));
  assign MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_534_nl = (readslicef_15_8_7(MultLoop_718_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_719_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_534_nl = nl_MultLoop_acc_534_nl[7:0];
  assign nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5791:5784]));
  assign MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5799:5792]));
  assign MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_531_nl = (readslicef_15_8_7(MultLoop_724_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_725_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_531_nl = nl_MultLoop_acc_531_nl[7:0];
  assign nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5807:5800]));
  assign MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5815:5808]));
  assign MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_530_nl = (readslicef_15_8_7(MultLoop_726_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_727_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_530_nl = nl_MultLoop_acc_530_nl[7:0];
  assign nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5855:5848]));
  assign MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5863:5856]));
  assign MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_527_nl = (readslicef_15_8_7(MultLoop_732_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_733_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_527_nl = nl_MultLoop_acc_527_nl[7:0];
  assign nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5871:5864]));
  assign MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[5879:5872]));
  assign MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_526_nl = (readslicef_15_8_7(MultLoop_734_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_735_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_526_nl = nl_MultLoop_acc_526_nl[7:0];
  assign nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6111:6104]));
  assign MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6119:6112]));
  assign MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_511_nl = (readslicef_15_8_7(MultLoop_764_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_765_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_511_nl = nl_MultLoop_acc_511_nl[7:0];
  assign nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6127:6120]));
  assign MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_7_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1))
      * $signed((w4_rsci_idat_mxwt[6135:6128]));
  assign MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[14:0];
  assign nl_MultLoop_acc_510_nl = (readslicef_15_8_7(MultLoop_766_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl))
      + (readslicef_15_8_7(MultLoop_767_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign MultLoop_acc_510_nl = nl_MultLoop_acc_510_nl[7:0];
  assign nl_MultLoop_acc_634_nl = MultLoop_acc_537_nl + MultLoop_acc_536_nl + MultLoop_acc_529_nl
      + MultLoop_acc_528_nl + MultLoop_acc_533_nl + MultLoop_acc_532_nl + MultLoop_acc_513_nl
      + MultLoop_acc_512_nl + MultLoop_acc_517_nl + MultLoop_acc_516_nl + MultLoop_acc_515_nl
      + MultLoop_acc_514_nl + MultLoop_acc_525_nl + MultLoop_acc_524_nl + MultLoop_acc_523_nl
      + MultLoop_acc_522_nl + MultLoop_acc_521_nl + MultLoop_acc_520_nl + MultLoop_acc_519_nl
      + MultLoop_acc_518_nl + MultLoop_acc_541_nl + MultLoop_acc_540_nl + MultLoop_acc_539_nl
      + MultLoop_acc_538_nl + MultLoop_acc_535_nl + MultLoop_acc_534_nl + MultLoop_acc_531_nl
      + MultLoop_acc_530_nl + MultLoop_acc_527_nl + MultLoop_acc_526_nl + MultLoop_acc_511_nl
      + MultLoop_acc_510_nl;
  assign MultLoop_acc_634_nl = nl_MultLoop_acc_634_nl[7:0];
  assign nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1 = MultLoop_acc_635_nl
      + MultLoop_acc_634_nl;
  assign nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1 = nl_nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1[7:0];
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_85_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_86_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_86_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_87_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_87_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_88_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_89_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_90_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_91_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_92_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_101_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_107_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_108_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_108_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, (AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[6:0]),
      (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2262_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_2262_nl = nl_AccumDotWidth_acc_2262_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2262_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2251_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_2251_nl = nl_AccumDotWidth_acc_2251_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2251_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2240_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_2240_nl = nl_AccumDotWidth_acc_2240_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2240_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2229_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_2229_nl = nl_AccumDotWidth_acc_2229_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2229_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2218_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_2218_nl = nl_AccumDotWidth_acc_2218_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2218_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2207_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_2207_nl = nl_AccumDotWidth_acc_2207_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2207_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2196_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_2196_nl = nl_AccumDotWidth_acc_2196_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2196_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2185_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_2185_nl = nl_AccumDotWidth_acc_2185_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2185_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2168_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_2168_nl = nl_AccumDotWidth_acc_2168_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2168_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2151_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_2151_nl = nl_AccumDotWidth_acc_2151_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2151_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2134_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_2134_nl = nl_AccumDotWidth_acc_2134_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2134_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2117_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_2117_nl = nl_AccumDotWidth_acc_2117_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2117_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2100_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_2100_nl = nl_AccumDotWidth_acc_2100_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2100_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2083_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_2083_nl = nl_AccumDotWidth_acc_2083_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2083_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2066_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_2066_nl = nl_AccumDotWidth_acc_2066_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2066_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2049_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_2049_nl = nl_AccumDotWidth_acc_2049_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2049_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2032_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_2032_nl = nl_AccumDotWidth_acc_2032_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2032_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_2015_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_2015_nl = nl_AccumDotWidth_acc_2015_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_2015_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1998_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1998_nl = nl_AccumDotWidth_acc_1998_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1998_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1981_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1981_nl = nl_AccumDotWidth_acc_1981_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1981_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1964_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1964_nl = nl_AccumDotWidth_acc_1964_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1964_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1947_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1947_nl = nl_AccumDotWidth_acc_1947_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1947_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1930_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1930_nl = nl_AccumDotWidth_acc_1930_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1930_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1913_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1913_nl = nl_AccumDotWidth_acc_1913_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1913_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1902_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1902_nl = nl_AccumDotWidth_acc_1902_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1902_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1891_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1891_nl = nl_AccumDotWidth_acc_1891_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1891_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1880_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1880_nl = nl_AccumDotWidth_acc_1880_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1880_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1869_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1869_nl = nl_AccumDotWidth_acc_1869_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1869_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1858_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1858_nl = nl_AccumDotWidth_acc_1858_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1858_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1847_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1847_nl = nl_AccumDotWidth_acc_1847_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1847_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1836_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1836_nl = nl_AccumDotWidth_acc_1836_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1836_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1825_nl = (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1825_nl = nl_AccumDotWidth_acc_1825_nl[7:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1825_nl + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_4_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_4_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1808_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1808_nl = nl_AccumDotWidth_acc_1808_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1808_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1791_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1791_nl = nl_AccumDotWidth_acc_1791_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1791_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1774_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1774_nl = nl_AccumDotWidth_acc_1774_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1774_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1757_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1757_nl = nl_AccumDotWidth_acc_1757_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1757_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1740_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1740_nl = nl_AccumDotWidth_acc_1740_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1740_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1723_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1723_nl = nl_AccumDotWidth_acc_1723_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1723_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1706_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1706_nl = nl_AccumDotWidth_acc_1706_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1706_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1689_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1689_nl = nl_AccumDotWidth_acc_1689_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1689_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_4_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1663_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1663_nl = nl_AccumDotWidth_acc_1663_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1663_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1637_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1637_nl = nl_AccumDotWidth_acc_1637_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1637_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1611_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1611_nl = nl_AccumDotWidth_acc_1611_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1611_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1585_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1585_nl = nl_AccumDotWidth_acc_1585_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1585_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1559_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1559_nl = nl_AccumDotWidth_acc_1559_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1559_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1533_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1533_nl = nl_AccumDotWidth_acc_1533_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1533_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1507_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1507_nl = nl_AccumDotWidth_acc_1507_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1507_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[367:360])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[375:368])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[383:376])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1481_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1481_nl = nl_AccumDotWidth_acc_1481_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1481_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1455_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1455_nl = nl_AccumDotWidth_acc_1455_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1455_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1429_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1429_nl = nl_AccumDotWidth_acc_1429_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1429_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1403_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1403_nl = nl_AccumDotWidth_acc_1403_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1403_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1377_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1377_nl = nl_AccumDotWidth_acc_1377_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1377_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1351_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1351_nl = nl_AccumDotWidth_acc_1351_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1351_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1325_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1325_nl = nl_AccumDotWidth_acc_1325_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1325_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1299_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1299_nl = nl_AccumDotWidth_acc_1299_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1299_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[343:336])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[351:344])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[359:352])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1273_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1273_nl = nl_AccumDotWidth_acc_1273_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_1273_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_2_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1256_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1256_nl = nl_AccumDotWidth_acc_1256_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1256_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_8_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1239_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1239_nl = nl_AccumDotWidth_acc_1239_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1239_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_7_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1222_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1222_nl = nl_AccumDotWidth_acc_1222_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1222_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_6_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1205_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1205_nl = nl_AccumDotWidth_acc_1205_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1205_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_5_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1188_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1188_nl = nl_AccumDotWidth_acc_1188_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1188_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_4_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1171_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1171_nl = nl_AccumDotWidth_acc_1171_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1171_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_3_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1154_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1154_nl = nl_AccumDotWidth_acc_1154_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1154_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[335:328])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1137_nl = (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1137_nl = nl_AccumDotWidth_acc_1137_nl[7:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[295:288])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[303:296])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[327:320])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[319:312])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[311:304])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = AccumDotWidth_acc_1137_nl + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_1_AccumFilt_1_AccumDotWidth_acc_ncse_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1120_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_1120_nl = nl_AccumDotWidth_acc_1120_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1 = AccumDotWidth_acc_1120_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_63_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1103_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_1103_nl = nl_AccumDotWidth_acc_1103_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1 = AccumDotWidth_acc_1103_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_62_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1086_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_1086_nl = nl_AccumDotWidth_acc_1086_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1 = AccumDotWidth_acc_1086_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_61_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1069_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_1069_nl = nl_AccumDotWidth_acc_1069_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = AccumDotWidth_acc_1069_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1052_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_1052_nl = nl_AccumDotWidth_acc_1052_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = AccumDotWidth_acc_1052_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1035_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_1035_nl = nl_AccumDotWidth_acc_1035_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1 = AccumDotWidth_acc_1035_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_58_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1018_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_1018_nl = nl_AccumDotWidth_acc_1018_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1 = AccumDotWidth_acc_1018_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_57_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_1001_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_1001_nl = nl_AccumDotWidth_acc_1001_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1 = AccumDotWidth_acc_1001_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_56_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_975_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_975_nl = nl_AccumDotWidth_acc_975_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_975_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_55_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_949_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_949_nl = nl_AccumDotWidth_acc_949_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_949_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_54_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_923_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_923_nl = nl_AccumDotWidth_acc_923_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_923_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_53_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_897_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_897_nl = nl_AccumDotWidth_acc_897_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_897_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_52_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_871_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_871_nl = nl_AccumDotWidth_acc_871_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_871_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_51_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_845_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_845_nl = nl_AccumDotWidth_acc_845_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_845_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_50_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_819_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_819_nl = nl_AccumDotWidth_acc_819_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_819_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_49_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[271:264])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[279:272])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[287:280])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_793_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_793_nl = nl_AccumDotWidth_acc_793_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_793_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_48_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[127:120]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[63:56]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_767_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_767_nl = nl_AccumDotWidth_acc_767_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[191:184]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_767_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_47_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[119:112]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[55:48]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_741_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_741_nl = nl_AccumDotWidth_acc_741_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[183:176]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_741_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_46_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[111:104]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[47:40]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_715_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_715_nl = nl_AccumDotWidth_acc_715_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[175:168]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_715_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_45_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[103:96]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[39:32]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_689_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_689_nl = nl_AccumDotWidth_acc_689_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[167:160]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_689_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_44_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[95:88]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[31:24]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_663_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_663_nl = nl_AccumDotWidth_acc_663_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[159:152]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_663_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_43_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[87:80]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[23:16]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_637_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_637_nl = nl_AccumDotWidth_acc_637_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[151:144]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_637_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_42_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[79:72]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[15:8]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_611_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_611_nl = nl_AccumDotWidth_acc_611_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[143:136]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_611_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_41_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[247:240])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[71:64]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[255:248])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[7:0]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[263:256])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_585_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_585_nl = nl_AccumDotWidth_acc_585_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[135:128]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1 = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + AccumDotWidth_acc_585_nl + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_40_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_568_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_568_nl = nl_AccumDotWidth_acc_568_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[255:248]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[447:440]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[383:376]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[319:312]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[511:504]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[575:568]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1 = AccumDotWidth_acc_568_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_39_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_551_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_551_nl = nl_AccumDotWidth_acc_551_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[247:240]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[439:432]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[375:368]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[311:304]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[503:496]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[567:560]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1 = AccumDotWidth_acc_551_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_38_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_534_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_534_nl = nl_AccumDotWidth_acc_534_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[239:232]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[431:424]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[367:360]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[303:296]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[495:488]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[559:552]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1 = AccumDotWidth_acc_534_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_37_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_517_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_517_nl = nl_AccumDotWidth_acc_517_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[231:224]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[423:416]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[359:352]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[295:288]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[487:480]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[551:544]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1 = AccumDotWidth_acc_517_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_36_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_500_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_500_nl = nl_AccumDotWidth_acc_500_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[223:216]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[415:408]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[351:344]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[287:280]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[479:472]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[543:536]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1 = AccumDotWidth_acc_500_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_35_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_483_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_483_nl = nl_AccumDotWidth_acc_483_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[215:208]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[407:400]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[343:336]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[279:272]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[471:464]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[535:528]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1 = AccumDotWidth_acc_483_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_34_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_466_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_466_nl = nl_AccumDotWidth_acc_466_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[207:200]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[399:392]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[335:328]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[271:264]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[463:456]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[527:520]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1 = AccumDotWidth_acc_466_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_33_sva_1[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[239:232])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_449_nl = (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_449_nl = nl_AccumDotWidth_acc_449_nl[7:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[199:192]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[391:384]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[199:192])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[207:200])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[231:224])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[327:320]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[223:216])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[263:256]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[455:448]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[519:512]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[215:208])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1 = AccumDotWidth_acc_449_nl
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_1_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_2_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_32_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_438_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_438_nl = nl_AccumDotWidth_acc_438_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1 = AccumDotWidth_acc_438_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_31_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_427_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_427_nl = nl_AccumDotWidth_acc_427_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1 = AccumDotWidth_acc_427_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_30_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_416_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_416_nl = nl_AccumDotWidth_acc_416_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1 = AccumDotWidth_acc_416_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_29_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_405_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_405_nl = nl_AccumDotWidth_acc_405_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1 = AccumDotWidth_acc_405_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_28_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_394_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_394_nl = nl_AccumDotWidth_acc_394_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1 = AccumDotWidth_acc_394_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_27_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_383_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_383_nl = nl_AccumDotWidth_acc_383_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1 = AccumDotWidth_acc_383_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_26_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_372_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_372_nl = nl_AccumDotWidth_acc_372_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1 = AccumDotWidth_acc_372_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_25_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_361_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_361_nl = nl_AccumDotWidth_acc_361_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1 = AccumDotWidth_acc_361_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_4_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_24_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_344_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_344_nl = nl_AccumDotWidth_acc_344_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1 = AccumDotWidth_acc_344_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_23_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_327_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_327_nl = nl_AccumDotWidth_acc_327_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1 = AccumDotWidth_acc_327_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_22_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_310_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_310_nl = nl_AccumDotWidth_acc_310_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1 = AccumDotWidth_acc_310_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_21_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_293_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_293_nl = nl_AccumDotWidth_acc_293_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1 = AccumDotWidth_acc_293_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_20_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_276_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_276_nl = nl_AccumDotWidth_acc_276_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1 = AccumDotWidth_acc_276_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_19_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_259_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_259_nl = nl_AccumDotWidth_acc_259_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1 = AccumDotWidth_acc_259_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_18_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_242_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_242_nl = nl_AccumDotWidth_acc_242_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1 = AccumDotWidth_acc_242_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_17_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[191:184])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_225_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_225_nl = nl_AccumDotWidth_acc_225_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[79:72])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[183:176])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[175:168])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[87:80])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[95:88])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1 = AccumDotWidth_acc_225_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_16_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_208_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_208_nl = nl_AccumDotWidth_acc_208_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[639:632]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1215:1208]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1279:1272]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[767:760]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[703:696]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1343:1336]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1 = AccumDotWidth_acc_208_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_15_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_191_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_191_nl = nl_AccumDotWidth_acc_191_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[631:624]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1207:1200]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1271:1264]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[759:752]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[695:688]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1335:1328]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1 = AccumDotWidth_acc_191_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_14_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_174_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_174_nl = nl_AccumDotWidth_acc_174_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[623:616]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1199:1192]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1263:1256]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[751:744]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[687:680]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1327:1320]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1 = AccumDotWidth_acc_174_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_13_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_157_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_157_nl = nl_AccumDotWidth_acc_157_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[615:608]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1191:1184]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1255:1248]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[743:736]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[679:672]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1319:1312]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1 = AccumDotWidth_acc_157_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_12_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_140_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_140_nl = nl_AccumDotWidth_acc_140_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[607:600]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1183:1176]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1247:1240]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[735:728]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[671:664]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1311:1304]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1 = AccumDotWidth_acc_140_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_11_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_123_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_123_nl = nl_AccumDotWidth_acc_123_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[599:592]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1175:1168]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1239:1232]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[727:720]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[663:656]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1303:1296]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1 = AccumDotWidth_acc_123_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_10_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_106_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_106_nl = nl_AccumDotWidth_acc_106_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[591:584]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1167:1160]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1231:1224]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[719:712]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[655:648]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1295:1288]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1 = AccumDotWidth_acc_106_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_9_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[167:160])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_89_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_89_nl = nl_AccumDotWidth_acc_89_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[583:576]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[55:48])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1159:1152]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1223:1216]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[159:152])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[711:704]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[151:144])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[647:640]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[63:56])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[71:64])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1287:1280]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1 = AccumDotWidth_acc_89_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_1_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_2_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_8_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1727:1720]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_78_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[55:49]);
  assign AccumDotWidth_acc_78_nl = nl_AccumDotWidth_acc_78_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[831:824]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1599:1592]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[895:888]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1087:1080]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1471:1464]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1663:1656]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[959:952]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1151:1144]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1535:1528]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[1023:1016]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1407:1400]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1 = AccumDotWidth_acc_78_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_8_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_7_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1719:1712]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_67_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[48:42]);
  assign AccumDotWidth_acc_67_nl = nl_AccumDotWidth_acc_67_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[823:816]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1591:1584]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[887:880]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1079:1072]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1463:1456]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1655:1648]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[951:944]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1143:1136]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1527:1520]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[1015:1008]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1399:1392]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1 = AccumDotWidth_acc_67_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_6_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1711:1704]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_56_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[41:35]);
  assign AccumDotWidth_acc_56_nl = nl_AccumDotWidth_acc_56_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[815:808]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1583:1576]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[879:872]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1071:1064]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1455:1448]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1647:1640]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[943:936]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1135:1128]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1519:1512]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[1007:1000]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1391:1384]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1 = AccumDotWidth_acc_56_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_5_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1703:1696]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_45_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[34:28]);
  assign AccumDotWidth_acc_45_nl = nl_AccumDotWidth_acc_45_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[807:800]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1575:1568]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[871:864]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1063:1056]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1447:1440]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1639:1632]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[935:928]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1127:1120]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1511:1504]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[999:992]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1383:1376]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1 = AccumDotWidth_acc_45_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_5_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_4_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1695:1688]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_34_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[27:21]);
  assign AccumDotWidth_acc_34_nl = nl_AccumDotWidth_acc_34_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[799:792]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1567:1560]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[863:856]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1055:1048]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1439:1432]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1631:1624]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[927:920]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1119:1112]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1503:1496]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[991:984]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1375:1368]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1 = AccumDotWidth_acc_34_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_4_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_3_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1687:1680]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_23_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[20:14]);
  assign AccumDotWidth_acc_23_nl = nl_AccumDotWidth_acc_23_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[791:784]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1559:1552]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[855:848]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1047:1040]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1431:1424]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1623:1616]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[919:912]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1111:1104]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1495:1488]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[983:976]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1367:1360]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1 = AccumDotWidth_acc_23_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_2_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1679:1672]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_12_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[13:7]);
  assign AccumDotWidth_acc_12_nl = nl_AccumDotWidth_acc_12_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[783:776]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1551:1544]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[847:840]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1039:1032]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1423:1416]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1615:1608]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[911:904]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1103:1096]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1487:1480]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[975:968]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1359:1352]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1 = AccumDotWidth_acc_12_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_1_sva_1[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[143:136])) * $signed((w2_rsci_idat_mxwt[1671:1664]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_AccumDotWidth_acc_7_nl = (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + conv_s2s_7_8(b2_rsci_idat_mxwt[6:0]);
  assign AccumDotWidth_acc_7_nl = nl_AccumDotWidth_acc_7_nl[7:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[7:0])) * $signed((w2_rsci_idat_mxwt[775:768]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[127:120])) * $signed((w2_rsci_idat_mxwt[1543:1536]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[15:8])) * $signed((w2_rsci_idat_mxwt[839:832]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[39:32])) * $signed((w2_rsci_idat_mxwt[1031:1024]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[111:104])) * $signed((w2_rsci_idat_mxwt[1415:1408]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[135:128])) * $signed((w2_rsci_idat_mxwt[1607:1600]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[23:16])) * $signed((w2_rsci_idat_mxwt[903:896]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[47:40])) * $signed((w2_rsci_idat_mxwt[1095:1088]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[119:112])) * $signed((w2_rsci_idat_mxwt[1479:1472]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[31:24])) * $signed((w2_rsci_idat_mxwt[967:960]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl[14:0];
  assign nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = $signed((input_1_rsci_idat_mxwt[103:96])) * $signed((w2_rsci_idat_mxwt[1351:1344]));
  assign ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl
      = nl_ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl[14:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1 = AccumDotWidth_acc_7_nl
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_2_ConvFiltHeight_3_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_3_else_mul_nl))
      + (readslicef_15_8_7(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_1_ConvChan_1_ConvFiltHeight_3_ConvFiltWidth_2_else_mul_nl));
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1[7:0];
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_8_9(nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl[8:0];
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_asn_1289 = MUX_v_7_2_2(7'b0000000,
      (nnet_conv_2d_input_t_layer2_t_config2_acc_0_sva_1[6:0]), (readslicef_9_1_8(nnet_relu_layer2_t_layer3_t_relu_config3_for_1_operator_8_2_true_AC_TRN_AC_WRAP_acc_nl)));
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_idat_6_0 <= 7'b0000000;
      layer5_out_rsci_idat_14_8 <= 7'b0000000;
      layer5_out_rsci_idat_22_16 <= 7'b0000000;
      layer5_out_rsci_idat_30_24 <= 7'b0000000;
      layer5_out_rsci_idat_38_32 <= 7'b0000000;
      layer5_out_rsci_idat_46_40 <= 7'b0000000;
      layer5_out_rsci_idat_54_48 <= 7'b0000000;
      layer5_out_rsci_idat_62_56 <= 7'b0000000;
      layer5_out_rsci_idat_70_64 <= 7'b0000000;
      layer5_out_rsci_idat_78_72 <= 7'b0000000;
    end
    else if ( nnet_relu_layer4_t_result_t_relu_config5_for_if_and_cse ) begin
      layer5_out_rsci_idat_6_0 <= MUX_v_7_2_2(7'b0000000, (layer4_out_0_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_14_8 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_22_16 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_30_24 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_38_32 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_46_40 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_54_48 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_62_56 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_70_64 <= MUX_v_7_2_2(7'b0000000, (nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
      layer5_out_rsci_idat_78_72 <= MUX_v_7_2_2(7'b0000000, (MultLoop_1280_MultLoop_acc_3_ncse_sva_1[6:0]),
          (readslicef_9_1_8(nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl)));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= 1'b1;
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= fsm_output[1];
    end
  end
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(layer4_out_0_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_1_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_2_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_3_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_4_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_5_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_6_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_7_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_7_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_8_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(nnet_dense_large_rf_leq_nin_layer3_t_layer4_t_config4_acc_8_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_8_9(MultLoop_1280_MultLoop_acc_3_ncse_sva_1);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_8_2_true_AC_TRN_AC_WRAP_1_acc_nl[8:0];

  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] readslicef_15_8_7;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_15_8_7 = tmp[7:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] conv_s2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10
// ------------------------------------------------------------------


module econ_4x4_d10 (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_rdy, input_1_rsc_triosy_lz,
      layer5_out_rsc_dat, layer5_out_rsc_vld, layer5_out_rsc_rdy, layer5_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_rdy,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_rdy, const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld,
      w2_rsc_rdy, w2_rsc_triosy_lz, b2_rsc_dat, b2_rsc_vld, b2_rsc_rdy, b2_rsc_triosy_lz,
      w4_rsc_dat, w4_rsc_vld, w4_rsc_rdy, w4_rsc_triosy_lz, b4_rsc_dat, b4_rsc_vld,
      b4_rsc_rdy, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [383:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_rdy;
  output input_1_rsc_triosy_lz;
  output [79:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input layer5_out_rsc_rdy;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input const_size_in_1_rsc_rdy;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input const_size_out_1_rsc_rdy;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_rdy;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_rdy;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_rdy;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_rdy;
  output b4_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  econ_4x4_d10_core econ_4x4_d10_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_rdy(input_1_rsc_rdy),
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_rdy(layer5_out_rsc_rdy),
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_rdy(const_size_in_1_rsc_rdy),
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_rdy(const_size_out_1_rsc_rdy),
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_rdy(w2_rsc_rdy),
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_rdy(b2_rsc_rdy),
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_rdy(w4_rsc_rdy),
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_rdy(b4_rsc_rdy),
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz)
    );
endmodule



