
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_vld_v1 (dat, vld, idat, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             vld;
  input  [width-1:0] idat;
  input              ivld;

  wire   [width-1:0] dat;
  wire               vld;

  assign dat = idat;
  assign vld = ivld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> ../td_ccore_solutions/nnet__relu_layer6_t_result_t_relu_config7__34efe21f6655c9bfc003c946efcef06b7604_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 17:54:16 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer6_t_result_t_relu_config7_core
// ------------------------------------------------------------------


module nnet_relu_layer6_t_result_t_relu_config7_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [53:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [53:0] data_rsci_idat;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;

  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [53:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18 , 1'b0
      , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd20),
  .width(32'sd54)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd21),
  .width(32'sd54)) res_rsci (
      .d(nl_res_rsci_d[53:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer6_t_result_t_relu_config7
// ------------------------------------------------------------------


module nnet_relu_layer6_t_result_t_relu_config7 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [53:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer6_t_result_t_relu_config7_core nnet_relu_layer6_t_result_t_relu_config7_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_layer5_t_layer6_t_config6__84b33fe340531fb85f7e6289891f4e23dd66_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 17:54:46 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer5_t_layer6_t_config6_core
// ------------------------------------------------------------------


module nnet_dense_large_layer5_t_layer6_t_config6_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [107:0] data_rsci_idat;
  reg [17:0] res_rsci_d_53_36;
  wire [18:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [18:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [18:0] nl_res_rsci_d_17_0;
  wire [18:0] Result_acc_54_cse_1;
  wire [19:0] nl_Result_acc_54_cse_1;
  wire [14:0] Result_acc_15_itm_24_10;
  wire [13:0] Result_acc_21_itm_18_5;

  wire[17:0] MultLoop_acc_8_nl;
  wire[19:0] nl_MultLoop_acc_8_nl;
  wire[17:0] MultLoop_acc_6_nl;
  wire[18:0] nl_MultLoop_acc_6_nl;
  wire[22:0] Result_acc_30_nl;
  wire[23:0] nl_Result_acc_30_nl;
  wire[19:0] Result_acc_47_nl;
  wire[20:0] nl_Result_acc_47_nl;
  wire[17:0] Result_acc_46_nl;
  wire[18:0] nl_Result_acc_46_nl;
  wire[22:0] Result_acc_28_nl;
  wire[23:0] nl_Result_acc_28_nl;
  wire[20:0] Result_acc_32_nl;
  wire[21:0] nl_Result_acc_32_nl;
  wire[17:0] Result_acc_31_nl;
  wire[18:0] nl_Result_acc_31_nl;
  wire[17:0] Result_acc_76_nl;
  wire[18:0] nl_Result_acc_76_nl;
  wire[22:0] Result_acc_41_nl;
  wire[24:0] nl_Result_acc_41_nl;
  wire[10:0] Result_acc_75_nl;
  wire[11:0] nl_Result_acc_75_nl;
  wire[13:0] MultLoop_acc_19_nl;
  wire[14:0] nl_MultLoop_acc_19_nl;
  wire[17:0] MultLoop_acc_7_nl;
  wire[18:0] nl_MultLoop_acc_7_nl;
  wire[17:0] Result_acc_79_nl;
  wire[18:0] nl_Result_acc_79_nl;
  wire[18:0] Result_acc_78_nl;
  wire[19:0] nl_Result_acc_78_nl;
  wire[23:0] Result_acc_35_nl;
  wire[25:0] nl_Result_acc_35_nl;
  wire[8:0] Result_acc_77_nl;
  wire[9:0] nl_Result_acc_77_nl;
  wire[24:0] Result_acc_29_nl;
  wire[25:0] nl_Result_acc_29_nl;
  wire[22:0] Result_acc_45_nl;
  wire[24:0] nl_Result_acc_45_nl;
  wire[17:0] Result_acc_43_nl;
  wire[18:0] nl_Result_acc_43_nl;
  wire[10:0] Result_acc_80_nl;
  wire[11:0] nl_Result_acc_80_nl;
  wire[17:0] MultLoop_acc_18_nl;
  wire[19:0] nl_MultLoop_acc_18_nl;
  wire[24:0] Result_acc_2_nl;
  wire[25:0] nl_Result_acc_2_nl;
  wire[22:0] Result_acc_61_nl;
  wire[23:0] nl_Result_acc_61_nl;
  wire[17:0] Result_acc_nl;
  wire[18:0] nl_Result_acc_nl;
  wire[21:0] Result_acc_60_nl;
  wire[23:0] nl_Result_acc_60_nl;
  wire[17:0] Result_acc_58_nl;
  wire[18:0] nl_Result_acc_58_nl;
  wire[10:0] Result_acc_72_nl;
  wire[11:0] nl_Result_acc_72_nl;
  wire[15:0] MultLoop_acc_15_nl;
  wire[16:0] nl_MultLoop_acc_15_nl;
  wire[24:0] Result_acc_3_nl;
  wire[26:0] nl_Result_acc_3_nl;
  wire[12:0] Result_acc_73_nl;
  wire[13:0] nl_Result_acc_73_nl;
  wire[11:0] MultLoop_acc_14_nl;
  wire[12:0] nl_MultLoop_acc_14_nl;
  wire[17:0] MultLoop_acc_17_nl;
  wire[18:0] nl_MultLoop_acc_17_nl;
  wire[24:0] Result_acc_19_nl;
  wire[25:0] nl_Result_acc_19_nl;
  wire[22:0] Result_acc_66_nl;
  wire[24:0] nl_Result_acc_66_nl;
  wire[18:0] Result_acc_74_nl;
  wire[19:0] nl_Result_acc_74_nl;
  wire[22:0] Result_acc_69_nl;
  wire[24:0] nl_Result_acc_69_nl;
  wire[17:0] Result_acc_67_nl;
  wire[18:0] nl_Result_acc_67_nl;
  wire[17:0] MultLoop_acc_13_nl;
  wire[18:0] nl_MultLoop_acc_13_nl;
  wire[17:0] MultLoop_acc_11_nl;
  wire[18:0] nl_MultLoop_acc_11_nl;
  wire[20:0] Result_acc_26_nl;
  wire[21:0] nl_Result_acc_26_nl;
  wire[17:0] Result_acc_56_nl;
  wire[18:0] nl_Result_acc_56_nl;
  wire[14:0] MultLoop_acc_10_nl;
  wire[15:0] nl_MultLoop_acc_10_nl;
  wire[13:0] MultLoop_acc_9_nl;
  wire[14:0] nl_MultLoop_acc_9_nl;
  wire[21:0] Result_acc_23_nl;
  wire[22:0] nl_Result_acc_23_nl;
  wire[18:0] Result_acc_51_nl;
  wire[19:0] nl_Result_acc_51_nl;
  wire[25:0] Result_acc_22_nl;
  wire[26:0] nl_Result_acc_22_nl;
  wire[22:0] Result_acc_50_nl;
  wire[24:0] nl_Result_acc_50_nl;
  wire[9:0] Result_acc_70_nl;
  wire[10:0] nl_Result_acc_70_nl;
  wire[17:0] MultLoop_acc_12_nl;
  wire[18:0] nl_MultLoop_acc_12_nl;
  wire[17:0] Result_acc_71_nl;
  wire[18:0] nl_Result_acc_71_nl;
  wire[20:0] Result_acc_53_nl;
  wire[21:0] nl_Result_acc_53_nl;
  wire[17:0] Result_acc_52_nl;
  wire[18:0] nl_Result_acc_52_nl;
  wire[21:0] Result_acc_25_nl;
  wire[22:0] nl_Result_acc_25_nl;
  wire[19:0] Result_acc_55_nl;
  wire[20:0] nl_Result_acc_55_nl;
  wire[24:0] Result_acc_15_nl;
  wire[26:0] nl_Result_acc_15_nl;
  wire[19:0] Result_acc_37_nl;
  wire[20:0] nl_Result_acc_37_nl;
  wire[18:0] Result_acc_21_nl;
  wire[19:0] nl_Result_acc_21_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [53:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_53_36 , res_rsci_d_35_18 , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd15),
  .width(32'sd108)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd16),
  .width(32'sd54)) res_rsci (
      .d(nl_res_rsci_d[53:0]),
      .z(res_rsc_z)
    );
  assign nl_Result_acc_37_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[53:36]));
  assign Result_acc_37_nl = nl_Result_acc_37_nl[19:0];
  assign nl_Result_acc_15_nl = conv_s2s_24_25({(data_rsci_idat[53:36]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[53:36]) , 4'b0000}) + conv_s2s_20_25(Result_acc_37_nl);
  assign Result_acc_15_nl = nl_Result_acc_15_nl[24:0];
  assign Result_acc_15_itm_24_10 = readslicef_25_15_10((Result_acc_15_nl));
  assign nl_Result_acc_21_nl = conv_s2u_16_19(data_rsci_idat[107:92]) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign Result_acc_21_nl = nl_Result_acc_21_nl[18:0];
  assign Result_acc_21_itm_18_5 = readslicef_19_14_5((Result_acc_21_nl));
  assign nl_Result_acc_54_cse_1 = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_15_19(data_rsci_idat[71:57]);
  assign Result_acc_54_cse_1 = nl_Result_acc_54_cse_1[18:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_53_36 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
    end
  end
  assign nl_Result_acc_46_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_13_18(data_rsci_idat[107:95]);
  assign Result_acc_46_nl = nl_Result_acc_46_nl[17:0];
  assign nl_Result_acc_47_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_18_20(Result_acc_46_nl);
  assign Result_acc_47_nl = nl_Result_acc_47_nl[19:0];
  assign nl_Result_acc_30_nl = conv_s2u_20_23(Result_acc_47_nl) + conv_s2u_22_23({(data_rsci_idat[107:90])
      , 4'b0000});
  assign Result_acc_30_nl = nl_Result_acc_30_nl[22:0];
  assign nl_Result_acc_31_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_14_18(data_rsci_idat[17:4]);
  assign Result_acc_31_nl = nl_Result_acc_31_nl[17:0];
  assign nl_Result_acc_32_nl = conv_s2s_20_21({(~ (data_rsci_idat[17:0])) , 2'b01})
      + conv_s2s_18_21(Result_acc_31_nl);
  assign Result_acc_32_nl = nl_Result_acc_32_nl[20:0];
  assign nl_Result_acc_28_nl = conv_s2u_21_23(Result_acc_32_nl) + ({(data_rsci_idat[17:0])
      , 5'b00100});
  assign Result_acc_28_nl = nl_Result_acc_28_nl[22:0];
  assign nl_MultLoop_acc_6_nl = (readslicef_23_18_5((Result_acc_30_nl))) + conv_s2s_17_18(readslicef_23_17_6((Result_acc_28_nl)));
  assign MultLoop_acc_6_nl = nl_MultLoop_acc_6_nl[17:0];
  assign nl_Result_acc_75_nl =  -conv_s2s_10_11(data_rsci_idat[71:62]);
  assign Result_acc_75_nl = nl_Result_acc_75_nl[10:0];
  assign nl_Result_acc_41_nl = ({(data_rsci_idat[71:54]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[71:54])) , 2'b01}) + conv_s2s_19_23({(Result_acc_75_nl) , (~
      (data_rsci_idat[61:54]))});
  assign Result_acc_41_nl = nl_Result_acc_41_nl[22:0];
  assign nl_Result_acc_76_nl = conv_s2u_15_18(readslicef_23_15_8((Result_acc_41_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign Result_acc_76_nl = nl_Result_acc_76_nl[17:0];
  assign nl_MultLoop_acc_19_nl = (Result_acc_15_itm_24_10[14:1]) + 14'b11111111011111;
  assign MultLoop_acc_19_nl = nl_MultLoop_acc_19_nl[13:0];
  assign nl_MultLoop_acc_8_nl = (MultLoop_acc_6_nl) + conv_s2s_17_18(readslicef_18_17_1((Result_acc_76_nl)))
      + conv_s2s_15_18({(MultLoop_acc_19_nl) , (Result_acc_15_itm_24_10[0])});
  assign MultLoop_acc_8_nl = nl_MultLoop_acc_8_nl[17:0];
  assign nl_Result_acc_77_nl =  -conv_s2s_8_9(data_rsci_idat[35:28]);
  assign Result_acc_77_nl = nl_Result_acc_77_nl[8:0];
  assign nl_Result_acc_35_nl = ({(data_rsci_idat[35:18]) , 6'b000100}) + conv_s2s_20_24({(~
      (data_rsci_idat[35:18])) , 2'b01}) + conv_s2s_19_24({(Result_acc_77_nl) , (~
      (data_rsci_idat[27:18]))});
  assign Result_acc_35_nl = nl_Result_acc_35_nl[23:0];
  assign nl_Result_acc_78_nl = conv_s2u_18_19(data_rsci_idat[35:18]) + conv_s2u_16_19(readslicef_24_16_8((Result_acc_35_nl)));
  assign Result_acc_78_nl = nl_Result_acc_78_nl[18:0];
  assign nl_Result_acc_79_nl = conv_s2u_17_18(readslicef_19_17_2((Result_acc_78_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign Result_acc_79_nl = nl_Result_acc_79_nl[17:0];
  assign nl_Result_acc_80_nl = conv_s2s_10_11(data_rsci_idat[89:80]) + 11'b00000000001;
  assign Result_acc_80_nl = nl_Result_acc_80_nl[10:0];
  assign nl_Result_acc_43_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_17_18({(Result_acc_80_nl)
      , (data_rsci_idat[79:74])});
  assign Result_acc_43_nl = nl_Result_acc_43_nl[17:0];
  assign nl_Result_acc_45_nl = conv_s2s_22_23({(~ (data_rsci_idat[89:72])) , 4'b0100})
      + conv_s2s_20_23({(~ (data_rsci_idat[89:72])) , 2'b01}) + conv_s2s_18_23(Result_acc_43_nl);
  assign Result_acc_45_nl = nl_Result_acc_45_nl[22:0];
  assign nl_Result_acc_29_nl = conv_s2u_23_25(Result_acc_45_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[89:72])) , 6'b010000});
  assign Result_acc_29_nl = nl_Result_acc_29_nl[24:0];
  assign nl_MultLoop_acc_7_nl = (Result_acc_79_nl) + (readslicef_25_18_7((Result_acc_29_nl)));
  assign MultLoop_acc_7_nl = nl_MultLoop_acc_7_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_8_nl) + (MultLoop_acc_7_nl);
  assign nl_Result_acc_61_nl = conv_s2s_22_23({(~ (data_rsci_idat[35:18])) , 4'b0001})
      + conv_s2s_18_23(~ (data_rsci_idat[35:18]));
  assign Result_acc_61_nl = nl_Result_acc_61_nl[22:0];
  assign nl_Result_acc_2_nl = conv_s2s_23_25(Result_acc_61_nl) + ({(data_rsci_idat[35:18])
      , 7'b0010000});
  assign Result_acc_2_nl = nl_Result_acc_2_nl[24:0];
  assign nl_Result_acc_72_nl = conv_s2s_10_11(data_rsci_idat[17:8]) + 11'b00000000001;
  assign Result_acc_72_nl = nl_Result_acc_72_nl[10:0];
  assign nl_Result_acc_58_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_17_18({(Result_acc_72_nl)
      , (data_rsci_idat[7:2])});
  assign Result_acc_58_nl = nl_Result_acc_58_nl[17:0];
  assign nl_Result_acc_60_nl = ({(data_rsci_idat[17:0]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[17:0])) , 2'b01}) + conv_s2s_18_22(Result_acc_58_nl);
  assign Result_acc_60_nl = nl_Result_acc_60_nl[21:0];
  assign nl_Result_acc_nl = conv_s2u_16_18(readslicef_22_16_6((Result_acc_60_nl)))
      + (~ (data_rsci_idat[17:0]));
  assign Result_acc_nl = nl_Result_acc_nl[17:0];
  assign nl_Result_acc_73_nl =  -conv_s2s_12_13(data_rsci_idat[53:42]);
  assign Result_acc_73_nl = nl_Result_acc_73_nl[12:0];
  assign nl_Result_acc_3_nl = conv_s2s_24_25({(~ (data_rsci_idat[53:36])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[53:36])) , 4'b0001}) + conv_s2s_19_25({(Result_acc_73_nl)
      , (~ (data_rsci_idat[41:36]))});
  assign Result_acc_3_nl = nl_Result_acc_3_nl[24:0];
  assign nl_MultLoop_acc_14_nl = conv_s2s_11_12(Result_acc_21_itm_18_5[13:3]) + 12'b000110111101;
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[11:0];
  assign nl_MultLoop_acc_15_nl = (readslicef_25_16_9((Result_acc_3_nl))) + conv_s2s_12_16(MultLoop_acc_14_nl);
  assign MultLoop_acc_15_nl = nl_MultLoop_acc_15_nl[15:0];
  assign nl_MultLoop_acc_18_nl = (readslicef_25_18_7((Result_acc_2_nl))) + conv_s2s_17_18(readslicef_18_17_1((Result_acc_nl)))
      + conv_s2s_16_18(MultLoop_acc_15_nl);
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[17:0];
  assign nl_Result_acc_66_nl = ({(~ (data_rsci_idat[71:54])) , 5'b00000}) + conv_s2s_21_23({(data_rsci_idat[71:54])
      , 3'b000}) + conv_s2s_19_23(Result_acc_54_cse_1);
  assign Result_acc_66_nl = nl_Result_acc_66_nl[22:0];
  assign nl_Result_acc_19_nl = conv_s2u_23_25(Result_acc_66_nl) + ({(data_rsci_idat[71:54])
      , 7'b0100000});
  assign Result_acc_19_nl = nl_Result_acc_19_nl[24:0];
  assign nl_Result_acc_67_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_16_18(data_rsci_idat[89:74]);
  assign Result_acc_67_nl = nl_Result_acc_67_nl[17:0];
  assign nl_Result_acc_69_nl = ({(data_rsci_idat[89:72]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[89:72])) , 3'b001}) + conv_s2s_18_23(Result_acc_67_nl);
  assign Result_acc_69_nl = nl_Result_acc_69_nl[22:0];
  assign nl_Result_acc_74_nl = conv_s2u_16_19(readslicef_23_16_7((Result_acc_69_nl)))
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign Result_acc_74_nl = nl_Result_acc_74_nl[18:0];
  assign nl_MultLoop_acc_17_nl = (readslicef_25_18_7((Result_acc_19_nl))) + (readslicef_19_18_1((Result_acc_74_nl)));
  assign MultLoop_acc_17_nl = nl_MultLoop_acc_17_nl[17:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_18_nl) + (MultLoop_acc_17_nl);
  assign nl_Result_acc_56_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_14_18(data_rsci_idat[89:76]);
  assign Result_acc_56_nl = nl_Result_acc_56_nl[17:0];
  assign nl_Result_acc_26_nl = conv_s2u_18_21(Result_acc_56_nl) + ({(data_rsci_idat[89:72])
      , 3'b001});
  assign Result_acc_26_nl = nl_Result_acc_26_nl[20:0];
  assign nl_MultLoop_acc_9_nl = Result_acc_21_itm_18_5 + 14'b11111110001111;
  assign MultLoop_acc_9_nl = nl_MultLoop_acc_9_nl[13:0];
  assign nl_Result_acc_51_nl = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_16_19(data_rsci_idat[35:20]);
  assign Result_acc_51_nl = nl_Result_acc_51_nl[18:0];
  assign nl_Result_acc_23_nl = conv_s2u_19_22(Result_acc_51_nl) + conv_s2u_21_22({(data_rsci_idat[35:18])
      , 3'b000});
  assign Result_acc_23_nl = nl_Result_acc_23_nl[21:0];
  assign nl_MultLoop_acc_10_nl = conv_s2s_14_15(MultLoop_acc_9_nl) + (readslicef_22_15_7((Result_acc_23_nl)));
  assign MultLoop_acc_10_nl = nl_MultLoop_acc_10_nl[14:0];
  assign nl_MultLoop_acc_11_nl = conv_s2s_17_18(readslicef_21_17_4((Result_acc_26_nl)))
      + conv_s2s_15_18(MultLoop_acc_10_nl);
  assign MultLoop_acc_11_nl = nl_MultLoop_acc_11_nl[17:0];
  assign nl_Result_acc_70_nl = conv_s2s_9_10(data_rsci_idat[17:9]) + 10'b0000000001;
  assign Result_acc_70_nl = nl_Result_acc_70_nl[9:0];
  assign nl_Result_acc_50_nl = ({(~ (data_rsci_idat[17:0])) , 5'b00000}) + conv_s2s_18_23(data_rsci_idat[17:0])
      + conv_s2s_17_23({(Result_acc_70_nl) , (data_rsci_idat[8:2])});
  assign Result_acc_50_nl = nl_Result_acc_50_nl[22:0];
  assign nl_Result_acc_22_nl = conv_s2u_23_26(Result_acc_50_nl) + conv_s2u_25_26({(~
      (data_rsci_idat[17:0])) , 7'b0100000});
  assign Result_acc_22_nl = nl_Result_acc_22_nl[25:0];
  assign nl_MultLoop_acc_13_nl = (MultLoop_acc_11_nl) + (readslicef_26_18_8((Result_acc_22_nl)));
  assign MultLoop_acc_13_nl = nl_MultLoop_acc_13_nl[17:0];
  assign nl_Result_acc_52_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_15_18(data_rsci_idat[53:39]);
  assign Result_acc_52_nl = nl_Result_acc_52_nl[17:0];
  assign nl_Result_acc_53_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_18_21(Result_acc_52_nl);
  assign Result_acc_53_nl = nl_Result_acc_53_nl[20:0];
  assign nl_Result_acc_71_nl = conv_s2u_15_18(readslicef_21_15_6((Result_acc_53_nl)))
      + (data_rsci_idat[53:36]);
  assign Result_acc_71_nl = nl_Result_acc_71_nl[17:0];
  assign nl_Result_acc_55_nl = ({(~ (data_rsci_idat[71:54])) , 2'b00}) + conv_s2s_19_20(Result_acc_54_cse_1);
  assign Result_acc_55_nl = nl_Result_acc_55_nl[19:0];
  assign nl_Result_acc_25_nl = conv_s2u_20_22(Result_acc_55_nl) + ({(data_rsci_idat[71:54])
      , 4'b0100});
  assign Result_acc_25_nl = nl_Result_acc_25_nl[21:0];
  assign nl_MultLoop_acc_12_nl = (Result_acc_71_nl) + conv_s2s_17_18(readslicef_22_17_5((Result_acc_25_nl)));
  assign MultLoop_acc_12_nl = nl_MultLoop_acc_12_nl[17:0];
  assign nl_res_rsci_d_35_18  = (MultLoop_acc_13_nl) + (MultLoop_acc_12_nl);

  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [13:0] readslicef_19_14_5;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_19_14_5 = tmp[13:0];
  end
  endfunction


  function automatic [16:0] readslicef_19_17_2;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_19_17_2 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [14:0] readslicef_21_15_6;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_21_15_6 = tmp[14:0];
  end
  endfunction


  function automatic [16:0] readslicef_21_17_4;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_21_17_4 = tmp[16:0];
  end
  endfunction


  function automatic [14:0] readslicef_22_15_7;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_22_15_7 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_22_16_6;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_22_16_6 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_22_17_5;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_22_17_5 = tmp[16:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_23_16_7;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_23_16_7 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_23_17_6;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_23_17_6 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_23_18_5;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_23_18_5 = tmp[17:0];
  end
  endfunction


  function automatic [15:0] readslicef_24_16_8;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_24_16_8 = tmp[15:0];
  end
  endfunction


  function automatic [14:0] readslicef_25_15_10;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_25_15_10 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_25_16_9;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_25_16_9 = tmp[15:0];
  end
  endfunction


  function automatic [17:0] readslicef_25_18_7;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_25_18_7 = tmp[17:0];
  end
  endfunction


  function automatic [17:0] readslicef_26_18_8;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_26_18_8 = tmp[17:0];
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_15 = {vector[13], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_17_23 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_23 = {{6{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_19_25 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_25 = {{6{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_23_26 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_26 = {{3{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2u_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2u_25_26 = {vector[24], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer5_t_layer6_t_config6
// ------------------------------------------------------------------


module nnet_dense_large_layer5_t_layer6_t_config6 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [53:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_layer5_t_layer6_t_config6_core nnet_dense_large_layer5_t_layer6_t_config6_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__relu_layer4_t_layer5_t_relu_config5__b4f43beadc57ef670128187311fd10ca9086_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 17:55:15 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer4_t_layer5_t_relu_config5_core
// ------------------------------------------------------------------


module nnet_relu_layer4_t_layer5_t_relu_config5_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [107:0] data_rsci_idat;
  reg [16:0] res_rsci_d_106_90;
  reg [16:0] res_rsci_d_88_72;
  reg [16:0] res_rsci_d_70_54;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;

  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [107:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_106_90 , 1'b0 , res_rsci_d_88_72 , 1'b0
      , res_rsci_d_70_54 , 1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18 , 1'b0
      , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd13),
  .width(32'sd108)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd14),
  .width(32'sd108)) res_rsci (
      .d(nl_res_rsci_d[107:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_106_90 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
      res_rsci_d_88_72 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_70_54 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_106_90 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[106:90]),
          (readslicef_19_1_18((for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_88_72 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[88:72]),
          (readslicef_19_1_18((for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_70_54 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[70:54]),
          (readslicef_19_1_18((for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[107:90]);
  assign for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[89:72]);
  assign for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[71:54]);
  assign for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer4_t_layer5_t_relu_config5
// ------------------------------------------------------------------


module nnet_relu_layer4_t_layer5_t_relu_config5 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [107:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer4_t_layer5_t_relu_config5_core nnet_relu_layer4_t_layer5_t_relu_config5_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_layer3_t_layer4_t_config4__d025c2976550a6e247a69155a3f8bdb2311e4_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 17:57:27 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4_core
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [431:0] data_rsci_idat;
  reg [17:0] res_rsci_d_107_90;
  wire [21:0] nl_res_rsci_d_107_90;
  reg [17:0] res_rsci_d_89_72;
  wire [20:0] nl_res_rsci_d_89_72;
  reg [17:0] res_rsci_d_71_54;
  wire [20:0] nl_res_rsci_d_71_54;
  reg [17:0] res_rsci_d_53_36;
  wire [20:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [20:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [20:0] nl_res_rsci_d_17_0;
  wire [17:0] MultLoop_acc_174_cse_1;
  wire [18:0] nl_MultLoop_acc_174_cse_1;
  wire [17:0] Result_acc_137_cse_1;
  wire [18:0] nl_Result_acc_137_cse_1;
  wire [18:0] Result_acc_131_cse_1;
  wire [19:0] nl_Result_acc_131_cse_1;
  wire [18:0] Result_acc_172_cse_1;
  wire [19:0] nl_Result_acc_172_cse_1;
  wire [19:0] MultLoop_acc_263_cse_1;
  wire [20:0] nl_MultLoop_acc_263_cse_1;
  wire [19:0] MultLoop_acc_76_cse_1;
  wire [20:0] nl_MultLoop_acc_76_cse_1;
  wire [19:0] MultLoop_acc_193_cse_1;
  wire [20:0] nl_MultLoop_acc_193_cse_1;
  wire [19:0] MultLoop_acc_395;
  wire [20:0] nl_MultLoop_acc_395;
  wire [12:0] MultLoop_MultLoop_conc_50_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_50_18_6;
  wire [16:0] MultLoop_acc_106_itm_22_6;
  wire [12:0] Result_acc_43_itm_17_5;
  wire [16:0] MultLoop_acc_72_itm_23_7;
  wire [16:0] MultLoop_acc_54_itm_21_5;

  wire[17:0] MultLoop_acc_139_nl;
  wire[20:0] nl_MultLoop_acc_139_nl;
  wire[24:0] Result_acc_84_nl;
  wire[25:0] nl_Result_acc_84_nl;
  wire[21:0] Result_acc_111_nl;
  wire[22:0] nl_Result_acc_111_nl;
  wire[19:0] Result_acc_110_nl;
  wire[20:0] nl_Result_acc_110_nl;
  wire[26:0] Result_acc_62_nl;
  wire[27:0] nl_Result_acc_62_nl;
  wire[24:0] Result_acc_113_nl;
  wire[26:0] nl_Result_acc_113_nl;
  wire[21:0] Result_acc_83_nl;
  wire[22:0] nl_Result_acc_83_nl;
  wire[17:0] Result_acc_100_nl;
  wire[18:0] nl_Result_acc_100_nl;
  wire[17:0] Result_acc_218_nl;
  wire[18:0] nl_Result_acc_218_nl;
  wire[23:0] Result_acc_103_nl;
  wire[25:0] nl_Result_acc_103_nl;
  wire[10:0] Result_acc_217_nl;
  wire[11:0] nl_Result_acc_217_nl;
  wire[17:0] Result_acc_220_nl;
  wire[18:0] nl_Result_acc_220_nl;
  wire[22:0] Result_acc_107_nl;
  wire[24:0] nl_Result_acc_107_nl;
  wire[10:0] Result_acc_219_nl;
  wire[11:0] nl_Result_acc_219_nl;
  wire[23:0] Result_acc_57_nl;
  wire[24:0] nl_Result_acc_57_nl;
  wire[21:0] Result_acc_88_nl;
  wire[22:0] nl_Result_acc_88_nl;
  wire[20:0] Result_acc_59_nl;
  wire[21:0] nl_Result_acc_59_nl;
  wire[18:0] Result_acc_90_nl;
  wire[19:0] nl_Result_acc_90_nl;
  wire[12:0] Result_acc_221_nl;
  wire[13:0] nl_Result_acc_221_nl;
  wire[17:0] MultLoop_acc_138_nl;
  wire[19:0] nl_MultLoop_acc_138_nl;
  wire[25:0] Result_acc_63_nl;
  wire[27:0] nl_Result_acc_63_nl;
  wire[11:0] Result_acc_223_nl;
  wire[12:0] nl_Result_acc_223_nl;
  wire[22:0] Result_acc_85_nl;
  wire[23:0] nl_Result_acc_85_nl;
  wire[17:0] Result_acc_117_nl;
  wire[18:0] nl_Result_acc_117_nl;
  wire[11:0] Result_acc_224_nl;
  wire[12:0] nl_Result_acc_224_nl;
  wire[17:0] Result_acc_226_nl;
  wire[18:0] nl_Result_acc_226_nl;
  wire[24:0] Result_acc_121_nl;
  wire[26:0] nl_Result_acc_121_nl;
  wire[19:0] Result_acc_119_nl;
  wire[20:0] nl_Result_acc_119_nl;
  wire[9:0] Result_acc_225_nl;
  wire[10:0] nl_Result_acc_225_nl;
  wire[20:0] Result_acc_229_nl;
  wire[21:0] nl_Result_acc_229_nl;
  wire[17:0] Result_acc_228_nl;
  wire[18:0] nl_Result_acc_228_nl;
  wire[20:0] Result_acc_123_nl;
  wire[21:0] nl_Result_acc_123_nl;
  wire[10:0] Result_acc_227_nl;
  wire[11:0] nl_Result_acc_227_nl;
  wire[22:0] Result_acc_82_nl;
  wire[23:0] nl_Result_acc_82_nl;
  wire[20:0] Result_acc_96_nl;
  wire[21:0] nl_Result_acc_96_nl;
  wire[24:0] Result_acc_65_nl;
  wire[26:0] nl_Result_acc_65_nl;
  wire[12:0] Result_acc_232_nl;
  wire[13:0] nl_Result_acc_232_nl;
  wire[18:0] Result_acc_230_nl;
  wire[19:0] nl_Result_acc_230_nl;
  wire[21:0] Result_acc_125_nl;
  wire[22:0] nl_Result_acc_125_nl;
  wire[26:0] Result_acc_74_nl;
  wire[27:0] nl_Result_acc_74_nl;
  wire[24:0] Result_acc_127_nl;
  wire[26:0] nl_Result_acc_127_nl;
  wire[23:0] Result_acc_86_nl;
  wire[24:0] nl_Result_acc_86_nl;
  wire[21:0] Result_acc_130_nl;
  wire[23:0] nl_Result_acc_130_nl;
  wire[17:0] Result_acc_73_nl;
  wire[18:0] nl_Result_acc_73_nl;
  wire[23:0] Result_acc_72_nl;
  wire[24:0] nl_Result_acc_72_nl;
  wire[20:0] Result_acc_91_nl;
  wire[21:0] nl_Result_acc_91_nl;
  wire[22:0] Result_acc_80_nl;
  wire[23:0] nl_Result_acc_80_nl;
  wire[20:0] Result_acc_94_nl;
  wire[21:0] nl_Result_acc_94_nl;
  wire[17:0] Result_acc_93_nl;
  wire[18:0] nl_Result_acc_93_nl;
  wire[12:0] Result_acc_231_nl;
  wire[13:0] nl_Result_acc_231_nl;
  wire[19:0] Result_acc_79_nl;
  wire[20:0] nl_Result_acc_79_nl;
  wire[11:0] MultLoop_acc_119_nl;
  wire[12:0] nl_MultLoop_acc_119_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl;
  wire[17:0] Result_acc_77_nl;
  wire[18:0] nl_Result_acc_77_nl;
  wire[17:0] MultLoop_acc_340_nl;
  wire[21:0] nl_MultLoop_acc_340_nl;
  wire[24:0] MultLoop_acc_97_nl;
  wire[25:0] nl_MultLoop_acc_97_nl;
  wire[22:0] MultLoop_acc_292_nl;
  wire[24:0] nl_MultLoop_acc_292_nl;
  wire[22:0] MultLoop_acc_90_nl;
  wire[23:0] nl_MultLoop_acc_90_nl;
  wire[20:0] MultLoop_acc_289_nl;
  wire[22:0] nl_MultLoop_acc_289_nl;
  wire[22:0] MultLoop_acc_28_nl;
  wire[23:0] nl_MultLoop_acc_28_nl;
  wire[21:0] MultLoop_acc_286_nl;
  wire[23:0] nl_MultLoop_acc_286_nl;
  wire[10:0] MultLoop_acc_375_nl;
  wire[11:0] nl_MultLoop_acc_375_nl;
  wire[18:0] MultLoop_acc_396_nl;
  wire[19:0] nl_MultLoop_acc_396_nl;
  wire[23:0] MultLoop_acc_14_nl;
  wire[24:0] nl_MultLoop_acc_14_nl;
  wire[20:0] MultLoop_acc_283_nl;
  wire[21:0] nl_MultLoop_acc_283_nl;
  wire[18:0] MultLoop_acc_96_nl;
  wire[19:0] nl_MultLoop_acc_96_nl;
  wire[18:0] MultLoop_acc_376_nl;
  wire[19:0] nl_MultLoop_acc_376_nl;
  wire[19:0] MultLoop_acc_287_nl;
  wire[20:0] nl_MultLoop_acc_287_nl;
  wire[17:0] MultLoop_acc_378_nl;
  wire[18:0] nl_MultLoop_acc_378_nl;
  wire[19:0] MultLoop_acc_279_nl;
  wire[20:0] nl_MultLoop_acc_279_nl;
  wire[20:0] MultLoop_acc_9_nl;
  wire[21:0] nl_MultLoop_acc_9_nl;
  wire[18:0] MultLoop_acc_277_nl;
  wire[19:0] nl_MultLoop_acc_277_nl;
  wire[13:0] MultLoop_acc_379_nl;
  wire[14:0] nl_MultLoop_acc_379_nl;
  wire[17:0] MultLoop_acc_339_nl;
  wire[19:0] nl_MultLoop_acc_339_nl;
  wire[18:0] MultLoop_acc_380_nl;
  wire[19:0] nl_MultLoop_acc_380_nl;
  wire[22:0] MultLoop_acc_293_nl;
  wire[23:0] nl_MultLoop_acc_293_nl;
  wire[19:0] MultLoop_acc_381_nl;
  wire[20:0] nl_MultLoop_acc_381_nl;
  wire[25:0] MultLoop_acc_295_nl;
  wire[27:0] nl_MultLoop_acc_295_nl;
  wire[24:0] MultLoop_acc_95_nl;
  wire[25:0] nl_MultLoop_acc_95_nl;
  wire[22:0] MultLoop_acc_298_nl;
  wire[23:0] nl_MultLoop_acc_298_nl;
  wire[19:0] MultLoop_acc_297_nl;
  wire[20:0] nl_MultLoop_acc_297_nl;
  wire[17:0] MultLoop_acc_296_nl;
  wire[18:0] nl_MultLoop_acc_296_nl;
  wire[17:0] MultLoop_acc_384_nl;
  wire[18:0] nl_MultLoop_acc_384_nl;
  wire[18:0] MultLoop_acc_383_nl;
  wire[19:0] nl_MultLoop_acc_383_nl;
  wire[23:0] MultLoop_acc_301_nl;
  wire[24:0] nl_MultLoop_acc_301_nl;
  wire[20:0] MultLoop_acc_300_nl;
  wire[21:0] nl_MultLoop_acc_300_nl;
  wire[9:0] MultLoop_acc_382_nl;
  wire[10:0] nl_MultLoop_acc_382_nl;
  wire[17:0] MultLoop_acc_337_nl;
  wire[20:0] nl_MultLoop_acc_337_nl;
  wire[23:0] MultLoop_acc_92_nl;
  wire[24:0] nl_MultLoop_acc_92_nl;
  wire[21:0] MultLoop_acc_314_nl;
  wire[23:0] nl_MultLoop_acc_314_nl;
  wire[24:0] MultLoop_acc_91_nl;
  wire[25:0] nl_MultLoop_acc_91_nl;
  wire[23:0] MultLoop_acc_316_nl;
  wire[24:0] nl_MultLoop_acc_316_nl;
  wire[17:0] MultLoop_acc_315_nl;
  wire[18:0] nl_MultLoop_acc_315_nl;
  wire[16:0] MultLoop_3_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_3_MultLoop_acc_3_nl;
  wire[16:0] MultLoop_acc_322_nl;
  wire[18:0] nl_MultLoop_acc_322_nl;
  wire[19:0] MultLoop_acc_7_nl;
  wire[20:0] nl_MultLoop_acc_7_nl;
  wire[18:0] MultLoop_acc_318_nl;
  wire[19:0] nl_MultLoop_acc_318_nl;
  wire[11:0] MultLoop_acc_390_nl;
  wire[12:0] nl_MultLoop_acc_390_nl;
  wire[18:0] MultLoop_acc_89_nl;
  wire[19:0] nl_MultLoop_acc_89_nl;
  wire[22:0] MultLoop_acc_6_nl;
  wire[23:0] nl_MultLoop_acc_6_nl;
  wire[17:0] MultLoop_acc_320_nl;
  wire[18:0] nl_MultLoop_acc_320_nl;
  wire[12:0] MultLoop_acc_391_nl;
  wire[13:0] nl_MultLoop_acc_391_nl;
  wire[17:0] MultLoop_acc_23_nl;
  wire[18:0] nl_MultLoop_acc_23_nl;
  wire[23:0] MultLoop_acc_21_nl;
  wire[25:0] nl_MultLoop_acc_21_nl;
  wire[13:0] MultLoop_acc_392_nl;
  wire[14:0] nl_MultLoop_acc_392_nl;
  wire[17:0] MultLoop_acc_386_nl;
  wire[18:0] nl_MultLoop_acc_386_nl;
  wire[22:0] MultLoop_acc_305_nl;
  wire[23:0] nl_MultLoop_acc_305_nl;
  wire[19:0] MultLoop_acc_304_nl;
  wire[20:0] nl_MultLoop_acc_304_nl;
  wire[12:0] MultLoop_acc_385_nl;
  wire[13:0] nl_MultLoop_acc_385_nl;
  wire[23:0] MultLoop_acc_94_nl;
  wire[24:0] nl_MultLoop_acc_94_nl;
  wire[17:0] MultLoop_acc_307_nl;
  wire[18:0] nl_MultLoop_acc_307_nl;
  wire[10:0] MultLoop_acc_387_nl;
  wire[11:0] nl_MultLoop_acc_387_nl;
  wire[17:0] MultLoop_acc_389_nl;
  wire[18:0] nl_MultLoop_acc_389_nl;
  wire[22:0] MultLoop_acc_310_nl;
  wire[24:0] nl_MultLoop_acc_310_nl;
  wire[10:0] MultLoop_acc_388_nl;
  wire[11:0] nl_MultLoop_acc_388_nl;
  wire[24:0] MultLoop_acc_93_nl;
  wire[25:0] nl_MultLoop_acc_93_nl;
  wire[20:0] MultLoop_acc_312_nl;
  wire[22:0] nl_MultLoop_acc_312_nl;
  wire[17:0] MultLoop_acc_162_nl;
  wire[20:0] nl_MultLoop_acc_162_nl;
  wire[17:0] MultLoop_acc_158_nl;
  wire[20:0] nl_MultLoop_acc_158_nl;
  wire[19:0] Result_acc_56_nl;
  wire[20:0] nl_Result_acc_56_nl;
  wire[17:0] Result_acc_169_nl;
  wire[18:0] nl_Result_acc_169_nl;
  wire[18:0] Result_acc_48_nl;
  wire[19:0] nl_Result_acc_48_nl;
  wire[24:0] Result_acc_32_nl;
  wire[25:0] nl_Result_acc_32_nl;
  wire[20:0] Result_acc_134_nl;
  wire[21:0] nl_Result_acc_134_nl;
  wire[24:0] Result_acc_29_nl;
  wire[26:0] nl_Result_acc_29_nl;
  wire[12:0] Result_acc_204_nl;
  wire[13:0] nl_Result_acc_204_nl;
  wire[18:0] Result_acc_233_nl;
  wire[19:0] nl_Result_acc_233_nl;
  wire[20:0] Result_acc_42_nl;
  wire[21:0] nl_Result_acc_42_nl;
  wire[18:0] Result_acc_136_nl;
  wire[19:0] nl_Result_acc_136_nl;
  wire[12:0] Result_acc_205_nl;
  wire[13:0] nl_Result_acc_205_nl;
  wire[12:0] MultLoop_acc_374_nl;
  wire[13:0] nl_MultLoop_acc_374_nl;
  wire[22:0] Result_acc_49_nl;
  wire[23:0] nl_Result_acc_49_nl;
  wire[21:0] Result_acc_138_nl;
  wire[22:0] nl_Result_acc_138_nl;
  wire[18:0] Result_acc_234_nl;
  wire[19:0] nl_Result_acc_234_nl;
  wire[22:0] Result_acc_37_nl;
  wire[23:0] nl_Result_acc_37_nl;
  wire[20:0] Result_acc_142_nl;
  wire[22:0] nl_Result_acc_142_nl;
  wire[11:0] Result_acc_206_nl;
  wire[12:0] nl_Result_acc_206_nl;
  wire[22:0] Result_acc_51_nl;
  wire[23:0] nl_Result_acc_51_nl;
  wire[20:0] Result_acc_144_nl;
  wire[21:0] nl_Result_acc_144_nl;
  wire[17:0] Result_acc_143_nl;
  wire[18:0] nl_Result_acc_143_nl;
  wire[17:0] MultLoop_acc_161_nl;
  wire[19:0] nl_MultLoop_acc_161_nl;
  wire[25:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl;
  wire[27:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl;
  wire[12:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl;
  wire[18:0] Result_acc_207_nl;
  wire[19:0] nl_Result_acc_207_nl;
  wire[21:0] Result_acc_145_nl;
  wire[22:0] nl_Result_acc_145_nl;
  wire[22:0] Result_acc_52_nl;
  wire[23:0] nl_Result_acc_52_nl;
  wire[17:0] Result_acc_147_nl;
  wire[18:0] nl_Result_acc_147_nl;
  wire[11:0] Result_acc_208_nl;
  wire[12:0] nl_Result_acc_208_nl;
  wire[19:0] Result_acc_209_nl;
  wire[20:0] nl_Result_acc_209_nl;
  wire[25:0] Result_acc_150_nl;
  wire[26:0] nl_Result_acc_150_nl;
  wire[22:0] Result_acc_149_nl;
  wire[23:0] nl_Result_acc_149_nl;
  wire[19:0] Result_acc_148_nl;
  wire[20:0] nl_Result_acc_148_nl;
  wire[17:0] MultLoop_acc_159_nl;
  wire[19:0] nl_MultLoop_acc_159_nl;
  wire[20:0] Result_acc_54_nl;
  wire[21:0] nl_Result_acc_54_nl;
  wire[18:0] Result_acc_160_nl;
  wire[19:0] nl_Result_acc_160_nl;
  wire[17:0] Result_acc_214_nl;
  wire[18:0] nl_Result_acc_214_nl;
  wire[22:0] Result_acc_163_nl;
  wire[24:0] nl_Result_acc_163_nl;
  wire[9:0] Result_acc_213_nl;
  wire[10:0] nl_Result_acc_213_nl;
  wire[22:0] Result_acc_41_nl;
  wire[23:0] nl_Result_acc_41_nl;
  wire[20:0] Result_acc_166_nl;
  wire[21:0] nl_Result_acc_166_nl;
  wire[17:0] Result_acc_165_nl;
  wire[18:0] nl_Result_acc_165_nl;
  wire[9:0] Result_acc_215_nl;
  wire[10:0] nl_Result_acc_215_nl;
  wire[21:0] Result_acc_55_nl;
  wire[22:0] nl_Result_acc_55_nl;
  wire[17:0] Result_acc_168_nl;
  wire[18:0] nl_Result_acc_168_nl;
  wire[13:0] Result_acc_216_nl;
  wire[14:0] nl_Result_acc_216_nl;
  wire[23:0] Result_acc_53_nl;
  wire[24:0] nl_Result_acc_53_nl;
  wire[20:0] Result_acc_152_nl;
  wire[21:0] nl_Result_acc_152_nl;
  wire[17:0] Result_acc_151_nl;
  wire[18:0] nl_Result_acc_151_nl;
  wire[17:0] Result_acc_211_nl;
  wire[18:0] nl_Result_acc_211_nl;
  wire[22:0] Result_acc_156_nl;
  wire[24:0] nl_Result_acc_156_nl;
  wire[9:0] Result_acc_210_nl;
  wire[10:0] nl_Result_acc_210_nl;
  wire[18:0] Result_acc_212_nl;
  wire[19:0] nl_Result_acc_212_nl;
  wire[18:0] Result_acc_235_nl;
  wire[19:0] nl_Result_acc_235_nl;
  wire[22:0] Result_acc_38_nl;
  wire[23:0] nl_Result_acc_38_nl;
  wire[19:0] Result_acc_159_nl;
  wire[20:0] nl_Result_acc_159_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl;
  wire[21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl;
  wire[18:0] MultLoop_acc_368_nl;
  wire[19:0] nl_MultLoop_acc_368_nl;
  wire[21:0] MultLoop_acc_101_nl;
  wire[22:0] nl_MultLoop_acc_101_nl;
  wire[17:0] MultLoop_acc_253_nl;
  wire[18:0] nl_MultLoop_acc_253_nl;
  wire[13:0] MultLoop_acc_369_nl;
  wire[14:0] nl_MultLoop_acc_369_nl;
  wire[24:0] MultLoop_acc_35_nl;
  wire[25:0] nl_MultLoop_acc_35_nl;
  wire[21:0] MultLoop_acc_243_nl;
  wire[22:0] nl_MultLoop_acc_243_nl;
  wire[17:0] MultLoop_acc_366_nl;
  wire[18:0] nl_MultLoop_acc_366_nl;
  wire[19:0] MultLoop_acc_245_nl;
  wire[20:0] nl_MultLoop_acc_245_nl;
  wire[12:0] MultLoop_acc_365_nl;
  wire[13:0] nl_MultLoop_acc_365_nl;
  wire[24:0] MultLoop_acc_50_nl;
  wire[25:0] nl_MultLoop_acc_50_nl;
  wire[21:0] MultLoop_acc_247_nl;
  wire[22:0] nl_MultLoop_acc_247_nl;
  wire[23:0] MultLoop_acc_104_nl;
  wire[24:0] nl_MultLoop_acc_104_nl;
  wire[17:0] MultLoop_acc_249_nl;
  wire[18:0] nl_MultLoop_acc_249_nl;
  wire[11:0] MultLoop_acc_367_nl;
  wire[12:0] nl_MultLoop_acc_367_nl;
  wire[25:0] MultLoop_acc_41_nl;
  wire[26:0] nl_MultLoop_acc_41_nl;
  wire[20:0] MultLoop_acc_254_nl;
  wire[21:0] nl_MultLoop_acc_254_nl;
  wire[25:0] MultLoop_acc_38_nl;
  wire[27:0] nl_MultLoop_acc_38_nl;
  wire[11:0] MultLoop_acc_370_nl;
  wire[12:0] nl_MultLoop_acc_370_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl;
  wire[24:0] MultLoop_acc_48_nl;
  wire[25:0] nl_MultLoop_acc_48_nl;
  wire[22:0] MultLoop_acc_258_nl;
  wire[23:0] nl_MultLoop_acc_258_nl;
  wire[20:0] MultLoop_acc_257_nl;
  wire[21:0] nl_MultLoop_acc_257_nl;
  wire[23:0] MultLoop_acc_45_nl;
  wire[24:0] nl_MultLoop_acc_45_nl;
  wire[21:0] MultLoop_acc_260_nl;
  wire[22:0] nl_MultLoop_acc_260_nl;
  wire[22:0] MultLoop_acc_103_nl;
  wire[23:0] nl_MultLoop_acc_103_nl;
  wire[19:0] MultLoop_acc_262_nl;
  wire[20:0] nl_MultLoop_acc_262_nl;
  wire[17:0] MultLoop_acc_261_nl;
  wire[18:0] nl_MultLoop_acc_261_nl;
  wire[22:0] MultLoop_acc_32_nl;
  wire[23:0] nl_MultLoop_acc_32_nl;
  wire[21:0] MultLoop_acc_105_nl;
  wire[22:0] nl_MultLoop_acc_105_nl;
  wire[18:0] MultLoop_acc_242_nl;
  wire[19:0] nl_MultLoop_acc_242_nl;
  wire[12:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl;
  wire[14:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl;
  wire[10:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl;
  wire[12:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl;
  wire[18:0] MultLoop_acc_102_nl;
  wire[19:0] nl_MultLoop_acc_102_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl;
  wire[26:0] MultLoop_acc_36_nl;
  wire[27:0] nl_MultLoop_acc_36_nl;
  wire[24:0] MultLoop_acc_272_nl;
  wire[25:0] nl_MultLoop_acc_272_nl;
  wire[22:0] MultLoop_acc_98_nl;
  wire[23:0] nl_MultLoop_acc_98_nl;
  wire[20:0] MultLoop_acc_275_nl;
  wire[21:0] nl_MultLoop_acc_275_nl;
  wire[17:0] MultLoop_acc_274_nl;
  wire[18:0] nl_MultLoop_acc_274_nl;
  wire[12:0] MultLoop_acc_373_nl;
  wire[13:0] nl_MultLoop_acc_373_nl;
  wire[18:0] MultLoop_acc_99_nl;
  wire[19:0] nl_MultLoop_acc_99_nl;
  wire[26:0] MultLoop_acc_42_nl;
  wire[27:0] nl_MultLoop_acc_42_nl;
  wire[21:0] MultLoop_acc_264_nl;
  wire[22:0] nl_MultLoop_acc_264_nl;
  wire[22:0] MultLoop_acc_100_nl;
  wire[23:0] nl_MultLoop_acc_100_nl;
  wire[20:0] MultLoop_acc_266_nl;
  wire[22:0] nl_MultLoop_acc_266_nl;
  wire[25:0] MultLoop_acc_40_nl;
  wire[27:0] nl_MultLoop_acc_40_nl;
  wire[11:0] MultLoop_acc_371_nl;
  wire[12:0] nl_MultLoop_acc_371_nl;
  wire[18:0] MultLoop_acc_372_nl;
  wire[19:0] nl_MultLoop_acc_372_nl;
  wire[23:0] MultLoop_acc_271_nl;
  wire[24:0] nl_MultLoop_acc_271_nl;
  wire[21:0] MultLoop_acc_270_nl;
  wire[22:0] nl_MultLoop_acc_270_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl;
  wire[20:0] Result_acc_198_nl;
  wire[21:0] nl_Result_acc_198_nl;
  wire[17:0] Result_acc_197_nl;
  wire[18:0] nl_Result_acc_197_nl;
  wire[19:0] Result_acc_194_nl;
  wire[20:0] nl_Result_acc_194_nl;
  wire[9:0] Result_acc_196_nl;
  wire[10:0] nl_Result_acc_196_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[20:0] Result_acc_16_nl;
  wire[21:0] nl_Result_acc_16_nl;
  wire[18:0] Result_acc_171_nl;
  wire[19:0] nl_Result_acc_171_nl;
  wire[23:0] Result_acc_17_nl;
  wire[24:0] nl_Result_acc_17_nl;
  wire[20:0] Result_acc_173_nl;
  wire[21:0] nl_Result_acc_173_nl;
  wire[22:0] Result_acc_18_nl;
  wire[23:0] nl_Result_acc_18_nl;
  wire[20:0] Result_acc_175_nl;
  wire[22:0] nl_Result_acc_175_nl;
  wire[17:0] Result_acc_200_nl;
  wire[18:0] nl_Result_acc_200_nl;
  wire[23:0] Result_acc_178_nl;
  wire[24:0] nl_Result_acc_178_nl;
  wire[20:0] Result_acc_177_nl;
  wire[21:0] nl_Result_acc_177_nl;
  wire[11:0] Result_acc_199_nl;
  wire[12:0] nl_Result_acc_199_nl;
  wire[20:0] Result_acc_19_nl;
  wire[21:0] nl_Result_acc_19_nl;
  wire[17:0] Result_acc_179_nl;
  wire[18:0] nl_Result_acc_179_nl;
  wire[20:0] Result_acc_20_nl;
  wire[21:0] nl_Result_acc_20_nl;
  wire[18:0] Result_acc_180_nl;
  wire[19:0] nl_Result_acc_180_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl;
  wire[22:0] Result_acc_21_nl;
  wire[23:0] nl_Result_acc_21_nl;
  wire[18:0] Result_acc_181_nl;
  wire[19:0] nl_Result_acc_181_nl;
  wire[25:0] Result_acc_3_nl;
  wire[26:0] nl_Result_acc_3_nl;
  wire[22:0] Result_acc_183_nl;
  wire[24:0] nl_Result_acc_183_nl;
  wire[22:0] Result_acc_22_nl;
  wire[23:0] nl_Result_acc_22_nl;
  wire[21:0] Result_acc_185_nl;
  wire[22:0] nl_Result_acc_185_nl;
  wire[17:0] Result_acc_184_nl;
  wire[18:0] nl_Result_acc_184_nl;
  wire[18:0] MultLoop_acc_114_nl;
  wire[19:0] nl_MultLoop_acc_114_nl;
  wire[22:0] Result_acc_nl;
  wire[23:0] nl_Result_acc_nl;
  wire[17:0] Result_acc_170_nl;
  wire[18:0] nl_Result_acc_170_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl;
  wire[17:0] MultLoop_acc_360_nl;
  wire[18:0] nl_MultLoop_acc_360_nl;
  wire[19:0] MultLoop_acc_169_nl;
  wire[20:0] nl_MultLoop_acc_169_nl;
  wire[9:0] MultLoop_acc_359_nl;
  wire[10:0] nl_MultLoop_acc_359_nl;
  wire[17:0] MultLoop_acc_362_nl;
  wire[18:0] nl_MultLoop_acc_362_nl;
  wire[23:0] MultLoop_acc_172_nl;
  wire[24:0] nl_MultLoop_acc_172_nl;
  wire[20:0] MultLoop_acc_171_nl;
  wire[21:0] nl_MultLoop_acc_171_nl;
  wire[11:0] MultLoop_acc_361_nl;
  wire[12:0] nl_MultLoop_acc_361_nl;
  wire[24:0] MultLoop_acc_113_nl;
  wire[25:0] nl_MultLoop_acc_113_nl;
  wire[20:0] MultLoop_acc_175_nl;
  wire[21:0] nl_MultLoop_acc_175_nl;
  wire[22:0] MultLoop_acc_78_nl;
  wire[23:0] nl_MultLoop_acc_78_nl;
  wire[20:0] MultLoop_acc_167_nl;
  wire[21:0] nl_MultLoop_acc_167_nl;
  wire[13:0] MultLoop_acc_364_nl;
  wire[14:0] nl_MultLoop_acc_364_nl;
  wire[22:0] MultLoop_acc_84_nl;
  wire[23:0] nl_MultLoop_acc_84_nl;
  wire[20:0] MultLoop_acc_165_nl;
  wire[21:0] nl_MultLoop_acc_165_nl;
  wire[17:0] MultLoop_acc_86_nl;
  wire[18:0] nl_MultLoop_acc_86_nl;
  wire[9:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl;
  wire[10:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl;
  wire[19:0] MultLoop_acc_80_nl;
  wire[20:0] nl_MultLoop_acc_80_nl;
  wire[23:0] Result_acc_23_nl;
  wire[24:0] nl_Result_acc_23_nl;
  wire[20:0] Result_acc_187_nl;
  wire[22:0] nl_Result_acc_187_nl;
  wire[25:0] Result_acc_11_nl;
  wire[26:0] nl_Result_acc_11_nl;
  wire[11:0] Result_acc_201_nl;
  wire[12:0] nl_Result_acc_201_nl;
  wire[19:0] Result_acc_202_nl;
  wire[20:0] nl_Result_acc_202_nl;
  wire[25:0] Result_acc_190_nl;
  wire[27:0] nl_Result_acc_190_nl;
  wire[20:0] Result_acc_24_nl;
  wire[21:0] nl_Result_acc_24_nl;
  wire[17:0] Result_acc_192_nl;
  wire[18:0] nl_Result_acc_192_nl;
  wire[13:0] Result_acc_203_nl;
  wire[14:0] nl_Result_acc_203_nl;
  wire[17:0] MultLoop_acc_238_nl;
  wire[20:0] nl_MultLoop_acc_238_nl;
  wire[25:0] MultLoop_acc_65_nl;
  wire[26:0] nl_MultLoop_acc_65_nl;
  wire[23:0] MultLoop_acc_192_nl;
  wire[25:0] nl_MultLoop_acc_192_nl;
  wire[18:0] MultLoop_acc_393_nl;
  wire[19:0] nl_MultLoop_acc_393_nl;
  wire[24:0] MultLoop_acc_68_nl;
  wire[26:0] nl_MultLoop_acc_68_nl;
  wire[12:0] MultLoop_acc_346_nl;
  wire[13:0] nl_MultLoop_acc_346_nl;
  wire[17:0] MultLoop_acc_348_nl;
  wire[18:0] nl_MultLoop_acc_348_nl;
  wire[21:0] MultLoop_acc_188_nl;
  wire[22:0] nl_MultLoop_acc_188_nl;
  wire[11:0] MultLoop_acc_347_nl;
  wire[12:0] nl_MultLoop_acc_347_nl;
  wire[24:0] MultLoop_acc_66_nl;
  wire[25:0] nl_MultLoop_acc_66_nl;
  wire[22:0] MultLoop_acc_190_nl;
  wire[23:0] nl_MultLoop_acc_190_nl;
  wire[20:0] MultLoop_acc_189_nl;
  wire[21:0] nl_MultLoop_acc_189_nl;
  wire[21:0] MultLoop_acc_108_nl;
  wire[22:0] nl_MultLoop_acc_108_nl;
  wire[17:0] MultLoop_acc_195_nl;
  wire[18:0] nl_MultLoop_acc_195_nl;
  wire[12:0] MultLoop_acc_349_nl;
  wire[13:0] nl_MultLoop_acc_349_nl;
  wire[24:0] MultLoop_acc_77_nl;
  wire[26:0] nl_MultLoop_acc_77_nl;
  wire[17:0] MultLoop_acc_236_nl;
  wire[19:0] nl_MultLoop_acc_236_nl;
  wire[23:0] MultLoop_acc_110_nl;
  wire[24:0] nl_MultLoop_acc_110_nl;
  wire[17:0] MultLoop_acc_206_nl;
  wire[18:0] nl_MultLoop_acc_206_nl;
  wire[11:0] MultLoop_acc_356_nl;
  wire[12:0] nl_MultLoop_acc_356_nl;
  wire[23:0] MultLoop_acc_109_nl;
  wire[24:0] nl_MultLoop_acc_109_nl;
  wire[22:0] MultLoop_acc_208_nl;
  wire[23:0] nl_MultLoop_acc_208_nl;
  wire[17:0] MultLoop_acc_207_nl;
  wire[18:0] nl_MultLoop_acc_207_nl;
  wire[17:0] MultLoop_acc_358_nl;
  wire[18:0] nl_MultLoop_acc_358_nl;
  wire[23:0] MultLoop_acc_212_nl;
  wire[25:0] nl_MultLoop_acc_212_nl;
  wire[9:0] MultLoop_acc_357_nl;
  wire[10:0] nl_MultLoop_acc_357_nl;
  wire[26:0] MultLoop_acc_57_nl;
  wire[27:0] nl_MultLoop_acc_57_nl;
  wire[24:0] MultLoop_acc_214_nl;
  wire[26:0] nl_MultLoop_acc_214_nl;
  wire[17:0] MultLoop_acc_235_nl;
  wire[18:0] nl_MultLoop_acc_235_nl;
  wire[17:0] MultLoop_acc_227_nl;
  wire[18:0] nl_MultLoop_acc_227_nl;
  wire[14:0] MultLoop_acc_53_nl;
  wire[15:0] nl_MultLoop_acc_53_nl;
  wire[18:0] MultLoop_acc_343_nl;
  wire[19:0] nl_MultLoop_acc_343_nl;
  wire[24:0] MultLoop_acc_217_nl;
  wire[25:0] nl_MultLoop_acc_217_nl;
  wire[22:0] MultLoop_acc_216_nl;
  wire[23:0] nl_MultLoop_acc_216_nl;
  wire[20:0] MultLoop_acc_215_nl;
  wire[21:0] nl_MultLoop_acc_215_nl;
  wire[17:0] MultLoop_acc_234_nl;
  wire[20:0] nl_MultLoop_acc_234_nl;
  wire[27:0] MultLoop_acc_64_nl;
  wire[29:0] nl_MultLoop_acc_64_nl;
  wire[9:0] MultLoop_acc_344_nl;
  wire[10:0] nl_MultLoop_acc_344_nl;
  wire[22:0] MultLoop_acc_58_nl;
  wire[23:0] nl_MultLoop_acc_58_nl;
  wire[21:0] MultLoop_acc_182_nl;
  wire[22:0] nl_MultLoop_acc_182_nl;
  wire[21:0] MultLoop_acc_107_nl;
  wire[22:0] nl_MultLoop_acc_107_nl;
  wire[20:0] MultLoop_acc_184_nl;
  wire[21:0] nl_MultLoop_acc_184_nl;
  wire[17:0] MultLoop_acc_183_nl;
  wire[18:0] nl_MultLoop_acc_183_nl;
  wire[22:0] MultLoop_acc_73_nl;
  wire[23:0] nl_MultLoop_acc_73_nl;
  wire[19:0] MultLoop_acc_177_nl;
  wire[20:0] nl_MultLoop_acc_177_nl;
  wire[13:0] MultLoop_acc_345_nl;
  wire[14:0] nl_MultLoop_acc_345_nl;
  wire[17:0] MultLoop_acc_353_nl;
  wire[18:0] nl_MultLoop_acc_353_nl;
  wire[18:0] MultLoop_acc_352_nl;
  wire[19:0] nl_MultLoop_acc_352_nl;
  wire[23:0] MultLoop_acc_198_nl;
  wire[24:0] nl_MultLoop_acc_198_nl;
  wire[20:0] MultLoop_acc_197_nl;
  wire[21:0] nl_MultLoop_acc_197_nl;
  wire[9:0] MultLoop_acc_351_nl;
  wire[10:0] nl_MultLoop_acc_351_nl;
  wire[17:0] MultLoop_acc_355_nl;
  wire[18:0] nl_MultLoop_acc_355_nl;
  wire[22:0] MultLoop_acc_202_nl;
  wire[23:0] nl_MultLoop_acc_202_nl;
  wire[19:0] MultLoop_acc_201_nl;
  wire[20:0] nl_MultLoop_acc_201_nl;
  wire[11:0] MultLoop_acc_354_nl;
  wire[12:0] nl_MultLoop_acc_354_nl;
  wire[22:0] MultLoop_acc_111_nl;
  wire[23:0] nl_MultLoop_acc_111_nl;
  wire[19:0] MultLoop_acc_204_nl;
  wire[20:0] nl_MultLoop_acc_204_nl;
  wire[17:0] MultLoop_acc_203_nl;
  wire[18:0] nl_MultLoop_acc_203_nl;
  wire[18:0] MultLoop_acc_112_nl;
  wire[19:0] nl_MultLoop_acc_112_nl;
  wire[10:0] MultLoop_acc_363_nl;
  wire[11:0] nl_MultLoop_acc_363_nl;
  wire[22:0] MultLoop_acc_106_nl;
  wire[23:0] nl_MultLoop_acc_106_nl;
  wire[17:0] MultLoop_acc_118_nl;
  wire[18:0] nl_MultLoop_acc_118_nl;
  wire[17:0] Result_acc_43_nl;
  wire[18:0] nl_Result_acc_43_nl;
  wire[23:0] MultLoop_acc_72_nl;
  wire[24:0] nl_MultLoop_acc_72_nl;
  wire[19:0] MultLoop_acc_181_nl;
  wire[20:0] nl_MultLoop_acc_181_nl;
  wire[21:0] MultLoop_acc_54_nl;
  wire[22:0] nl_MultLoop_acc_54_nl;
  wire[20:0] MultLoop_acc_117_nl;
  wire[21:0] nl_MultLoop_acc_117_nl;
  wire[17:0] MultLoop_acc_116_nl;
  wire[18:0] nl_MultLoop_acc_116_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [107:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_107_90 , res_rsci_d_89_72 , res_rsci_d_71_54
      , res_rsci_d_53_36 , res_rsci_d_35_18 , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd432)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd108)) res_rsci (
      .d(nl_res_rsci_d[107:0]),
      .z(res_rsc_z)
    );
  assign nl_MultLoop_acc_363_nl = conv_s2s_10_11(data_rsci_idat[71:62]) + 11'b00000000001;
  assign MultLoop_acc_363_nl = nl_MultLoop_acc_363_nl[10:0];
  assign nl_MultLoop_acc_174_cse_1 = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({(MultLoop_acc_363_nl)
      , (data_rsci_idat[61:56])});
  assign MultLoop_acc_174_cse_1 = nl_MultLoop_acc_174_cse_1[17:0];
  assign nl_Result_acc_137_cse_1 = (~ (data_rsci_idat[89:72])) + conv_s2s_15_18(data_rsci_idat[89:75]);
  assign Result_acc_137_cse_1 = nl_Result_acc_137_cse_1[17:0];
  assign nl_MultLoop_acc_118_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18(data_rsci_idat[35:20]);
  assign MultLoop_acc_118_nl = nl_MultLoop_acc_118_nl[17:0];
  assign nl_MultLoop_acc_106_nl = conv_s2u_18_23(MultLoop_acc_118_nl) + ({(data_rsci_idat[35:18])
      , 5'b00001});
  assign MultLoop_acc_106_nl = nl_MultLoop_acc_106_nl[22:0];
  assign MultLoop_acc_106_itm_22_6 = readslicef_23_17_6((MultLoop_acc_106_nl));
  assign nl_Result_acc_131_cse_1 = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_15_19(data_rsci_idat[161:147]);
  assign Result_acc_131_cse_1 = nl_Result_acc_131_cse_1[18:0];
  assign nl_Result_acc_43_nl = conv_s2u_13_18(data_rsci_idat[377:365]) - (data_rsci_idat[377:360]);
  assign Result_acc_43_nl = nl_Result_acc_43_nl[17:0];
  assign Result_acc_43_itm_17_5 = readslicef_18_13_5((Result_acc_43_nl));
  assign nl_Result_acc_172_cse_1 = conv_s2s_18_19(data_rsci_idat[215:198]) + conv_s2s_16_19(data_rsci_idat[215:200]);
  assign Result_acc_172_cse_1 = nl_Result_acc_172_cse_1[18:0];
  assign nl_MultLoop_acc_263_cse_1 = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[251:234]));
  assign MultLoop_acc_263_cse_1 = nl_MultLoop_acc_263_cse_1[19:0];
  assign nl_MultLoop_acc_76_cse_1 = conv_s2s_18_20(~ (data_rsci_idat[413:396])) +
      ({(data_rsci_idat[413:396]) , 2'b01});
  assign MultLoop_acc_76_cse_1 = nl_MultLoop_acc_76_cse_1[19:0];
  assign nl_MultLoop_acc_181_nl = ({(data_rsci_idat[341:324]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[341:324]));
  assign MultLoop_acc_181_nl = nl_MultLoop_acc_181_nl[19:0];
  assign nl_MultLoop_acc_72_nl = conv_s2s_20_24(MultLoop_acc_181_nl) + conv_s2s_23_24({(data_rsci_idat[341:324])
      , 5'b00000});
  assign MultLoop_acc_72_nl = nl_MultLoop_acc_72_nl[23:0];
  assign MultLoop_acc_72_itm_23_7 = readslicef_24_17_7((MultLoop_acc_72_nl));
  assign nl_MultLoop_acc_193_cse_1 = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_193_cse_1 = nl_MultLoop_acc_193_cse_1[19:0];
  assign nl_MultLoop_acc_116_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_15_18(data_rsci_idat[17:3]);
  assign MultLoop_acc_116_nl = nl_MultLoop_acc_116_nl[17:0];
  assign nl_MultLoop_acc_117_nl = conv_s2s_20_21({(~ (data_rsci_idat[17:0])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_116_nl);
  assign MultLoop_acc_117_nl = nl_MultLoop_acc_117_nl[20:0];
  assign nl_MultLoop_acc_54_nl = conv_s2u_21_22(MultLoop_acc_117_nl) + ({(data_rsci_idat[17:0])
      , 4'b0100});
  assign MultLoop_acc_54_nl = nl_MultLoop_acc_54_nl[21:0];
  assign MultLoop_acc_54_itm_21_5 = readslicef_22_17_5((MultLoop_acc_54_nl));
  assign nl_MultLoop_MultLoop_conc_50_18_6 =  -conv_s2s_12_13(data_rsci_idat[431:420]);
  assign MultLoop_MultLoop_conc_50_18_6 = nl_MultLoop_MultLoop_conc_50_18_6[12:0];
  assign nl_MultLoop_acc_395 = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[305:288]));
  assign MultLoop_acc_395 = nl_MultLoop_acc_395[19:0];
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_107_90 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_89_72 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
      res_rsci_d_71_54 <= 18'b000000000000000000;
      res_rsci_d_53_36 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_107_90 <= nl_res_rsci_d_107_90[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_89_72 <= nl_res_rsci_d_89_72[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
      res_rsci_d_71_54 <= nl_res_rsci_d_71_54[17:0];
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
    end
  end
  assign nl_Result_acc_110_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_174_cse_1);
  assign Result_acc_110_nl = nl_Result_acc_110_nl[19:0];
  assign nl_Result_acc_111_nl = ({(~ (data_rsci_idat[71:54])) , 4'b0000}) + conv_s2s_20_22(Result_acc_110_nl);
  assign Result_acc_111_nl = nl_Result_acc_111_nl[21:0];
  assign nl_Result_acc_84_nl = conv_s2u_22_25(Result_acc_111_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[71:54])) , 6'b010000});
  assign Result_acc_84_nl = nl_Result_acc_84_nl[24:0];
  assign nl_Result_acc_113_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[107:90])) , 4'b0001}) + conv_s2s_18_25(~
      (data_rsci_idat[107:90]));
  assign Result_acc_113_nl = nl_Result_acc_113_nl[24:0];
  assign nl_Result_acc_62_nl = conv_s2s_25_27(Result_acc_113_nl) + ({(data_rsci_idat[107:90])
      , 9'b001000000});
  assign Result_acc_62_nl = nl_Result_acc_62_nl[26:0];
  assign nl_Result_acc_100_nl = (~ (data_rsci_idat[215:198])) + conv_s2s_16_18(data_rsci_idat[215:200]);
  assign Result_acc_100_nl = nl_Result_acc_100_nl[17:0];
  assign nl_Result_acc_83_nl = conv_s2u_18_22(Result_acc_100_nl) + ({(data_rsci_idat[215:198])
      , 4'b0001});
  assign Result_acc_83_nl = nl_Result_acc_83_nl[21:0];
  assign nl_Result_acc_217_nl =  -conv_s2s_10_11(data_rsci_idat[305:296]);
  assign Result_acc_217_nl = nl_Result_acc_217_nl[10:0];
  assign nl_Result_acc_103_nl = ({(data_rsci_idat[305:288]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[305:288])) , 4'b0001}) + conv_s2s_19_24({(Result_acc_217_nl)
      , (~ (data_rsci_idat[295:288]))});
  assign Result_acc_103_nl = nl_Result_acc_103_nl[23:0];
  assign nl_Result_acc_218_nl = conv_s2u_16_18(readslicef_24_16_8((Result_acc_103_nl)))
      + (~ (data_rsci_idat[305:288]));
  assign Result_acc_218_nl = nl_Result_acc_218_nl[17:0];
  assign nl_Result_acc_219_nl = conv_s2s_10_11(data_rsci_idat[431:422]) + 11'b00000000001;
  assign Result_acc_219_nl = nl_Result_acc_219_nl[10:0];
  assign nl_Result_acc_107_nl = conv_s2s_22_23({(data_rsci_idat[431:414]) , 4'b0000})
      + conv_s2s_20_23({(data_rsci_idat[431:414]) , 2'b00}) + conv_s2s_18_23(data_rsci_idat[431:414])
      + conv_s2s_17_23({(Result_acc_219_nl) , (data_rsci_idat[421:416])});
  assign Result_acc_107_nl = nl_Result_acc_107_nl[22:0];
  assign nl_Result_acc_220_nl = conv_s2u_17_18(readslicef_23_17_6((Result_acc_107_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign Result_acc_220_nl = nl_Result_acc_220_nl[17:0];
  assign nl_Result_acc_88_nl = conv_s2s_21_22({(~ (data_rsci_idat[17:0])) , 3'b001})
      + conv_s2s_18_22(~ (data_rsci_idat[17:0]));
  assign Result_acc_88_nl = nl_Result_acc_88_nl[21:0];
  assign nl_Result_acc_57_nl = conv_s2s_22_24(Result_acc_88_nl) + ({(data_rsci_idat[17:0])
      , 6'b001000});
  assign Result_acc_57_nl = nl_Result_acc_57_nl[23:0];
  assign nl_Result_acc_221_nl = conv_s2s_12_13(data_rsci_idat[53:42]) + 13'b0000000000001;
  assign Result_acc_221_nl = nl_Result_acc_221_nl[12:0];
  assign nl_Result_acc_90_nl = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_16_19({(Result_acc_221_nl)
      , (data_rsci_idat[41:39])});
  assign Result_acc_90_nl = nl_Result_acc_90_nl[18:0];
  assign nl_Result_acc_59_nl = conv_s2u_19_21(Result_acc_90_nl) + ({(~ (data_rsci_idat[53:36]))
      , 3'b000});
  assign Result_acc_59_nl = nl_Result_acc_59_nl[20:0];
  assign nl_MultLoop_acc_139_nl = conv_s2s_17_18(readslicef_25_17_8((Result_acc_84_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((Result_acc_62_nl))) + conv_s2s_16_18(readslicef_22_16_6((Result_acc_83_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((Result_acc_218_nl))) + conv_s2s_16_18(readslicef_18_16_2((Result_acc_220_nl)))
      + conv_s2s_14_18(readslicef_24_14_10((Result_acc_57_nl))) + conv_s2s_14_18(readslicef_21_14_7((Result_acc_59_nl)));
  assign MultLoop_acc_139_nl = nl_MultLoop_acc_139_nl[17:0];
  assign nl_Result_acc_223_nl =  -conv_s2s_11_12(data_rsci_idat[125:115]);
  assign Result_acc_223_nl = nl_Result_acc_223_nl[11:0];
  assign nl_Result_acc_63_nl = conv_s2s_25_26({(~ (data_rsci_idat[125:108])) , 7'b0100000})
      + conv_s2s_23_26({(~ (data_rsci_idat[125:108])) , 5'b00001}) + conv_s2s_19_26({(Result_acc_223_nl)
      , (~ (data_rsci_idat[114:108]))});
  assign Result_acc_63_nl = nl_Result_acc_63_nl[25:0];
  assign nl_Result_acc_224_nl = conv_s2s_11_12(data_rsci_idat[233:223]) + 12'b000000000001;
  assign Result_acc_224_nl = nl_Result_acc_224_nl[11:0];
  assign nl_Result_acc_117_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_16_18({(Result_acc_224_nl)
      , (data_rsci_idat[222:219])});
  assign Result_acc_117_nl = nl_Result_acc_117_nl[17:0];
  assign nl_Result_acc_85_nl = conv_s2u_18_23(Result_acc_117_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[233:216])) , 4'b0001});
  assign Result_acc_85_nl = nl_Result_acc_85_nl[22:0];
  assign nl_Result_acc_225_nl =  -conv_s2s_9_10(data_rsci_idat[251:243]);
  assign Result_acc_225_nl = nl_Result_acc_225_nl[9:0];
  assign nl_Result_acc_119_nl = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_19_20({(Result_acc_225_nl)
      , (~ (data_rsci_idat[242:234]))});
  assign Result_acc_119_nl = nl_Result_acc_119_nl[19:0];
  assign nl_Result_acc_121_nl = conv_s2s_24_25({(data_rsci_idat[251:234]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[251:234]) , 4'b0000}) + conv_s2s_20_25(Result_acc_119_nl);
  assign Result_acc_121_nl = nl_Result_acc_121_nl[24:0];
  assign nl_Result_acc_226_nl = conv_s2u_16_18(readslicef_25_16_9((Result_acc_121_nl)))
      + (~ (data_rsci_idat[251:234]));
  assign Result_acc_226_nl = nl_Result_acc_226_nl[17:0];
  assign nl_Result_acc_227_nl =  -conv_s2s_10_11(data_rsci_idat[269:260]);
  assign Result_acc_227_nl = nl_Result_acc_227_nl[10:0];
  assign nl_Result_acc_123_nl = ({(data_rsci_idat[269:252]) , 3'b001}) + conv_s2s_19_21({(Result_acc_227_nl)
      , (~ (data_rsci_idat[259:252]))});
  assign Result_acc_123_nl = nl_Result_acc_123_nl[20:0];
  assign nl_Result_acc_228_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_15_18(readslicef_21_15_6((Result_acc_123_nl)));
  assign Result_acc_228_nl = nl_Result_acc_228_nl[17:0];
  assign nl_Result_acc_229_nl = conv_s2u_18_21(Result_acc_228_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[269:252])) , 2'b01});
  assign Result_acc_229_nl = nl_Result_acc_229_nl[20:0];
  assign nl_MultLoop_acc_138_nl = conv_s2s_17_18(readslicef_26_17_9((Result_acc_63_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((Result_acc_85_nl))) + conv_s2s_17_18(readslicef_18_17_1((Result_acc_226_nl)))
      + conv_s2s_17_18(readslicef_21_17_4((Result_acc_229_nl)));
  assign MultLoop_acc_138_nl = nl_MultLoop_acc_138_nl[17:0];
  assign nl_Result_acc_96_nl = conv_s2s_20_21({(data_rsci_idat[161:144]) , 2'b00})
      + conv_s2s_19_21(Result_acc_131_cse_1);
  assign Result_acc_96_nl = nl_Result_acc_96_nl[20:0];
  assign nl_Result_acc_82_nl = conv_s2u_21_23(Result_acc_96_nl) + conv_s2u_22_23({(data_rsci_idat[161:144])
      , 4'b0000});
  assign Result_acc_82_nl = nl_Result_acc_82_nl[22:0];
  assign nl_Result_acc_232_nl =  -conv_s2s_12_13(data_rsci_idat[197:186]);
  assign Result_acc_232_nl = nl_Result_acc_232_nl[12:0];
  assign nl_Result_acc_65_nl = conv_s2s_24_25({(~ (data_rsci_idat[197:180])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[197:180])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[197:180])) , 2'b01}) + conv_s2s_19_25({(Result_acc_232_nl)
      , (~ (data_rsci_idat[185:180]))});
  assign Result_acc_65_nl = nl_Result_acc_65_nl[24:0];
  assign nl_Result_acc_125_nl = ({(data_rsci_idat[287:270]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[287:270]));
  assign Result_acc_125_nl = nl_Result_acc_125_nl[21:0];
  assign nl_Result_acc_230_nl = conv_s2u_15_19(readslicef_22_15_7((Result_acc_125_nl)))
      + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign Result_acc_230_nl = nl_Result_acc_230_nl[18:0];
  assign nl_Result_acc_127_nl = conv_s2s_24_25({(~ (data_rsci_idat[359:342])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[359:342])) , 4'b0001}) + conv_s2s_18_25(~
      (data_rsci_idat[359:342]));
  assign Result_acc_127_nl = nl_Result_acc_127_nl[24:0];
  assign nl_Result_acc_74_nl = conv_s2s_25_27(Result_acc_127_nl) + ({(data_rsci_idat[359:342])
      , 9'b001000000});
  assign Result_acc_74_nl = nl_Result_acc_74_nl[26:0];
  assign nl_Result_acc_130_nl = ({(~ (data_rsci_idat[377:360])) , 4'b0000}) + conv_s2s_20_22({(data_rsci_idat[377:360])
      , 2'b00}) + conv_s2s_18_22(data_rsci_idat[377:360]) + conv_s2s_15_22(data_rsci_idat[377:363]);
  assign Result_acc_130_nl = nl_Result_acc_130_nl[21:0];
  assign nl_Result_acc_86_nl = conv_s2u_22_24(Result_acc_130_nl) + ({(data_rsci_idat[377:360])
      , 6'b010000});
  assign Result_acc_86_nl = nl_Result_acc_86_nl[23:0];
  assign nl_Result_acc_73_nl = conv_s2u_12_18(data_rsci_idat[341:330]) - (data_rsci_idat[341:324]);
  assign Result_acc_73_nl = nl_Result_acc_73_nl[17:0];
  assign nl_Result_acc_91_nl = conv_s2s_20_21({(~ (data_rsci_idat[323:306])) , 2'b01})
      + conv_s2s_18_21(~ (data_rsci_idat[323:306]));
  assign Result_acc_91_nl = nl_Result_acc_91_nl[20:0];
  assign nl_Result_acc_72_nl = conv_s2s_21_24(Result_acc_91_nl) + ({(data_rsci_idat[323:306])
      , 6'b000100});
  assign Result_acc_72_nl = nl_Result_acc_72_nl[23:0];
  assign nl_Result_acc_231_nl = conv_s2s_12_13(data_rsci_idat[395:384]) + 13'b0000000000001;
  assign Result_acc_231_nl = nl_Result_acc_231_nl[12:0];
  assign nl_Result_acc_93_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_17_18({(Result_acc_231_nl)
      , (data_rsci_idat[383:380])});
  assign Result_acc_93_nl = nl_Result_acc_93_nl[17:0];
  assign nl_Result_acc_94_nl = conv_s2s_20_21({(~ (data_rsci_idat[395:378])) , 2'b01})
      + conv_s2s_18_21(Result_acc_93_nl);
  assign Result_acc_94_nl = nl_Result_acc_94_nl[20:0];
  assign nl_Result_acc_80_nl = conv_s2u_21_23(Result_acc_94_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[395:378])) , 4'b0100});
  assign Result_acc_80_nl = nl_Result_acc_80_nl[22:0];
  assign nl_Result_acc_79_nl = conv_s2u_18_20(Result_acc_137_cse_1) + ({(data_rsci_idat[89:72])
      , 2'b01});
  assign Result_acc_79_nl = nl_Result_acc_79_nl[19:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl = ~((data_rsci_idat[168:162]!=7'b0000000));
  assign nl_MultLoop_acc_119_nl = conv_u2s_6_12({5'b10100 , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl)})
      - conv_s2s_11_12(data_rsci_idat[179:169]);
  assign MultLoop_acc_119_nl = nl_MultLoop_acc_119_nl[11:0];
  assign nl_Result_acc_77_nl = conv_s2u_14_18(data_rsci_idat[413:400]) - (data_rsci_idat[413:396]);
  assign Result_acc_77_nl = nl_Result_acc_77_nl[17:0];
  assign nl_res_rsci_d_107_90  = (MultLoop_acc_139_nl) + (MultLoop_acc_138_nl) +
      conv_s2s_16_18(MultLoop_acc_106_itm_22_6[16:1]) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_82_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((Result_acc_65_nl))) + conv_s2s_17_18(readslicef_19_17_2((Result_acc_230_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((Result_acc_74_nl))) + conv_s2s_17_18(readslicef_24_17_7((Result_acc_86_nl)))
      + conv_s2s_15_18(readslicef_18_15_3((Result_acc_73_nl))) + conv_s2s_14_18(data_rsci_idat[143:130])
      + conv_s2s_14_18(readslicef_24_14_10((Result_acc_72_nl))) + conv_s2s_15_18(readslicef_23_15_8((Result_acc_80_nl)))
      + conv_s2s_13_18(readslicef_20_13_7((Result_acc_79_nl))) + conv_s2s_12_18(MultLoop_acc_119_nl)
      + conv_s2s_12_18(readslicef_18_12_6((Result_acc_77_nl)));
  assign nl_MultLoop_acc_292_nl = ({(~ (data_rsci_idat[395:378])) , 5'b00000}) +
      conv_s2s_21_23({(data_rsci_idat[395:378]) , 3'b000}) + conv_s2s_18_23(data_rsci_idat[395:378])
      + conv_s2s_16_23(data_rsci_idat[395:380]);
  assign MultLoop_acc_292_nl = nl_MultLoop_acc_292_nl[22:0];
  assign nl_MultLoop_acc_97_nl = conv_s2u_23_25(MultLoop_acc_292_nl) + ({(data_rsci_idat[395:378])
      , 7'b0100000});
  assign MultLoop_acc_97_nl = nl_MultLoop_acc_97_nl[24:0];
  assign nl_MultLoop_acc_289_nl = conv_s2s_20_21({(data_rsci_idat[89:72]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[89:72]) + conv_s2s_16_21(data_rsci_idat[89:74]);
  assign MultLoop_acc_289_nl = nl_MultLoop_acc_289_nl[20:0];
  assign nl_MultLoop_acc_90_nl = conv_s2u_21_23(MultLoop_acc_289_nl) + conv_s2u_22_23({(data_rsci_idat[89:72])
      , 4'b0000});
  assign MultLoop_acc_90_nl = nl_MultLoop_acc_90_nl[22:0];
  assign nl_MultLoop_acc_375_nl = conv_s2s_10_11(data_rsci_idat[413:404]) + 11'b00000000001;
  assign MultLoop_acc_375_nl = nl_MultLoop_acc_375_nl[10:0];
  assign nl_MultLoop_acc_286_nl = conv_s2s_21_22({(data_rsci_idat[413:396]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[413:396]) + conv_s2s_16_22({(MultLoop_acc_375_nl)
      , (data_rsci_idat[403:399])});
  assign MultLoop_acc_286_nl = nl_MultLoop_acc_286_nl[21:0];
  assign nl_MultLoop_acc_28_nl = conv_s2u_22_23(MultLoop_acc_286_nl) + ({(~ (data_rsci_idat[413:396]))
      , 5'b00000});
  assign MultLoop_acc_28_nl = nl_MultLoop_acc_28_nl[22:0];
  assign nl_MultLoop_acc_396_nl = conv_s2u_14_19(MultLoop_acc_395[19:6]) + conv_s2u_18_19(data_rsci_idat[305:288]);
  assign MultLoop_acc_396_nl = nl_MultLoop_acc_396_nl[18:0];
  assign nl_MultLoop_acc_283_nl = conv_s2s_20_21({(~ (data_rsci_idat[161:144])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_283_nl = nl_MultLoop_acc_283_nl[20:0];
  assign nl_MultLoop_acc_14_nl = conv_s2s_21_24(MultLoop_acc_283_nl) + ({(data_rsci_idat[161:144])
      , 6'b000100});
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[23:0];
  assign nl_MultLoop_acc_96_nl = conv_s2u_13_19(data_rsci_idat[377:365]) + conv_s2u_18_19(data_rsci_idat[377:360]);
  assign MultLoop_acc_96_nl = nl_MultLoop_acc_96_nl[18:0];
  assign nl_MultLoop_acc_287_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_287_nl = nl_MultLoop_acc_287_nl[19:0];
  assign nl_MultLoop_acc_376_nl = conv_s2u_13_19(readslicef_20_13_7((MultLoop_acc_287_nl)))
      + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_376_nl = nl_MultLoop_acc_376_nl[18:0];
  assign nl_MultLoop_acc_279_nl = ({(data_rsci_idat[431:414]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_50_18_6
      , (~ (data_rsci_idat[419:414]))});
  assign MultLoop_acc_279_nl = nl_MultLoop_acc_279_nl[19:0];
  assign nl_MultLoop_acc_378_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_279_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_378_nl = nl_MultLoop_acc_378_nl[17:0];
  assign nl_MultLoop_acc_379_nl = conv_s2s_13_14(data_rsci_idat[71:59]) + 14'b00000000000001;
  assign MultLoop_acc_379_nl = nl_MultLoop_acc_379_nl[13:0];
  assign nl_MultLoop_acc_277_nl = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_17_19({(MultLoop_acc_379_nl)
      , (data_rsci_idat[58:56])});
  assign MultLoop_acc_277_nl = nl_MultLoop_acc_277_nl[18:0];
  assign nl_MultLoop_acc_9_nl = conv_s2u_19_21(MultLoop_acc_277_nl) + ({(~ (data_rsci_idat[71:54]))
      , 3'b000});
  assign MultLoop_acc_9_nl = nl_MultLoop_acc_9_nl[20:0];
  assign nl_MultLoop_acc_340_nl = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_97_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_90_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_28_nl)))
      + conv_s2s_15_18(readslicef_19_15_4((MultLoop_acc_396_nl))) + conv_s2s_15_18(readslicef_24_15_9((MultLoop_acc_14_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_96_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_376_nl)))
      + conv_s2s_14_18(readslicef_18_14_4((MultLoop_acc_378_nl))) + conv_s2s_13_18(readslicef_21_13_8((MultLoop_acc_9_nl)));
  assign MultLoop_acc_340_nl = nl_MultLoop_acc_340_nl[17:0];
  assign nl_MultLoop_acc_293_nl = ({(data_rsci_idat[359:342]) , 5'b00001}) + conv_s2s_18_23(~
      (data_rsci_idat[359:342]));
  assign MultLoop_acc_293_nl = nl_MultLoop_acc_293_nl[22:0];
  assign nl_MultLoop_acc_380_nl = conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_293_nl)))
      + conv_s2u_18_19(data_rsci_idat[359:342]);
  assign MultLoop_acc_380_nl = nl_MultLoop_acc_380_nl[18:0];
  assign nl_MultLoop_acc_295_nl = conv_s2s_25_26({(~ (data_rsci_idat[341:324])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[341:324])) , 5'b00001}) +
      conv_s2s_18_26(~ (data_rsci_idat[341:324]));
  assign MultLoop_acc_295_nl = nl_MultLoop_acc_295_nl[25:0];
  assign nl_MultLoop_acc_381_nl = conv_s2u_19_20(readslicef_26_19_7((MultLoop_acc_295_nl)))
      + ({(data_rsci_idat[341:324]) , 2'b01});
  assign MultLoop_acc_381_nl = nl_MultLoop_acc_381_nl[19:0];
  assign nl_MultLoop_acc_296_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_16_18(data_rsci_idat[251:236]);
  assign MultLoop_acc_296_nl = nl_MultLoop_acc_296_nl[17:0];
  assign nl_MultLoop_acc_297_nl = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_296_nl);
  assign MultLoop_acc_297_nl = nl_MultLoop_acc_297_nl[19:0];
  assign nl_MultLoop_acc_298_nl = conv_s2s_22_23({(data_rsci_idat[251:234]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_297_nl);
  assign MultLoop_acc_298_nl = nl_MultLoop_acc_298_nl[22:0];
  assign nl_MultLoop_acc_95_nl = conv_s2u_23_25(MultLoop_acc_298_nl) + conv_s2u_24_25({(data_rsci_idat[251:234])
      , 6'b000000});
  assign MultLoop_acc_95_nl = nl_MultLoop_acc_95_nl[24:0];
  assign nl_MultLoop_acc_382_nl =  -conv_s2s_9_10(data_rsci_idat[269:261]);
  assign MultLoop_acc_382_nl = nl_MultLoop_acc_382_nl[9:0];
  assign nl_MultLoop_acc_300_nl = ({(data_rsci_idat[269:252]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_382_nl)
      , (~ (data_rsci_idat[260:252]))});
  assign MultLoop_acc_300_nl = nl_MultLoop_acc_300_nl[20:0];
  assign nl_MultLoop_acc_301_nl = conv_s2s_23_24({(data_rsci_idat[269:252]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_300_nl);
  assign MultLoop_acc_301_nl = nl_MultLoop_acc_301_nl[23:0];
  assign nl_MultLoop_acc_383_nl = conv_s2u_18_19(data_rsci_idat[269:252]) + conv_s2u_17_19(readslicef_24_17_7((MultLoop_acc_301_nl)));
  assign MultLoop_acc_383_nl = nl_MultLoop_acc_383_nl[18:0];
  assign nl_MultLoop_acc_384_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_383_nl)))
      + (~ (data_rsci_idat[269:252]));
  assign MultLoop_acc_384_nl = nl_MultLoop_acc_384_nl[17:0];
  assign nl_MultLoop_acc_339_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_380_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_381_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_95_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_384_nl)));
  assign MultLoop_acc_339_nl = nl_MultLoop_acc_339_nl[17:0];
  assign nl_MultLoop_acc_314_nl = ({(~ (data_rsci_idat[143:126])) , 4'b0000}) + conv_s2s_18_22(data_rsci_idat[143:126])
      + conv_s2s_16_22(data_rsci_idat[143:128]);
  assign MultLoop_acc_314_nl = nl_MultLoop_acc_314_nl[21:0];
  assign nl_MultLoop_acc_92_nl = conv_s2u_22_24(MultLoop_acc_314_nl) + ({(data_rsci_idat[143:126])
      , 6'b010000});
  assign MultLoop_acc_92_nl = nl_MultLoop_acc_92_nl[23:0];
  assign nl_MultLoop_acc_315_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_16_18(data_rsci_idat[125:110]);
  assign MultLoop_acc_315_nl = nl_MultLoop_acc_315_nl[17:0];
  assign nl_MultLoop_acc_316_nl = conv_s2s_23_24({(~ (data_rsci_idat[125:108])) ,
      5'b00001}) + conv_s2s_18_24(MultLoop_acc_315_nl);
  assign MultLoop_acc_316_nl = nl_MultLoop_acc_316_nl[23:0];
  assign nl_MultLoop_acc_91_nl = conv_s2u_24_25(MultLoop_acc_316_nl) + ({(data_rsci_idat[125:108])
      , 7'b0100000});
  assign MultLoop_acc_91_nl = nl_MultLoop_acc_91_nl[24:0];
  assign nl_MultLoop_acc_390_nl = conv_s2s_11_12(data_rsci_idat[35:25]) + 12'b000000000001;
  assign MultLoop_acc_390_nl = nl_MultLoop_acc_390_nl[11:0];
  assign nl_MultLoop_acc_318_nl = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_14_19({(MultLoop_acc_390_nl)
      , (data_rsci_idat[24:23])});
  assign MultLoop_acc_318_nl = nl_MultLoop_acc_318_nl[18:0];
  assign nl_MultLoop_acc_7_nl = conv_s2u_19_20(MultLoop_acc_318_nl) + ({(~ (data_rsci_idat[35:18]))
      , 2'b00});
  assign MultLoop_acc_7_nl = nl_MultLoop_acc_7_nl[19:0];
  assign nl_MultLoop_acc_89_nl = conv_s2u_15_19(data_rsci_idat[53:39]) + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_89_nl = nl_MultLoop_acc_89_nl[18:0];
  assign nl_MultLoop_acc_322_nl = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_7_nl)))
      + conv_s2s_13_17(readslicef_19_13_6((MultLoop_acc_89_nl))) + 17'b11111111101011011;
  assign MultLoop_acc_322_nl = nl_MultLoop_acc_322_nl[16:0];
  assign nl_MultLoop_acc_391_nl = conv_s2s_12_13(data_rsci_idat[17:6]) + 13'b0000000000001;
  assign MultLoop_acc_391_nl = nl_MultLoop_acc_391_nl[12:0];
  assign nl_MultLoop_acc_320_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_17_18({(MultLoop_acc_391_nl)
      , (data_rsci_idat[5:2])});
  assign MultLoop_acc_320_nl = nl_MultLoop_acc_320_nl[17:0];
  assign nl_MultLoop_acc_6_nl = conv_s2u_18_23(MultLoop_acc_320_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[17:0])) , 4'b0001});
  assign MultLoop_acc_6_nl = nl_MultLoop_acc_6_nl[22:0];
  assign nl_MultLoop_3_MultLoop_acc_3_nl = (MultLoop_acc_322_nl) + (readslicef_23_17_6((MultLoop_acc_6_nl)));
  assign MultLoop_3_MultLoop_acc_3_nl = nl_MultLoop_3_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_23_nl = conv_s2u_16_18(data_rsci_idat[323:308]) - (data_rsci_idat[323:306]);
  assign MultLoop_acc_23_nl = nl_MultLoop_acc_23_nl[17:0];
  assign nl_MultLoop_acc_392_nl =  -conv_s2s_13_14(data_rsci_idat[287:275]);
  assign MultLoop_acc_392_nl = nl_MultLoop_acc_392_nl[13:0];
  assign nl_MultLoop_acc_21_nl = conv_s2s_23_24({(~ (data_rsci_idat[287:270])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[287:270])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_392_nl)
      , (~ (data_rsci_idat[274:270]))});
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[23:0];
  assign nl_MultLoop_acc_337_nl = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_92_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_91_nl))) + conv_s2s_17_18(MultLoop_3_MultLoop_acc_3_nl)
      + conv_s2s_15_18(readslicef_18_15_3((MultLoop_acc_23_nl))) + conv_s2s_15_18(readslicef_24_15_9((MultLoop_acc_21_nl)));
  assign MultLoop_acc_337_nl = nl_MultLoop_acc_337_nl[17:0];
  assign nl_MultLoop_acc_385_nl =  -conv_s2s_12_13(data_rsci_idat[215:204]);
  assign MultLoop_acc_385_nl = nl_MultLoop_acc_385_nl[12:0];
  assign nl_MultLoop_acc_304_nl = ({(data_rsci_idat[215:198]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_385_nl)
      , (~ (data_rsci_idat[203:198]))});
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[19:0];
  assign nl_MultLoop_acc_305_nl = conv_s2s_22_23({(data_rsci_idat[215:198]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_304_nl);
  assign MultLoop_acc_305_nl = nl_MultLoop_acc_305_nl[22:0];
  assign nl_MultLoop_acc_386_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_305_nl)))
      + (~ (data_rsci_idat[215:198]));
  assign MultLoop_acc_386_nl = nl_MultLoop_acc_386_nl[17:0];
  assign nl_MultLoop_acc_387_nl = conv_s2s_10_11(data_rsci_idat[233:224]) + 11'b00000000001;
  assign MultLoop_acc_387_nl = nl_MultLoop_acc_387_nl[10:0];
  assign nl_MultLoop_acc_307_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_16_18({(MultLoop_acc_387_nl)
      , (data_rsci_idat[223:219])});
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[17:0];
  assign nl_MultLoop_acc_94_nl = conv_s2u_18_24(MultLoop_acc_307_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[233:216])) , 5'b00001});
  assign MultLoop_acc_94_nl = nl_MultLoop_acc_94_nl[23:0];
  assign nl_MultLoop_acc_388_nl =  -conv_s2s_10_11(data_rsci_idat[179:170]);
  assign MultLoop_acc_388_nl = nl_MultLoop_acc_388_nl[10:0];
  assign nl_MultLoop_acc_310_nl = ({(data_rsci_idat[179:162]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_388_nl)
      , (~ (data_rsci_idat[169:162]))});
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[22:0];
  assign nl_MultLoop_acc_389_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_310_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_389_nl = nl_MultLoop_acc_389_nl[17:0];
  assign nl_MultLoop_acc_312_nl = ({(~ (data_rsci_idat[197:180])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[197:180])
      + conv_s2s_16_21(data_rsci_idat[197:182]);
  assign MultLoop_acc_312_nl = nl_MultLoop_acc_312_nl[20:0];
  assign nl_MultLoop_acc_93_nl = conv_s2u_21_25(MultLoop_acc_312_nl) + ({(data_rsci_idat[197:180])
      , 7'b0001000});
  assign MultLoop_acc_93_nl = nl_MultLoop_acc_93_nl[24:0];
  assign nl_res_rsci_d_17_0  = (MultLoop_acc_340_nl) + (MultLoop_acc_339_nl) + (MultLoop_acc_337_nl)
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_386_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_94_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_389_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_93_nl)));
  assign nl_Result_acc_169_nl = (~ (data_rsci_idat[413:396])) + conv_s2s_15_18(data_rsci_idat[413:399]);
  assign Result_acc_169_nl = nl_Result_acc_169_nl[17:0];
  assign nl_Result_acc_56_nl = conv_s2u_18_20(Result_acc_169_nl) + ({(data_rsci_idat[413:396])
      , 2'b01});
  assign Result_acc_56_nl = nl_Result_acc_56_nl[19:0];
  assign nl_Result_acc_48_nl = conv_s2u_14_19(data_rsci_idat[143:130]) + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign Result_acc_48_nl = nl_Result_acc_48_nl[18:0];
  assign nl_Result_acc_134_nl = ({(data_rsci_idat[179:162]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[179:162]));
  assign Result_acc_134_nl = nl_Result_acc_134_nl[20:0];
  assign nl_Result_acc_32_nl = conv_s2s_21_25(Result_acc_134_nl) + conv_s2s_24_25({(data_rsci_idat[179:162])
      , 6'b000000});
  assign Result_acc_32_nl = nl_Result_acc_32_nl[24:0];
  assign nl_Result_acc_204_nl =  -conv_s2s_12_13(data_rsci_idat[107:96]);
  assign Result_acc_204_nl = nl_Result_acc_204_nl[12:0];
  assign nl_Result_acc_29_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[107:90])) , 4'b0001}) + conv_s2s_19_25({(Result_acc_204_nl)
      , (~ (data_rsci_idat[95:90]))});
  assign Result_acc_29_nl = nl_Result_acc_29_nl[24:0];
  assign nl_Result_acc_233_nl = conv_s2u_17_19(Result_acc_131_cse_1[18:2]) + conv_s2u_18_19(data_rsci_idat[161:144]);
  assign Result_acc_233_nl = nl_Result_acc_233_nl[18:0];
  assign nl_Result_acc_205_nl = conv_s2s_12_13(data_rsci_idat[359:348]) + 13'b0000000000001;
  assign Result_acc_205_nl = nl_Result_acc_205_nl[12:0];
  assign nl_Result_acc_136_nl = conv_s2s_18_19(data_rsci_idat[359:342]) + conv_s2s_16_19({(Result_acc_205_nl)
      , (data_rsci_idat[347:345])});
  assign Result_acc_136_nl = nl_Result_acc_136_nl[18:0];
  assign nl_Result_acc_42_nl = conv_s2u_19_21(Result_acc_136_nl) + ({(~ (data_rsci_idat[359:342]))
      , 3'b000});
  assign Result_acc_42_nl = nl_Result_acc_42_nl[20:0];
  assign nl_MultLoop_acc_374_nl = conv_s2s_12_13(Result_acc_43_itm_17_5[12:1]) +
      13'b0000011110011;
  assign MultLoop_acc_374_nl = nl_MultLoop_acc_374_nl[12:0];
  assign nl_MultLoop_acc_158_nl = conv_s2s_17_18(readslicef_20_17_3((Result_acc_56_nl)))
      + conv_s2s_15_18(readslicef_19_15_4((Result_acc_48_nl))) + conv_s2s_15_18(readslicef_25_15_10((Result_acc_32_nl)))
      + conv_s2s_15_18(readslicef_25_15_10((Result_acc_29_nl))) + conv_s2s_14_18(data_rsci_idat[125:112])
      + conv_s2s_14_18(readslicef_19_14_5((Result_acc_233_nl))) + conv_s2s_15_18(readslicef_21_15_6((Result_acc_42_nl)))
      + conv_s2s_14_18({(MultLoop_acc_374_nl) , (Result_acc_43_itm_17_5[0])});
  assign MultLoop_acc_158_nl = nl_MultLoop_acc_158_nl[17:0];
  assign nl_Result_acc_138_nl = conv_s2s_21_22({(~ (data_rsci_idat[89:72])) , 3'b001})
      + conv_s2s_18_22(Result_acc_137_cse_1);
  assign Result_acc_138_nl = nl_Result_acc_138_nl[21:0];
  assign nl_Result_acc_49_nl = conv_s2u_22_23(Result_acc_138_nl) + ({(data_rsci_idat[89:72])
      , 5'b01000});
  assign Result_acc_49_nl = nl_Result_acc_49_nl[22:0];
  assign nl_Result_acc_234_nl = conv_s2u_15_19(Result_acc_172_cse_1[18:4]) + conv_s2u_18_19(data_rsci_idat[215:198]);
  assign Result_acc_234_nl = nl_Result_acc_234_nl[18:0];
  assign nl_Result_acc_206_nl = conv_s2s_11_12(data_rsci_idat[269:259]) + 12'b000000000001;
  assign Result_acc_206_nl = nl_Result_acc_206_nl[11:0];
  assign nl_Result_acc_142_nl = conv_s2s_20_21({(data_rsci_idat[269:252]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[269:252]) + conv_s2s_17_21({(Result_acc_206_nl)
      , (data_rsci_idat[258:254])});
  assign Result_acc_142_nl = nl_Result_acc_142_nl[20:0];
  assign nl_Result_acc_37_nl = conv_s2u_21_23(Result_acc_142_nl) + ({(~ (data_rsci_idat[269:252]))
      , 5'b00000});
  assign Result_acc_37_nl = nl_Result_acc_37_nl[22:0];
  assign nl_Result_acc_143_nl = (~ (data_rsci_idat[431:414])) + conv_s2s_15_18(data_rsci_idat[431:417]);
  assign Result_acc_143_nl = nl_Result_acc_143_nl[17:0];
  assign nl_Result_acc_144_nl = conv_s2s_20_21({(~ (data_rsci_idat[431:414])) , 2'b01})
      + conv_s2s_18_21(Result_acc_143_nl);
  assign Result_acc_144_nl = nl_Result_acc_144_nl[20:0];
  assign nl_Result_acc_51_nl = conv_s2u_21_23(Result_acc_144_nl) + ({(data_rsci_idat[431:414])
      , 5'b00100});
  assign Result_acc_51_nl = nl_Result_acc_51_nl[22:0];
  assign nl_MultLoop_acc_162_nl = (MultLoop_acc_158_nl) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_49_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((Result_acc_234_nl))) + conv_s2s_16_18(readslicef_23_16_7((Result_acc_37_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_51_nl)));
  assign MultLoop_acc_162_nl = nl_MultLoop_acc_162_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl =  -conv_s2s_11_12(data_rsci_idat[17:7]);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl[11:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl = conv_s2s_25_26({(~
      (data_rsci_idat[17:0])) , 7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[17:0]))
      , 5'b00001}) + conv_s2s_19_26({(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_nl)
      , (~ (data_rsci_idat[6:0]))});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl[25:0];
  assign nl_Result_acc_145_nl = ({(data_rsci_idat[35:18]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[35:18]));
  assign Result_acc_145_nl = nl_Result_acc_145_nl[21:0];
  assign nl_Result_acc_207_nl = conv_s2u_15_19(readslicef_22_15_7((Result_acc_145_nl)))
      + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign Result_acc_207_nl = nl_Result_acc_207_nl[18:0];
  assign nl_Result_acc_208_nl = conv_s2s_11_12(data_rsci_idat[53:43]) + 12'b000000000001;
  assign Result_acc_208_nl = nl_Result_acc_208_nl[11:0];
  assign nl_Result_acc_147_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18({(Result_acc_208_nl)
      , (data_rsci_idat[42:39])});
  assign Result_acc_147_nl = nl_Result_acc_147_nl[17:0];
  assign nl_Result_acc_52_nl = conv_s2u_18_23(Result_acc_147_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[53:36])) , 4'b0001});
  assign Result_acc_52_nl = nl_Result_acc_52_nl[22:0];
  assign nl_Result_acc_148_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[71:54]));
  assign Result_acc_148_nl = nl_Result_acc_148_nl[19:0];
  assign nl_Result_acc_149_nl = ({(~ (data_rsci_idat[71:54])) , 5'b00000}) + conv_s2s_20_23(Result_acc_148_nl);
  assign Result_acc_149_nl = nl_Result_acc_149_nl[22:0];
  assign nl_Result_acc_150_nl = conv_s2s_25_26({(~ (data_rsci_idat[71:54])) , 7'b0100000})
      + conv_s2s_23_26(Result_acc_149_nl);
  assign Result_acc_150_nl = nl_Result_acc_150_nl[25:0];
  assign nl_Result_acc_209_nl = conv_s2u_19_20(readslicef_26_19_7((Result_acc_150_nl)))
      + ({(data_rsci_idat[71:54]) , 2'b01});
  assign Result_acc_209_nl = nl_Result_acc_209_nl[19:0];
  assign nl_MultLoop_acc_161_nl = conv_s2s_17_18(readslicef_26_17_9((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_1_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((Result_acc_207_nl))) + conv_s2s_17_18(readslicef_23_17_6((Result_acc_52_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((Result_acc_209_nl)));
  assign MultLoop_acc_161_nl = nl_MultLoop_acc_161_nl[17:0];
  assign nl_Result_acc_160_nl = conv_s2s_18_19(data_rsci_idat[305:288]) + conv_s2s_15_19(data_rsci_idat[305:291]);
  assign Result_acc_160_nl = nl_Result_acc_160_nl[18:0];
  assign nl_Result_acc_54_nl = conv_s2u_19_21(Result_acc_160_nl) + conv_s2u_20_21({(data_rsci_idat[305:288])
      , 2'b00});
  assign Result_acc_54_nl = nl_Result_acc_54_nl[20:0];
  assign nl_Result_acc_213_nl = conv_s2s_9_10(data_rsci_idat[323:315]) + 10'b0000000001;
  assign Result_acc_213_nl = nl_Result_acc_213_nl[9:0];
  assign nl_Result_acc_163_nl = conv_s2s_22_23({(data_rsci_idat[323:306]) , 4'b0000})
      + conv_s2s_18_23(data_rsci_idat[323:306]) + conv_s2s_16_23({(Result_acc_213_nl)
      , (data_rsci_idat[314:309])});
  assign Result_acc_163_nl = nl_Result_acc_163_nl[22:0];
  assign nl_Result_acc_214_nl = conv_s2u_17_18(readslicef_23_17_6((Result_acc_163_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign Result_acc_214_nl = nl_Result_acc_214_nl[17:0];
  assign nl_Result_acc_215_nl = conv_s2s_9_10(data_rsci_idat[341:333]) + 10'b0000000001;
  assign Result_acc_215_nl = nl_Result_acc_215_nl[9:0];
  assign nl_Result_acc_165_nl = (~ (data_rsci_idat[341:324])) + conv_s2s_15_18({(Result_acc_215_nl)
      , (data_rsci_idat[332:328])});
  assign Result_acc_165_nl = nl_Result_acc_165_nl[17:0];
  assign nl_Result_acc_166_nl = ({(data_rsci_idat[341:324]) , 3'b001}) + conv_s2s_18_21(Result_acc_165_nl);
  assign Result_acc_166_nl = nl_Result_acc_166_nl[20:0];
  assign nl_Result_acc_41_nl = conv_s2u_21_23(Result_acc_166_nl) + ({(~ (data_rsci_idat[341:324]))
      , 5'b00000});
  assign Result_acc_41_nl = nl_Result_acc_41_nl[22:0];
  assign nl_Result_acc_216_nl = conv_s2s_13_14(data_rsci_idat[395:383]) + 14'b00000000000001;
  assign Result_acc_216_nl = nl_Result_acc_216_nl[13:0];
  assign nl_Result_acc_168_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_17_18({(Result_acc_216_nl)
      , (data_rsci_idat[382:380])});
  assign Result_acc_168_nl = nl_Result_acc_168_nl[17:0];
  assign nl_Result_acc_55_nl = conv_s2u_18_22(Result_acc_168_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[395:378])) , 3'b001});
  assign Result_acc_55_nl = nl_Result_acc_55_nl[21:0];
  assign nl_MultLoop_acc_159_nl = conv_s2s_17_18(readslicef_21_17_4((Result_acc_54_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((Result_acc_214_nl))) + conv_s2s_17_18(readslicef_23_17_6((Result_acc_41_nl)))
      + conv_s2s_17_18(readslicef_22_17_5((Result_acc_55_nl)));
  assign MultLoop_acc_159_nl = nl_MultLoop_acc_159_nl[17:0];
  assign nl_Result_acc_151_nl = (~ (data_rsci_idat[197:180])) + conv_s2s_16_18(data_rsci_idat[197:182]);
  assign Result_acc_151_nl = nl_Result_acc_151_nl[17:0];
  assign nl_Result_acc_152_nl = ({(data_rsci_idat[197:180]) , 3'b001}) + conv_s2s_18_21(Result_acc_151_nl);
  assign Result_acc_152_nl = nl_Result_acc_152_nl[20:0];
  assign nl_Result_acc_53_nl = conv_s2u_21_24(Result_acc_152_nl) + conv_s2u_23_24({(data_rsci_idat[197:180])
      , 5'b00000});
  assign Result_acc_53_nl = nl_Result_acc_53_nl[23:0];
  assign nl_Result_acc_210_nl = conv_s2s_9_10(data_rsci_idat[233:225]) + 10'b0000000001;
  assign Result_acc_210_nl = nl_Result_acc_210_nl[9:0];
  assign nl_Result_acc_156_nl = conv_s2s_22_23({(data_rsci_idat[233:216]) , 4'b0000})
      + conv_s2s_20_23({(data_rsci_idat[233:216]) , 2'b00}) + conv_s2s_18_23(data_rsci_idat[233:216])
      + conv_s2s_16_23({(Result_acc_210_nl) , (data_rsci_idat[224:219])});
  assign Result_acc_156_nl = nl_Result_acc_156_nl[22:0];
  assign nl_Result_acc_211_nl = conv_s2u_17_18(readslicef_23_17_6((Result_acc_156_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign Result_acc_211_nl = nl_Result_acc_211_nl[17:0];
  assign nl_Result_acc_235_nl = conv_s2u_18_19(data_rsci_idat[251:234]) + conv_s2u_15_19(MultLoop_acc_263_cse_1[19:5]);
  assign Result_acc_235_nl = nl_Result_acc_235_nl[18:0];
  assign nl_Result_acc_212_nl = conv_s2u_17_19(readslicef_19_17_2((Result_acc_235_nl)))
      + conv_s2u_18_19(data_rsci_idat[251:234]);
  assign Result_acc_212_nl = nl_Result_acc_212_nl[18:0];
  assign nl_Result_acc_159_nl = ({(data_rsci_idat[287:270]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[287:270]));
  assign Result_acc_159_nl = nl_Result_acc_159_nl[19:0];
  assign nl_Result_acc_38_nl = conv_s2s_20_23(Result_acc_159_nl) + conv_s2s_22_23({(data_rsci_idat[287:270])
      , 4'b0000});
  assign Result_acc_38_nl = nl_Result_acc_38_nl[22:0];
  assign nl_res_rsci_d_89_72  = (MultLoop_acc_162_nl) + (MultLoop_acc_161_nl) + (MultLoop_acc_159_nl)
      + conv_s2s_17_18(readslicef_24_17_7((Result_acc_53_nl))) + conv_s2s_17_18(readslicef_18_17_1((Result_acc_211_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((Result_acc_212_nl))) + conv_s2s_17_18(readslicef_23_17_6((Result_acc_38_nl)));
  assign nl_MultLoop_acc_368_nl = conv_s2u_17_19(MultLoop_acc_72_itm_23_7) + conv_s2u_18_19(data_rsci_idat[341:324]);
  assign MultLoop_acc_368_nl = nl_MultLoop_acc_368_nl[18:0];
  assign nl_MultLoop_acc_369_nl = conv_s2s_13_14(data_rsci_idat[269:257]) + 14'b00000000000001;
  assign MultLoop_acc_369_nl = nl_MultLoop_acc_369_nl[13:0];
  assign nl_MultLoop_acc_253_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_17_18({(MultLoop_acc_369_nl)
      , (data_rsci_idat[256:254])});
  assign MultLoop_acc_253_nl = nl_MultLoop_acc_253_nl[17:0];
  assign nl_MultLoop_acc_101_nl = conv_s2u_18_22(MultLoop_acc_253_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[269:252])) , 3'b001});
  assign MultLoop_acc_101_nl = nl_MultLoop_acc_101_nl[21:0];
  assign nl_MultLoop_acc_243_nl = conv_s2s_21_22({(~ (data_rsci_idat[107:90])) ,
      3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_243_nl = nl_MultLoop_acc_243_nl[21:0];
  assign nl_MultLoop_acc_35_nl = conv_s2s_22_25(MultLoop_acc_243_nl) + ({(data_rsci_idat[107:90])
      , 7'b0001000});
  assign MultLoop_acc_35_nl = nl_MultLoop_acc_35_nl[24:0];
  assign nl_MultLoop_acc_365_nl =  -conv_s2s_12_13(data_rsci_idat[17:6]);
  assign MultLoop_acc_365_nl = nl_MultLoop_acc_365_nl[12:0];
  assign nl_MultLoop_acc_245_nl = ({(data_rsci_idat[17:0]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_365_nl)
      , (~ (data_rsci_idat[5:0]))});
  assign MultLoop_acc_245_nl = nl_MultLoop_acc_245_nl[19:0];
  assign nl_MultLoop_acc_366_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_245_nl)))
      + (~ (data_rsci_idat[17:0]));
  assign MultLoop_acc_366_nl = nl_MultLoop_acc_366_nl[17:0];
  assign nl_MultLoop_acc_247_nl = ({(~ (data_rsci_idat[413:396])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_76_cse_1);
  assign MultLoop_acc_247_nl = nl_MultLoop_acc_247_nl[21:0];
  assign nl_MultLoop_acc_50_nl = conv_s2s_22_25(MultLoop_acc_247_nl) + ({(data_rsci_idat[413:396])
      , 7'b0010000});
  assign MultLoop_acc_50_nl = nl_MultLoop_acc_50_nl[24:0];
  assign nl_MultLoop_acc_367_nl = conv_s2s_11_12(data_rsci_idat[377:367]) + 12'b000000000001;
  assign MultLoop_acc_367_nl = nl_MultLoop_acc_367_nl[11:0];
  assign nl_MultLoop_acc_249_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_17_18({(MultLoop_acc_367_nl)
      , (data_rsci_idat[366:362])});
  assign MultLoop_acc_249_nl = nl_MultLoop_acc_249_nl[17:0];
  assign nl_MultLoop_acc_104_nl = conv_s2u_18_24(MultLoop_acc_249_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[377:360])) , 5'b00001});
  assign MultLoop_acc_104_nl = nl_MultLoop_acc_104_nl[23:0];
  assign nl_MultLoop_acc_254_nl = conv_s2s_20_21({(~ (data_rsci_idat[233:216])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_254_nl = nl_MultLoop_acc_254_nl[20:0];
  assign nl_MultLoop_acc_41_nl = conv_s2s_21_26(MultLoop_acc_254_nl) + ({(data_rsci_idat[233:216])
      , 8'b00000100});
  assign MultLoop_acc_41_nl = nl_MultLoop_acc_41_nl[25:0];
  assign nl_MultLoop_acc_370_nl =  -conv_s2s_11_12(data_rsci_idat[179:169]);
  assign MultLoop_acc_370_nl = nl_MultLoop_acc_370_nl[11:0];
  assign nl_MultLoop_acc_38_nl = conv_s2s_25_26({(~ (data_rsci_idat[179:162])) ,
      7'b0000100}) + conv_s2s_20_26({(~ (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_26({(MultLoop_acc_370_nl)
      , (~ (data_rsci_idat[168:162]))});
  assign MultLoop_acc_38_nl = nl_MultLoop_acc_38_nl[25:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_368_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_101_nl))) + conv_s2s_15_18(~
      (data_rsci_idat[53:39])) + conv_s2s_15_18(~ (data_rsci_idat[125:111])) + conv_s2s_15_18(readslicef_25_15_10((MultLoop_acc_35_nl)))
      + conv_s2s_15_18(readslicef_18_15_3((MultLoop_acc_366_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_50_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_104_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_41_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_38_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl[17:0];
  assign nl_MultLoop_acc_257_nl = ({(data_rsci_idat[359:342]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[359:342]));
  assign MultLoop_acc_257_nl = nl_MultLoop_acc_257_nl[20:0];
  assign nl_MultLoop_acc_258_nl = ({(~ (data_rsci_idat[359:342])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_257_nl);
  assign MultLoop_acc_258_nl = nl_MultLoop_acc_258_nl[22:0];
  assign nl_MultLoop_acc_48_nl = conv_s2s_23_25(MultLoop_acc_258_nl) + ({(data_rsci_idat[359:342])
      , 7'b0100000});
  assign MultLoop_acc_48_nl = nl_MultLoop_acc_48_nl[24:0];
  assign nl_MultLoop_acc_260_nl = ({(~ (data_rsci_idat[305:288])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_395);
  assign MultLoop_acc_260_nl = nl_MultLoop_acc_260_nl[21:0];
  assign nl_MultLoop_acc_45_nl = conv_s2s_22_24(MultLoop_acc_260_nl) + ({(data_rsci_idat[305:288])
      , 6'b010000});
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[23:0];
  assign nl_MultLoop_acc_261_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_16_18(data_rsci_idat[323:308]);
  assign MultLoop_acc_261_nl = nl_MultLoop_acc_261_nl[17:0];
  assign nl_MultLoop_acc_262_nl = ({(data_rsci_idat[323:306]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_261_nl);
  assign MultLoop_acc_262_nl = nl_MultLoop_acc_262_nl[19:0];
  assign nl_MultLoop_acc_103_nl = conv_s2u_20_23(MultLoop_acc_262_nl) + conv_s2u_22_23({(data_rsci_idat[323:306])
      , 4'b0000});
  assign MultLoop_acc_103_nl = nl_MultLoop_acc_103_nl[22:0];
  assign nl_MultLoop_acc_32_nl = conv_s2s_18_23(~ (data_rsci_idat[35:18])) + ({(data_rsci_idat[35:18])
      , 5'b00001});
  assign MultLoop_acc_32_nl = nl_MultLoop_acc_32_nl[22:0];
  assign nl_MultLoop_acc_242_nl = conv_s2s_18_19(data_rsci_idat[431:414]) + conv_s2s_16_19(data_rsci_idat[431:416]);
  assign MultLoop_acc_242_nl = nl_MultLoop_acc_242_nl[18:0];
  assign nl_MultLoop_acc_105_nl = conv_s2u_19_22(MultLoop_acc_242_nl) + conv_s2u_21_22({(data_rsci_idat[431:414])
      , 3'b000});
  assign MultLoop_acc_105_nl = nl_MultLoop_acc_105_nl[21:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl = ~((data_rsci_idat[385:378]!=8'b00000000));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl = ~((data_rsci_idat[110:108]!=3'b000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl = conv_u2u_10_11({9'b100001110
      , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl)}) + conv_s2u_10_11(~
      (data_rsci_idat[395:386])) + conv_u2u_1_11(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl[10:0];
  assign nl_MultLoop_acc_102_nl = conv_s2u_16_19(data_rsci_idat[287:272]) + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_102_nl = nl_MultLoop_acc_102_nl[18:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl = ~((data_rsci_idat[38:36]!=3'b000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl = conv_u2s_11_13(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_27_nl)
      + conv_s2s_11_13(readslicef_19_11_8((MultLoop_acc_102_nl))) + conv_u2s_1_13(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl[12:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_48_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_45_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_103_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_32_nl))) + conv_s2s_14_18(readslicef_22_14_8((MultLoop_acc_105_nl)))
      + conv_s2s_13_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_28_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl[17:0];
  assign nl_MultLoop_acc_272_nl = conv_s2s_24_25({(~ (data_rsci_idat[143:126])) ,
      6'b000001}) + conv_s2s_18_25(~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_272_nl = nl_MultLoop_acc_272_nl[24:0];
  assign nl_MultLoop_acc_36_nl = conv_s2s_25_27(MultLoop_acc_272_nl) + ({(data_rsci_idat[143:126])
      , 9'b001000000});
  assign MultLoop_acc_36_nl = nl_MultLoop_acc_36_nl[26:0];
  assign nl_MultLoop_acc_373_nl = conv_s2s_12_13(data_rsci_idat[71:60]) + 13'b0000000000001;
  assign MultLoop_acc_373_nl = nl_MultLoop_acc_373_nl[12:0];
  assign nl_MultLoop_acc_274_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({(MultLoop_acc_373_nl)
      , (data_rsci_idat[59:56])});
  assign MultLoop_acc_274_nl = nl_MultLoop_acc_274_nl[17:0];
  assign nl_MultLoop_acc_275_nl = conv_s2s_20_21({(~ (data_rsci_idat[71:54])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_274_nl);
  assign MultLoop_acc_275_nl = nl_MultLoop_acc_275_nl[20:0];
  assign nl_MultLoop_acc_98_nl = conv_s2u_21_23(MultLoop_acc_275_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[71:54])) , 4'b0100});
  assign MultLoop_acc_98_nl = nl_MultLoop_acc_98_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_36_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_98_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl[17:0];
  assign nl_MultLoop_acc_99_nl = conv_s2u_9_19(data_rsci_idat[89:81]) + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_99_nl = nl_MultLoop_acc_99_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_37_nl)
      + (readslicef_19_18_1((MultLoop_acc_99_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl[17:0];
  assign nl_MultLoop_acc_264_nl = ({(~ (data_rsci_idat[251:234])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_263_cse_1);
  assign MultLoop_acc_264_nl = nl_MultLoop_acc_264_nl[21:0];
  assign nl_MultLoop_acc_42_nl = conv_s2s_22_27(MultLoop_acc_264_nl) + ({(data_rsci_idat[251:234])
      , 9'b000010000});
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[26:0];
  assign nl_MultLoop_acc_266_nl = ({(~ (data_rsci_idat[197:180])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[197:180])
      + conv_s2s_14_21(data_rsci_idat[197:184]);
  assign MultLoop_acc_266_nl = nl_MultLoop_acc_266_nl[20:0];
  assign nl_MultLoop_acc_100_nl = conv_s2u_21_23(MultLoop_acc_266_nl) + ({(data_rsci_idat[197:180])
      , 5'b01000});
  assign MultLoop_acc_100_nl = nl_MultLoop_acc_100_nl[22:0];
  assign nl_MultLoop_acc_371_nl =  -conv_s2s_11_12(data_rsci_idat[215:205]);
  assign MultLoop_acc_371_nl = nl_MultLoop_acc_371_nl[11:0];
  assign nl_MultLoop_acc_40_nl = conv_s2s_25_26({(~ (data_rsci_idat[215:198])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[215:198])) , 5'b00001}) +
      conv_s2s_19_26({(MultLoop_acc_371_nl) , (~ (data_rsci_idat[204:198]))});
  assign MultLoop_acc_40_nl = nl_MultLoop_acc_40_nl[25:0];
  assign nl_MultLoop_acc_270_nl = ({(~ (data_rsci_idat[161:144])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_193_cse_1);
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[21:0];
  assign nl_MultLoop_acc_271_nl = ({(data_rsci_idat[161:144]) , 6'b010000}) + conv_s2s_22_24(MultLoop_acc_270_nl);
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[23:0];
  assign nl_MultLoop_acc_372_nl = conv_s2u_16_19(readslicef_24_16_8((MultLoop_acc_271_nl)))
      + conv_s2u_18_19(data_rsci_idat[161:144]);
  assign MultLoop_acc_372_nl = nl_MultLoop_acc_372_nl[18:0];
  assign nl_res_rsci_d_35_18  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_46_nl) + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_44_nl)
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_42_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_100_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_40_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_372_nl)));
  assign nl_Result_acc_196_nl =  -conv_s2s_9_10(data_rsci_idat[395:387]);
  assign Result_acc_196_nl = nl_Result_acc_196_nl[9:0];
  assign nl_Result_acc_194_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_19_20({(Result_acc_196_nl)
      , (~ (data_rsci_idat[386:378]))});
  assign Result_acc_194_nl = nl_Result_acc_194_nl[19:0];
  assign nl_Result_acc_197_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_13_18(readslicef_20_13_7((Result_acc_194_nl)));
  assign Result_acc_197_nl = nl_Result_acc_197_nl[17:0];
  assign nl_Result_acc_198_nl = conv_s2u_18_21(Result_acc_197_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[395:378])) , 2'b01});
  assign Result_acc_198_nl = nl_Result_acc_198_nl[20:0];
  assign nl_Result_acc_171_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_16_19(data_rsci_idat[161:146]);
  assign Result_acc_171_nl = nl_Result_acc_171_nl[18:0];
  assign nl_Result_acc_16_nl = conv_s2u_19_21(Result_acc_171_nl) + conv_s2u_20_21({(data_rsci_idat[161:144])
      , 2'b00});
  assign Result_acc_16_nl = nl_Result_acc_16_nl[20:0];
  assign nl_Result_acc_173_nl = ({(~ (data_rsci_idat[215:198])) , 3'b000}) + conv_s2s_19_21(Result_acc_172_cse_1);
  assign Result_acc_173_nl = nl_Result_acc_173_nl[20:0];
  assign nl_Result_acc_17_nl = conv_s2u_21_24(Result_acc_173_nl) + ({(data_rsci_idat[215:198])
      , 6'b001000});
  assign Result_acc_17_nl = nl_Result_acc_17_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = conv_s2s_16_17(readslicef_21_16_5((Result_acc_16_nl)))
      + conv_s2s_16_17(readslicef_24_16_8((Result_acc_17_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl = (readslicef_21_18_3((Result_acc_198_nl)))
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl[17:0];
  assign nl_Result_acc_175_nl = ({(~ (data_rsci_idat[251:234])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[251:234])
      + conv_s2s_15_21(data_rsci_idat[251:237]);
  assign Result_acc_175_nl = nl_Result_acc_175_nl[20:0];
  assign nl_Result_acc_18_nl = conv_s2u_21_23(Result_acc_175_nl) + ({(data_rsci_idat[251:234])
      , 5'b01000});
  assign Result_acc_18_nl = nl_Result_acc_18_nl[22:0];
  assign nl_Result_acc_199_nl =  -conv_s2s_11_12(data_rsci_idat[269:259]);
  assign Result_acc_199_nl = nl_Result_acc_199_nl[11:0];
  assign nl_Result_acc_177_nl = ({(data_rsci_idat[269:252]) , 3'b001}) + conv_s2s_19_21({(Result_acc_199_nl)
      , (~ (data_rsci_idat[258:252]))});
  assign Result_acc_177_nl = nl_Result_acc_177_nl[20:0];
  assign nl_Result_acc_178_nl = conv_s2s_23_24({(data_rsci_idat[269:252]) , 5'b00000})
      + conv_s2s_21_24(Result_acc_177_nl);
  assign Result_acc_178_nl = nl_Result_acc_178_nl[23:0];
  assign nl_Result_acc_200_nl = conv_s2u_17_18(readslicef_24_17_7((Result_acc_178_nl)))
      + (~ (data_rsci_idat[269:252]));
  assign Result_acc_200_nl = nl_Result_acc_200_nl[17:0];
  assign nl_Result_acc_179_nl = (~ (data_rsci_idat[287:270])) + conv_s2s_15_18(data_rsci_idat[287:273]);
  assign Result_acc_179_nl = nl_Result_acc_179_nl[17:0];
  assign nl_Result_acc_19_nl = conv_s2u_18_21(Result_acc_179_nl) + ({(data_rsci_idat[287:270])
      , 3'b001});
  assign Result_acc_19_nl = nl_Result_acc_19_nl[20:0];
  assign nl_Result_acc_180_nl = conv_s2s_18_19(data_rsci_idat[431:414]) + conv_s2s_15_19(data_rsci_idat[431:417]);
  assign Result_acc_180_nl = nl_Result_acc_180_nl[18:0];
  assign nl_Result_acc_20_nl = conv_s2u_19_21(Result_acc_180_nl) + conv_s2u_20_21({(data_rsci_idat[431:414])
      , 2'b00});
  assign Result_acc_20_nl = nl_Result_acc_20_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl)
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_18_nl))) + conv_s2s_16_18(readslicef_18_16_2((Result_acc_200_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((Result_acc_19_nl))) + conv_s2s_16_18(readslicef_21_16_5((Result_acc_20_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl[17:0];
  assign nl_Result_acc_181_nl = conv_s2s_18_19(data_rsci_idat[179:162]) + conv_s2s_14_19(data_rsci_idat[179:166]);
  assign Result_acc_181_nl = nl_Result_acc_181_nl[18:0];
  assign nl_Result_acc_21_nl = conv_s2u_19_23(Result_acc_181_nl) + conv_s2u_22_23({(data_rsci_idat[179:162])
      , 4'b0000});
  assign Result_acc_21_nl = nl_Result_acc_21_nl[22:0];
  assign nl_Result_acc_183_nl = conv_s2s_22_23({(~ (data_rsci_idat[197:180])) , 4'b0100})
      + conv_s2s_20_23({(~ (data_rsci_idat[197:180])) , 2'b01}) + conv_s2s_18_23(~
      (data_rsci_idat[197:180]));
  assign Result_acc_183_nl = nl_Result_acc_183_nl[22:0];
  assign nl_Result_acc_3_nl = conv_s2s_23_26(Result_acc_183_nl) + ({(data_rsci_idat[197:180])
      , 8'b00010000});
  assign Result_acc_3_nl = nl_Result_acc_3_nl[25:0];
  assign nl_Result_acc_184_nl = (~ (data_rsci_idat[305:288])) + conv_s2s_16_18(data_rsci_idat[305:290]);
  assign Result_acc_184_nl = nl_Result_acc_184_nl[17:0];
  assign nl_Result_acc_185_nl = conv_s2s_21_22({(~ (data_rsci_idat[305:288])) , 3'b001})
      + conv_s2s_18_22(Result_acc_184_nl);
  assign Result_acc_185_nl = nl_Result_acc_185_nl[21:0];
  assign nl_Result_acc_22_nl = conv_s2u_22_23(Result_acc_185_nl) + ({(data_rsci_idat[305:288])
      , 5'b01000});
  assign Result_acc_22_nl = nl_Result_acc_22_nl[22:0];
  assign nl_MultLoop_acc_114_nl = conv_s2u_14_19(data_rsci_idat[89:76]) + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_114_nl = nl_MultLoop_acc_114_nl[18:0];
  assign nl_Result_acc_170_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_16_18(data_rsci_idat[233:218]);
  assign Result_acc_170_nl = nl_Result_acc_170_nl[17:0];
  assign nl_Result_acc_nl = conv_s2u_18_23(Result_acc_170_nl) + ({(data_rsci_idat[233:216])
      , 5'b00001});
  assign Result_acc_nl = nl_Result_acc_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl = conv_s2s_17_18(readslicef_23_17_6((Result_acc_21_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((Result_acc_3_nl))) + conv_s2s_17_18(readslicef_23_17_6((Result_acc_22_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_114_nl))) + conv_s2s_15_18(readslicef_23_15_8((Result_acc_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl[17:0];
  assign nl_MultLoop_acc_359_nl =  -conv_s2s_9_10(data_rsci_idat[125:117]);
  assign MultLoop_acc_359_nl = nl_MultLoop_acc_359_nl[9:0];
  assign nl_MultLoop_acc_169_nl = ({(data_rsci_idat[125:108]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_359_nl)
      , (~ (data_rsci_idat[116:108]))});
  assign MultLoop_acc_169_nl = nl_MultLoop_acc_169_nl[19:0];
  assign nl_MultLoop_acc_360_nl = conv_s2u_11_18(readslicef_20_11_9((MultLoop_acc_169_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_360_nl = nl_MultLoop_acc_360_nl[17:0];
  assign nl_MultLoop_acc_361_nl =  -conv_s2s_11_12(data_rsci_idat[53:43]);
  assign MultLoop_acc_361_nl = nl_MultLoop_acc_361_nl[11:0];
  assign nl_MultLoop_acc_171_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_361_nl)
      , (~ (data_rsci_idat[42:36]))});
  assign MultLoop_acc_171_nl = nl_MultLoop_acc_171_nl[20:0];
  assign nl_MultLoop_acc_172_nl = conv_s2s_23_24({(data_rsci_idat[53:36]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_171_nl);
  assign MultLoop_acc_172_nl = nl_MultLoop_acc_172_nl[23:0];
  assign nl_MultLoop_acc_362_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_172_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_362_nl = nl_MultLoop_acc_362_nl[17:0];
  assign nl_MultLoop_acc_175_nl = conv_s2s_20_21({(~ (data_rsci_idat[71:54])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_174_cse_1);
  assign MultLoop_acc_175_nl = nl_MultLoop_acc_175_nl[20:0];
  assign nl_MultLoop_acc_113_nl = conv_s2u_21_25(MultLoop_acc_175_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[71:54])) , 6'b000100});
  assign MultLoop_acc_113_nl = nl_MultLoop_acc_113_nl[24:0];
  assign nl_MultLoop_acc_364_nl =  -conv_s2s_13_14(data_rsci_idat[17:5]);
  assign MultLoop_acc_364_nl = nl_MultLoop_acc_364_nl[13:0];
  assign nl_MultLoop_acc_167_nl = ({(data_rsci_idat[17:0]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_364_nl)
      , (~ (data_rsci_idat[4:0]))});
  assign MultLoop_acc_167_nl = nl_MultLoop_acc_167_nl[20:0];
  assign nl_MultLoop_acc_78_nl = conv_s2s_21_23(MultLoop_acc_167_nl) + ({(~ (data_rsci_idat[17:0]))
      , 5'b00000});
  assign MultLoop_acc_78_nl = nl_MultLoop_acc_78_nl[22:0];
  assign nl_MultLoop_acc_165_nl = conv_s2s_20_21({(~ (data_rsci_idat[107:90])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_165_nl = nl_MultLoop_acc_165_nl[20:0];
  assign nl_MultLoop_acc_84_nl = conv_s2s_21_23(MultLoop_acc_165_nl) + ({(data_rsci_idat[107:90])
      , 5'b00100});
  assign MultLoop_acc_84_nl = nl_MultLoop_acc_84_nl[22:0];
  assign nl_MultLoop_acc_86_nl = conv_s2u_15_18(data_rsci_idat[143:129]) - (data_rsci_idat[143:126]);
  assign MultLoop_acc_86_nl = nl_MultLoop_acc_86_nl[17:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl = ~((data_rsci_idat[350:342]!=9'b000000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl = conv_s2s_9_10(~
      (data_rsci_idat[359:351])) + conv_u2s_8_10({7'b1110010 , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl)});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl[9:0];
  assign nl_MultLoop_acc_80_nl = conv_s2s_18_20(~ (data_rsci_idat[35:18])) + ({(data_rsci_idat[35:18])
      , 2'b01});
  assign MultLoop_acc_80_nl = nl_MultLoop_acc_80_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl = conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_360_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_362_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_113_nl)))
      + conv_s2s_15_18(readslicef_23_15_8((MultLoop_acc_78_nl))) + conv_s2s_13_18(readslicef_23_13_10((MultLoop_acc_84_nl)))
      + conv_s2s_11_18(readslicef_18_11_7((MultLoop_acc_86_nl))) + conv_s2s_10_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_4_nl)
      + conv_s2s_10_18(readslicef_20_10_10((MultLoop_acc_80_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl[17:0];
  assign nl_Result_acc_187_nl = conv_s2s_20_21({(data_rsci_idat[323:306]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[323:306]) + conv_s2s_15_21(data_rsci_idat[323:309]);
  assign Result_acc_187_nl = nl_Result_acc_187_nl[20:0];
  assign nl_Result_acc_23_nl = conv_s2u_21_24(Result_acc_187_nl) + conv_s2u_23_24({(data_rsci_idat[323:306])
      , 5'b00000});
  assign Result_acc_23_nl = nl_Result_acc_23_nl[23:0];
  assign nl_Result_acc_201_nl =  -conv_s2s_11_12(data_rsci_idat[341:331]);
  assign Result_acc_201_nl = nl_Result_acc_201_nl[11:0];
  assign nl_Result_acc_11_nl = conv_s2s_19_26({(Result_acc_201_nl) , (~ (data_rsci_idat[330:324]))})
      + conv_s2s_25_26({(~ (data_rsci_idat[341:324])) , 7'b0000001});
  assign Result_acc_11_nl = nl_Result_acc_11_nl[25:0];
  assign nl_Result_acc_190_nl = conv_s2s_25_26({(~ (data_rsci_idat[377:360])) , 7'b0001000})
      + conv_s2s_21_26({(~ (data_rsci_idat[377:360])) , 3'b001}) + conv_s2s_18_26(~
      (data_rsci_idat[377:360]));
  assign Result_acc_190_nl = nl_Result_acc_190_nl[25:0];
  assign nl_Result_acc_202_nl = conv_s2u_19_20(readslicef_26_19_7((Result_acc_190_nl)))
      + ({(data_rsci_idat[377:360]) , 2'b01});
  assign Result_acc_202_nl = nl_Result_acc_202_nl[19:0];
  assign nl_Result_acc_203_nl = conv_s2s_13_14(data_rsci_idat[413:401]) + 14'b00000000000001;
  assign Result_acc_203_nl = nl_Result_acc_203_nl[13:0];
  assign nl_Result_acc_192_nl = (~ (data_rsci_idat[413:396])) + conv_s2s_16_18({(Result_acc_203_nl)
      , (data_rsci_idat[400:399])});
  assign Result_acc_192_nl = nl_Result_acc_192_nl[17:0];
  assign nl_Result_acc_24_nl = conv_s2u_18_21(Result_acc_192_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[413:396])) , 2'b01});
  assign Result_acc_24_nl = nl_Result_acc_24_nl[20:0];
  assign nl_res_rsci_d_71_54  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_24_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_nl) + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_21_nl)
      + conv_s2s_17_18(readslicef_24_17_7((Result_acc_23_nl))) + conv_s2s_17_18(readslicef_26_17_9((Result_acc_11_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((Result_acc_202_nl))) + conv_s2s_17_18(readslicef_21_17_4((Result_acc_24_nl)));
  assign nl_MultLoop_acc_192_nl = conv_s2s_23_24({(~ (data_rsci_idat[215:198])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[215:198])) , 2'b01}) + conv_s2s_18_24(~
      (data_rsci_idat[215:198]));
  assign MultLoop_acc_192_nl = nl_MultLoop_acc_192_nl[23:0];
  assign nl_MultLoop_acc_65_nl = conv_s2s_24_26(MultLoop_acc_192_nl) + ({(data_rsci_idat[215:198])
      , 8'b00100000});
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[25:0];
  assign nl_MultLoop_acc_393_nl = conv_s2u_15_19(MultLoop_acc_193_cse_1[19:5]) +
      conv_s2u_18_19(data_rsci_idat[161:144]);
  assign MultLoop_acc_393_nl = nl_MultLoop_acc_393_nl[18:0];
  assign nl_MultLoop_acc_346_nl =  -conv_s2s_12_13(data_rsci_idat[269:258]);
  assign MultLoop_acc_346_nl = nl_MultLoop_acc_346_nl[12:0];
  assign nl_MultLoop_acc_68_nl = conv_s2s_24_25({(~ (data_rsci_idat[269:252])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[269:252])) , 3'b001}) + conv_s2s_19_25({(MultLoop_acc_346_nl)
      , (~ (data_rsci_idat[257:252]))});
  assign MultLoop_acc_68_nl = nl_MultLoop_acc_68_nl[24:0];
  assign nl_MultLoop_acc_347_nl =  -conv_s2s_11_12(data_rsci_idat[287:277]);
  assign MultLoop_acc_347_nl = nl_MultLoop_acc_347_nl[11:0];
  assign nl_MultLoop_acc_188_nl = ({(data_rsci_idat[287:270]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_347_nl)
      , (~ (data_rsci_idat[276:270]))});
  assign MultLoop_acc_188_nl = nl_MultLoop_acc_188_nl[21:0];
  assign nl_MultLoop_acc_348_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_188_nl)))
      + (~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_348_nl = nl_MultLoop_acc_348_nl[17:0];
  assign nl_MultLoop_acc_189_nl = ({(data_rsci_idat[233:216]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[233:216]));
  assign MultLoop_acc_189_nl = nl_MultLoop_acc_189_nl[20:0];
  assign nl_MultLoop_acc_190_nl = ({(~ (data_rsci_idat[233:216])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_189_nl);
  assign MultLoop_acc_190_nl = nl_MultLoop_acc_190_nl[22:0];
  assign nl_MultLoop_acc_66_nl = conv_s2s_23_25(MultLoop_acc_190_nl) + ({(data_rsci_idat[233:216])
      , 7'b0100000});
  assign MultLoop_acc_66_nl = nl_MultLoop_acc_66_nl[24:0];
  assign nl_MultLoop_acc_349_nl = conv_s2s_12_13(data_rsci_idat[143:132]) + 13'b0000000000001;
  assign MultLoop_acc_349_nl = nl_MultLoop_acc_349_nl[12:0];
  assign nl_MultLoop_acc_195_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_16_18({(MultLoop_acc_349_nl)
      , (data_rsci_idat[131:129])});
  assign MultLoop_acc_195_nl = nl_MultLoop_acc_195_nl[17:0];
  assign nl_MultLoop_acc_108_nl = conv_s2u_18_22(MultLoop_acc_195_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[143:126])) , 3'b001});
  assign MultLoop_acc_108_nl = nl_MultLoop_acc_108_nl[21:0];
  assign nl_MultLoop_acc_77_nl = conv_s2s_24_25({(~ (data_rsci_idat[431:414])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[431:414])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[431:414])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_50_18_6
      , (~ (data_rsci_idat[419:414]))});
  assign MultLoop_acc_77_nl = nl_MultLoop_acc_77_nl[24:0];
  assign nl_MultLoop_acc_238_nl = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_65_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_393_nl))) + conv_s2s_16_18(MultLoop_acc_76_cse_1[19:4])
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_68_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_348_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_66_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_108_nl)))
      + conv_s2s_15_18(readslicef_25_15_10((MultLoop_acc_77_nl)));
  assign MultLoop_acc_238_nl = nl_MultLoop_acc_238_nl[17:0];
  assign nl_MultLoop_acc_356_nl = conv_s2s_11_12(data_rsci_idat[251:241]) + 12'b000000000001;
  assign MultLoop_acc_356_nl = nl_MultLoop_acc_356_nl[11:0];
  assign nl_MultLoop_acc_206_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_17_18({(MultLoop_acc_356_nl)
      , (data_rsci_idat[240:236])});
  assign MultLoop_acc_206_nl = nl_MultLoop_acc_206_nl[17:0];
  assign nl_MultLoop_acc_110_nl = conv_s2u_18_24(MultLoop_acc_206_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[251:234])) , 5'b00001});
  assign MultLoop_acc_110_nl = nl_MultLoop_acc_110_nl[23:0];
  assign nl_MultLoop_acc_207_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18(data_rsci_idat[179:164]);
  assign MultLoop_acc_207_nl = nl_MultLoop_acc_207_nl[17:0];
  assign nl_MultLoop_acc_208_nl = conv_s2s_22_23({(~ (data_rsci_idat[179:162])) ,
      4'b0001}) + conv_s2s_18_23(MultLoop_acc_207_nl);
  assign MultLoop_acc_208_nl = nl_MultLoop_acc_208_nl[22:0];
  assign nl_MultLoop_acc_109_nl = conv_s2u_23_24(MultLoop_acc_208_nl) + ({(data_rsci_idat[179:162])
      , 6'b010000});
  assign MultLoop_acc_109_nl = nl_MultLoop_acc_109_nl[23:0];
  assign nl_MultLoop_acc_357_nl =  -conv_s2s_9_10(data_rsci_idat[107:99]);
  assign MultLoop_acc_357_nl = nl_MultLoop_acc_357_nl[9:0];
  assign nl_MultLoop_acc_212_nl = ({(data_rsci_idat[107:90]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[107:90])) , 4'b0100}) + conv_s2s_20_24({(~ (data_rsci_idat[107:90]))
      , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_357_nl) , (~ (data_rsci_idat[98:90]))});
  assign MultLoop_acc_212_nl = nl_MultLoop_acc_212_nl[23:0];
  assign nl_MultLoop_acc_358_nl = conv_s2u_15_18(readslicef_24_15_9((MultLoop_acc_212_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_358_nl = nl_MultLoop_acc_358_nl[17:0];
  assign nl_MultLoop_acc_214_nl = conv_s2s_24_25({(~ (data_rsci_idat[71:54])) , 6'b010000})
      + conv_s2s_22_25({(~ (data_rsci_idat[71:54])) , 4'b0001}) + conv_s2s_18_25(~
      (data_rsci_idat[71:54]));
  assign MultLoop_acc_214_nl = nl_MultLoop_acc_214_nl[24:0];
  assign nl_MultLoop_acc_57_nl = conv_s2s_25_27(MultLoop_acc_214_nl) + ({(data_rsci_idat[71:54])
      , 9'b001000000});
  assign MultLoop_acc_57_nl = nl_MultLoop_acc_57_nl[26:0];
  assign nl_MultLoop_acc_236_nl = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_110_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_109_nl))) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_358_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_57_nl)));
  assign MultLoop_acc_236_nl = nl_MultLoop_acc_236_nl[17:0];
  assign nl_MultLoop_acc_53_nl = (MultLoop_acc_54_itm_21_5[16:2]) + 15'b000000000101101;
  assign MultLoop_acc_53_nl = nl_MultLoop_acc_53_nl[14:0];
  assign nl_MultLoop_acc_227_nl = conv_s2s_17_18(MultLoop_acc_106_itm_22_6) + conv_s2s_17_18({(MultLoop_acc_53_nl)
      , (MultLoop_acc_54_itm_21_5[1:0])});
  assign MultLoop_acc_227_nl = nl_MultLoop_acc_227_nl[17:0];
  assign nl_MultLoop_acc_215_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[125:108]));
  assign MultLoop_acc_215_nl = nl_MultLoop_acc_215_nl[20:0];
  assign nl_MultLoop_acc_216_nl = ({(~ (data_rsci_idat[125:108])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_215_nl);
  assign MultLoop_acc_216_nl = nl_MultLoop_acc_216_nl[22:0];
  assign nl_MultLoop_acc_217_nl = ({(data_rsci_idat[125:108]) , 7'b0100000}) + conv_s2s_23_25(MultLoop_acc_216_nl);
  assign MultLoop_acc_217_nl = nl_MultLoop_acc_217_nl[24:0];
  assign nl_MultLoop_acc_343_nl = conv_s2u_16_19(readslicef_25_16_9((MultLoop_acc_217_nl)))
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_343_nl = nl_MultLoop_acc_343_nl[18:0];
  assign nl_MultLoop_acc_235_nl = (MultLoop_acc_227_nl) + (readslicef_19_18_1((MultLoop_acc_343_nl)));
  assign MultLoop_acc_235_nl = nl_MultLoop_acc_235_nl[17:0];
  assign nl_MultLoop_acc_344_nl =  -conv_s2s_9_10(data_rsci_idat[197:189]);
  assign MultLoop_acc_344_nl = nl_MultLoop_acc_344_nl[9:0];
  assign nl_MultLoop_acc_64_nl = conv_s2s_27_28({(~ (data_rsci_idat[197:180])) ,
      9'b000010000}) + conv_s2s_22_28({(~ (data_rsci_idat[197:180])) , 4'b0001})
      + conv_s2s_19_28({(MultLoop_acc_344_nl) , (~ (data_rsci_idat[188:180]))});
  assign MultLoop_acc_64_nl = nl_MultLoop_acc_64_nl[27:0];
  assign nl_MultLoop_acc_182_nl = conv_s2s_21_22({(~ (data_rsci_idat[89:72])) , 3'b001})
      + conv_s2s_18_22(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_182_nl = nl_MultLoop_acc_182_nl[21:0];
  assign nl_MultLoop_acc_58_nl = conv_s2s_22_23(MultLoop_acc_182_nl) + ({(data_rsci_idat[89:72])
      , 5'b01000});
  assign MultLoop_acc_58_nl = nl_MultLoop_acc_58_nl[22:0];
  assign nl_MultLoop_acc_183_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_15_18(data_rsci_idat[53:39]);
  assign MultLoop_acc_183_nl = nl_MultLoop_acc_183_nl[17:0];
  assign nl_MultLoop_acc_184_nl = conv_s2s_20_21({(~ (data_rsci_idat[53:36])) , 2'b01})
      + conv_s2s_18_21(MultLoop_acc_183_nl);
  assign MultLoop_acc_184_nl = nl_MultLoop_acc_184_nl[20:0];
  assign nl_MultLoop_acc_107_nl = conv_s2u_21_22(MultLoop_acc_184_nl) + ({(data_rsci_idat[53:36])
      , 4'b0100});
  assign MultLoop_acc_107_nl = nl_MultLoop_acc_107_nl[21:0];
  assign nl_MultLoop_acc_345_nl =  -conv_s2s_13_14(data_rsci_idat[359:347]);
  assign MultLoop_acc_345_nl = nl_MultLoop_acc_345_nl[13:0];
  assign nl_MultLoop_acc_177_nl = ({(data_rsci_idat[359:342]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_345_nl)
      , (~ (data_rsci_idat[346:342]))});
  assign MultLoop_acc_177_nl = nl_MultLoop_acc_177_nl[19:0];
  assign nl_MultLoop_acc_73_nl = conv_s2s_20_23(MultLoop_acc_177_nl) + ({(~ (data_rsci_idat[359:342]))
      , 5'b00000});
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[22:0];
  assign nl_MultLoop_acc_234_nl = (readslicef_28_18_10((MultLoop_acc_64_nl))) + conv_s2s_15_18(MultLoop_acc_72_itm_23_7[16:2])
      + conv_s2s_15_18(readslicef_23_15_8((MultLoop_acc_58_nl))) + conv_s2s_15_18(readslicef_22_15_7((MultLoop_acc_107_nl)))
      + conv_s2s_13_18(readslicef_23_13_10((MultLoop_acc_73_nl)));
  assign MultLoop_acc_234_nl = nl_MultLoop_acc_234_nl[17:0];
  assign nl_MultLoop_acc_351_nl =  -conv_s2s_9_10(data_rsci_idat[377:369]);
  assign MultLoop_acc_351_nl = nl_MultLoop_acc_351_nl[9:0];
  assign nl_MultLoop_acc_197_nl = ({(data_rsci_idat[377:360]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_351_nl)
      , (~ (data_rsci_idat[368:360]))});
  assign MultLoop_acc_197_nl = nl_MultLoop_acc_197_nl[20:0];
  assign nl_MultLoop_acc_198_nl = conv_s2s_23_24({(data_rsci_idat[377:360]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_197_nl);
  assign MultLoop_acc_198_nl = nl_MultLoop_acc_198_nl[23:0];
  assign nl_MultLoop_acc_352_nl = conv_s2u_18_19(data_rsci_idat[377:360]) + conv_s2u_17_19(readslicef_24_17_7((MultLoop_acc_198_nl)));
  assign MultLoop_acc_352_nl = nl_MultLoop_acc_352_nl[18:0];
  assign nl_MultLoop_acc_353_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_352_nl)))
      + (~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_353_nl = nl_MultLoop_acc_353_nl[17:0];
  assign nl_MultLoop_acc_354_nl =  -conv_s2s_11_12(data_rsci_idat[395:385]);
  assign MultLoop_acc_354_nl = nl_MultLoop_acc_354_nl[11:0];
  assign nl_MultLoop_acc_201_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_354_nl)
      , (~ (data_rsci_idat[384:378]))});
  assign MultLoop_acc_201_nl = nl_MultLoop_acc_201_nl[19:0];
  assign nl_MultLoop_acc_202_nl = conv_s2s_22_23({(data_rsci_idat[395:378]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_201_nl);
  assign MultLoop_acc_202_nl = nl_MultLoop_acc_202_nl[22:0];
  assign nl_MultLoop_acc_355_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_202_nl)))
      + (~ (data_rsci_idat[395:378]));
  assign MultLoop_acc_355_nl = nl_MultLoop_acc_355_nl[17:0];
  assign nl_MultLoop_acc_203_nl = (~ (data_rsci_idat[305:288])) + conv_s2s_14_18(data_rsci_idat[305:292]);
  assign MultLoop_acc_203_nl = nl_MultLoop_acc_203_nl[17:0];
  assign nl_MultLoop_acc_204_nl = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_203_nl);
  assign MultLoop_acc_204_nl = nl_MultLoop_acc_204_nl[19:0];
  assign nl_MultLoop_acc_111_nl = conv_s2u_20_23(MultLoop_acc_204_nl) + conv_s2u_22_23({(data_rsci_idat[305:288])
      , 4'b0000});
  assign MultLoop_acc_111_nl = nl_MultLoop_acc_111_nl[22:0];
  assign nl_MultLoop_acc_112_nl = conv_s2u_16_19(data_rsci_idat[323:308]) + conv_s2u_18_19(data_rsci_idat[323:306]);
  assign MultLoop_acc_112_nl = nl_MultLoop_acc_112_nl[18:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_238_nl) + (MultLoop_acc_236_nl) + (MultLoop_acc_235_nl)
      + (MultLoop_acc_234_nl) + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_353_nl)))
      + conv_s2s_17_18(readslicef_18_17_1((MultLoop_acc_355_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_111_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_112_nl)));

  function automatic [10:0] readslicef_18_11_7;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_18_11_7 = tmp[10:0];
  end
  endfunction


  function automatic [11:0] readslicef_18_12_6;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_18_12_6 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_18_13_5;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_18_13_5 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_18_14_4;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_18_14_4 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_18_15_3;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_18_15_3 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_18_16_2;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_18_16_2 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_18_17_1;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_18_17_1 = tmp[16:0];
  end
  endfunction


  function automatic [10:0] readslicef_19_11_8;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_19_11_8 = tmp[10:0];
  end
  endfunction


  function automatic [12:0] readslicef_19_13_6;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_19_13_6 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_19_14_5;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_19_14_5 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_19_15_4;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_19_15_4 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_19_16_3;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_19_16_3 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_19_17_2;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_19_17_2 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_19_18_1;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_19_18_1 = tmp[17:0];
  end
  endfunction


  function automatic [9:0] readslicef_20_10_10;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_20_10_10 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_20_11_9;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_20_11_9 = tmp[10:0];
  end
  endfunction


  function automatic [12:0] readslicef_20_13_7;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_20_13_7 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_20_14_6;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_20_14_6 = tmp[13:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_20_17_3;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_20_17_3 = tmp[16:0];
  end
  endfunction


  function automatic [12:0] readslicef_21_13_8;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_21_13_8 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_21_14_7;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_21_14_7 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_21_15_6;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_21_15_6 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_21_16_5;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_21_16_5 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_21_17_4;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_21_17_4 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_21_18_3;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_21_18_3 = tmp[17:0];
  end
  endfunction


  function automatic [13:0] readslicef_22_14_8;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_22_14_8 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_22_15_7;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_22_15_7 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_22_16_6;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_22_16_6 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_22_17_5;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_22_17_5 = tmp[16:0];
  end
  endfunction


  function automatic [12:0] readslicef_23_13_10;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_23_13_10 = tmp[12:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_23_16_7;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_23_16_7 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_23_17_6;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_23_17_6 = tmp[16:0];
  end
  endfunction


  function automatic [13:0] readslicef_24_14_10;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_24_14_10 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_24_15_9;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_24_15_9 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_24_16_8;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_24_16_8 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_24_17_7;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_24_17_7 = tmp[16:0];
  end
  endfunction


  function automatic [14:0] readslicef_25_15_10;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_25_15_10 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_25_16_9;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_25_16_9 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_25_17_8;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_25_17_8 = tmp[16:0];
  end
  endfunction


  function automatic [15:0] readslicef_26_16_10;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_26_16_10 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_26_17_9;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_26_17_9 = tmp[16:0];
  end
  endfunction


  function automatic [18:0] readslicef_26_19_7;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_26_19_7 = tmp[18:0];
  end
  endfunction


  function automatic [16:0] readslicef_27_17_10;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_27_17_10 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_28_18_10;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_28_18_10 = tmp[17:0];
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_10_18 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_18 = {{8{vector[9]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_13 = {{2{vector[10]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_13_17 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_17 = {{4{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_14_21 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_21 = {{7{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_15_21 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_21 = {{6{vector[14]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_15_22 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_22 = {{7{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_16_21 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_21 = {{5{vector[15]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_16_22 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_22 = {{6{vector[15]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_16_23 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_23 = {{7{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_17_21 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_21 = {{4{vector[16]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_17_23 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_23 = {{6{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_18_26 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_26 = {{8{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_19_25 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_25 = {{6{vector[18]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_19_26 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_26 = {{7{vector[18]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_19_28 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_28 = {{9{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_20_26 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_26 = {{6{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_21_25 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_25 = {{4{vector[20]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_21_26 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_26 = {{5{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_22_27 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_27 = {{5{vector[21]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_22_28 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_28 = {{6{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_23_26 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_26 = {{3{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_24_26 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_26 = {{2{vector[23]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_25_27 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_27 = {{2{vector[24]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2s_27_28 ;
    input [26:0]  vector ;
  begin
    conv_s2s_27_28 = {vector[26], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_9_19 ;
    input [8:0]  vector ;
  begin
    conv_s2u_9_19 = {{10{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_13_19 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_19 = {{6{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_21_25 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_25 = {{4{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_1_13 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_13 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_6_12 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_12 = {{6{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_10 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_11_13 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_13 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_1_11 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_layer3_t_layer4_t_config4
// ------------------------------------------------------------------


module nnet_dense_large_layer3_t_layer4_t_config4 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [107:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_layer3_t_layer4_t_config4_core nnet_dense_large_layer3_t_layer4_t_config4_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__relu_layer2_t_layer3_t_relu_config3__430e59af967157760564c6a2a3bbc91d13521_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 17:58:13 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3_core
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [431:0] data_rsci_idat;
  reg [16:0] res_rsci_d_412_396;
  reg [16:0] res_rsci_d_394_378;
  reg [16:0] res_rsci_d_376_360;
  reg [16:0] res_rsci_d_358_342;
  reg [16:0] res_rsci_d_340_324;
  reg [16:0] res_rsci_d_322_306;
  reg [16:0] res_rsci_d_304_288;
  reg [16:0] res_rsci_d_286_270;
  reg [16:0] res_rsci_d_268_252;
  reg [16:0] res_rsci_d_250_234;
  reg [16:0] res_rsci_d_232_216;
  reg [16:0] res_rsci_d_214_198;
  reg [16:0] res_rsci_d_196_180;
  reg [16:0] res_rsci_d_178_162;
  reg [16:0] res_rsci_d_160_144;
  reg [16:0] res_rsci_d_142_126;
  reg [16:0] res_rsci_d_124_108;
  reg [16:0] res_rsci_d_106_90;
  reg [16:0] res_rsci_d_88_72;
  reg [16:0] res_rsci_d_70_54;
  reg [16:0] res_rsci_d_52_36;
  reg [16:0] res_rsci_d_34_18;
  reg [16:0] res_rsci_d_16_0;
  reg [16:0] res_rsci_d_430_414;

  wire[18:0] for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[18:0] for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;
  wire[19:0] nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [431:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {1'b0 , res_rsci_d_430_414 , 1'b0 , res_rsci_d_412_396 ,
      1'b0 , res_rsci_d_394_378 , 1'b0 , res_rsci_d_376_360 , 1'b0 , res_rsci_d_358_342
      , 1'b0 , res_rsci_d_340_324 , 1'b0 , res_rsci_d_322_306 , 1'b0 , res_rsci_d_304_288
      , 1'b0 , res_rsci_d_286_270 , 1'b0 , res_rsci_d_268_252 , 1'b0 , res_rsci_d_250_234
      , 1'b0 , res_rsci_d_232_216 , 1'b0 , res_rsci_d_214_198 , 1'b0 , res_rsci_d_196_180
      , 1'b0 , res_rsci_d_178_162 , 1'b0 , res_rsci_d_160_144 , 1'b0 , res_rsci_d_142_126
      , 1'b0 , res_rsci_d_124_108 , 1'b0 , res_rsci_d_106_90 , 1'b0 , res_rsci_d_88_72
      , 1'b0 , res_rsci_d_70_54 , 1'b0 , res_rsci_d_52_36 , 1'b0 , res_rsci_d_34_18
      , 1'b0 , res_rsci_d_16_0};
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd432)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd432)) res_rsci (
      .d(nl_res_rsci_d[431:0]),
      .z(res_rsc_z)
    );
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_430_414 <= 17'b00000000000000000;
      res_rsci_d_16_0 <= 17'b00000000000000000;
      res_rsci_d_412_396 <= 17'b00000000000000000;
      res_rsci_d_34_18 <= 17'b00000000000000000;
      res_rsci_d_394_378 <= 17'b00000000000000000;
      res_rsci_d_52_36 <= 17'b00000000000000000;
      res_rsci_d_376_360 <= 17'b00000000000000000;
      res_rsci_d_70_54 <= 17'b00000000000000000;
      res_rsci_d_358_342 <= 17'b00000000000000000;
      res_rsci_d_88_72 <= 17'b00000000000000000;
      res_rsci_d_340_324 <= 17'b00000000000000000;
      res_rsci_d_106_90 <= 17'b00000000000000000;
      res_rsci_d_322_306 <= 17'b00000000000000000;
      res_rsci_d_124_108 <= 17'b00000000000000000;
      res_rsci_d_304_288 <= 17'b00000000000000000;
      res_rsci_d_142_126 <= 17'b00000000000000000;
      res_rsci_d_286_270 <= 17'b00000000000000000;
      res_rsci_d_160_144 <= 17'b00000000000000000;
      res_rsci_d_268_252 <= 17'b00000000000000000;
      res_rsci_d_178_162 <= 17'b00000000000000000;
      res_rsci_d_250_234 <= 17'b00000000000000000;
      res_rsci_d_196_180 <= 17'b00000000000000000;
      res_rsci_d_232_216 <= 17'b00000000000000000;
      res_rsci_d_214_198 <= 17'b00000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_430_414 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[430:414]),
          (readslicef_19_1_18((for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_16_0 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[16:0]),
          (readslicef_19_1_18((for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_412_396 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[412:396]),
          (readslicef_19_1_18((for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_34_18 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[34:18]),
          (readslicef_19_1_18((for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_394_378 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[394:378]),
          (readslicef_19_1_18((for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_52_36 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[52:36]),
          (readslicef_19_1_18((for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_376_360 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[376:360]),
          (readslicef_19_1_18((for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_70_54 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[70:54]),
          (readslicef_19_1_18((for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_358_342 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[358:342]),
          (readslicef_19_1_18((for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_88_72 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[88:72]),
          (readslicef_19_1_18((for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_340_324 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[340:324]),
          (readslicef_19_1_18((for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_106_90 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[106:90]),
          (readslicef_19_1_18((for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_322_306 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[322:306]),
          (readslicef_19_1_18((for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_124_108 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[124:108]),
          (readslicef_19_1_18((for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_304_288 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[304:288]),
          (readslicef_19_1_18((for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_142_126 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[142:126]),
          (readslicef_19_1_18((for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_286_270 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[286:270]),
          (readslicef_19_1_18((for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_160_144 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[160:144]),
          (readslicef_19_1_18((for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_268_252 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[268:252]),
          (readslicef_19_1_18((for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_178_162 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[178:162]),
          (readslicef_19_1_18((for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_250_234 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[250:234]),
          (readslicef_19_1_18((for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_196_180 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[196:180]),
          (readslicef_19_1_18((for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_232_216 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[232:216]),
          (readslicef_19_1_18((for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
      res_rsci_d_214_198 <= MUX_v_17_2_2(17'b00000000000000000, (data_rsci_idat[214:198]),
          (readslicef_19_1_18((for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl))));
    end
  end
  assign nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[431:414]);
  assign for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_24_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[17:0]);
  assign for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_1_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[413:396]);
  assign for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_23_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[35:18]);
  assign for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_2_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[395:378]);
  assign for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_22_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[53:36]);
  assign for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_3_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[377:360]);
  assign for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_21_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[71:54]);
  assign for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_4_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[359:342]);
  assign for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_20_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[89:72]);
  assign for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_5_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[341:324]);
  assign for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_19_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[107:90]);
  assign for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_6_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[323:306]);
  assign for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_18_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[125:108]);
  assign for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_7_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[305:288]);
  assign for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_17_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[143:126]);
  assign for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_8_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[287:270]);
  assign for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_16_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[161:144]);
  assign for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_9_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[269:252]);
  assign for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_15_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[179:162]);
  assign for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_10_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[251:234]);
  assign for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_14_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[197:180]);
  assign for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_11_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[233:216]);
  assign for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_13_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];
  assign nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl =  -conv_s2s_18_19(data_rsci_idat[215:198]);
  assign for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl = nl_for_12_operator_18_8_true_AC_TRN_AC_WRAP_acc_nl[18:0];

  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_19_1_18;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 18;
    readslicef_19_1_18 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_relu_layer2_t_layer3_t_relu_config3
// ------------------------------------------------------------------


module nnet_relu_layer2_t_layer3_t_relu_config3 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [431:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_relu_layer2_t_layer3_t_relu_config3_core nnet_relu_layer2_t_layer3_t_relu_config3_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ../td_ccore_solutions/nnet__dense_large_input_t_layer2_t_config2__1b7d9c734a4863f65ab961b20e6a3a0210dab8_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Fri Feb  7 18:09:23 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2_core
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2_core (
  data_rsc_dat, res_rsc_z, ccs_ccore_clk, ccs_ccore_srst, ccs_ccore_en
);
  input [863:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [863:0] data_rsci_idat;
  reg [17:0] res_rsci_d_431_414;
  wire [20:0] nl_res_rsci_d_431_414;
  reg [17:0] res_rsci_d_413_396;
  wire [20:0] nl_res_rsci_d_413_396;
  reg [17:0] res_rsci_d_395_378;
  wire [20:0] nl_res_rsci_d_395_378;
  reg [17:0] res_rsci_d_377_360;
  wire [21:0] nl_res_rsci_d_377_360;
  reg [17:0] res_rsci_d_359_342;
  wire [20:0] nl_res_rsci_d_359_342;
  reg [17:0] res_rsci_d_341_324;
  wire [20:0] nl_res_rsci_d_341_324;
  reg [17:0] res_rsci_d_323_306;
  wire [20:0] nl_res_rsci_d_323_306;
  reg [17:0] res_rsci_d_305_288;
  wire [20:0] nl_res_rsci_d_305_288;
  reg [17:0] res_rsci_d_287_270;
  wire [20:0] nl_res_rsci_d_287_270;
  reg [17:0] res_rsci_d_269_252;
  wire [20:0] nl_res_rsci_d_269_252;
  reg [17:0] res_rsci_d_251_234;
  wire [20:0] nl_res_rsci_d_251_234;
  reg [17:0] res_rsci_d_233_216;
  wire [20:0] nl_res_rsci_d_233_216;
  reg [17:0] res_rsci_d_215_198;
  wire [19:0] nl_res_rsci_d_215_198;
  reg [17:0] res_rsci_d_197_180;
  wire [20:0] nl_res_rsci_d_197_180;
  reg [17:0] res_rsci_d_179_162;
  wire [20:0] nl_res_rsci_d_179_162;
  reg [17:0] res_rsci_d_161_144;
  wire [20:0] nl_res_rsci_d_161_144;
  reg [17:0] res_rsci_d_143_126;
  wire [20:0] nl_res_rsci_d_143_126;
  reg [17:0] res_rsci_d_125_108;
  wire [20:0] nl_res_rsci_d_125_108;
  reg [17:0] res_rsci_d_107_90;
  wire [20:0] nl_res_rsci_d_107_90;
  reg [17:0] res_rsci_d_89_72;
  wire [20:0] nl_res_rsci_d_89_72;
  reg [17:0] res_rsci_d_71_54;
  wire [20:0] nl_res_rsci_d_71_54;
  reg [17:0] res_rsci_d_53_36;
  wire [20:0] nl_res_rsci_d_53_36;
  reg [17:0] res_rsci_d_35_18;
  wire [20:0] nl_res_rsci_d_35_18;
  reg [17:0] res_rsci_d_17_0;
  wire [19:0] nl_res_rsci_d_17_0;
  wire [18:0] MultLoop_acc_3283_cse;
  wire [19:0] nl_MultLoop_acc_3283_cse;
  wire [18:0] MultLoop_acc_3105_cse;
  wire [19:0] nl_MultLoop_acc_3105_cse;
  reg [17:0] MultLoop_acc_1588_itm_1;
  wire [20:0] nl_MultLoop_acc_1588_itm_1;
  reg [17:0] MultLoop_acc_1578_itm_1;
  wire [18:0] nl_MultLoop_acc_1578_itm_1;
  reg [15:0] MultLoop_acc_1562_itm_1;
  wire [17:0] nl_MultLoop_acc_1562_itm_1;
  reg [15:0] MultLoop_acc_1561_itm_1;
  wire [17:0] nl_MultLoop_acc_1561_itm_1;
  reg [16:0] MultLoop_acc_1576_itm_1;
  wire [18:0] nl_MultLoop_acc_1576_itm_1;
  reg [16:0] MultLoop_acc_1575_itm_1;
  wire [18:0] nl_MultLoop_acc_1575_itm_1;
  reg [17:0] MultLoop_acc_1585_itm_1;
  wire [20:0] nl_MultLoop_acc_1585_itm_1;
  reg [17:0] MultLoop_acc_1590_itm_1;
  wire [20:0] nl_MultLoop_acc_1590_itm_1;
  reg [17:0] MultLoop_acc_1582_itm_1;
  wire [19:0] nl_MultLoop_acc_1582_itm_1;
  reg [17:0] MultLoop_acc_1581_itm_1;
  wire [19:0] nl_MultLoop_acc_1581_itm_1;
  reg [17:0] MultLoop_acc_1683_itm_1;
  wire [19:0] nl_MultLoop_acc_1683_itm_1;
  reg [17:0] MultLoop_acc_1673_itm_1;
  wire [18:0] nl_MultLoop_acc_1673_itm_1;
  reg [15:0] MultLoop_acc_1659_itm_1;
  wire [17:0] nl_MultLoop_acc_1659_itm_1;
  reg [15:0] MultLoop_acc_1658_itm_1;
  wire [17:0] nl_MultLoop_acc_1658_itm_1;
  reg [16:0] MultLoop_acc_1671_itm_1;
  wire [19:0] nl_MultLoop_acc_1671_itm_1;
  reg [16:0] MultLoop_acc_1670_itm_1;
  wire [18:0] nl_MultLoop_acc_1670_itm_1;
  reg [16:0] MultLoop_acc_1669_itm_1;
  wire [18:0] nl_MultLoop_acc_1669_itm_1;
  reg [16:0] MultLoop_acc_1668_itm_1;
  wire [19:0] nl_MultLoop_acc_1668_itm_1;
  reg [17:0] MultLoop_acc_1685_itm_1;
  wire [20:0] nl_MultLoop_acc_1685_itm_1;
  reg [17:0] MultLoop_acc_1677_itm_1;
  wire [19:0] nl_MultLoop_acc_1677_itm_1;
  reg [17:0] MultLoop_acc_1676_itm_1;
  wire [19:0] nl_MultLoop_acc_1676_itm_1;
  reg [17:0] MultLoop_acc_1800_itm_1;
  wire [20:0] nl_MultLoop_acc_1800_itm_1;
  reg [15:0] MultLoop_acc_1772_itm_1;
  wire [18:0] nl_MultLoop_acc_1772_itm_1;
  reg [15:0] MultLoop_acc_1771_itm_1;
  wire [17:0] nl_MultLoop_acc_1771_itm_1;
  reg [16:0] MultLoop_acc_1783_itm_1;
  wire [19:0] nl_MultLoop_acc_1783_itm_1;
  reg [16:0] MultLoop_acc_1782_itm_1;
  wire [18:0] nl_MultLoop_acc_1782_itm_1;
  reg [16:0] MultLoop_acc_1781_itm_1;
  wire [18:0] nl_MultLoop_acc_1781_itm_1;
  reg [16:0] MultLoop_acc_1780_itm_1;
  wire [18:0] nl_MultLoop_acc_1780_itm_1;
  reg [16:0] MultLoop_acc_1779_itm_1;
  wire [17:0] nl_MultLoop_acc_1779_itm_1;
  reg [17:0] MultLoop_acc_1791_itm_1;
  wire [19:0] nl_MultLoop_acc_1791_itm_1;
  reg [17:0] MultLoop_acc_1797_itm_1;
  wire [20:0] nl_MultLoop_acc_1797_itm_1;
  reg [17:0] MultLoop_acc_1911_itm_1;
  wire [19:0] nl_MultLoop_acc_1911_itm_1;
  reg [17:0] MultLoop_acc_1910_itm_1;
  wire [19:0] nl_MultLoop_acc_1910_itm_1;
  reg [17:0] MultLoop_acc_1918_itm_1;
  wire [20:0] nl_MultLoop_acc_1918_itm_1;
  reg [17:0] MultLoop_acc_1917_itm_1;
  wire [19:0] nl_MultLoop_acc_1917_itm_1;
  reg [17:0] MultLoop_acc_1916_itm_1;
  wire [19:0] nl_MultLoop_acc_1916_itm_1;
  reg [15:0] MultLoop_acc_1889_itm_1;
  wire [17:0] nl_MultLoop_acc_1889_itm_1;
  reg [15:0] MultLoop_acc_1888_itm_1;
  wire [16:0] nl_MultLoop_acc_1888_itm_1;
  reg [16:0] MultLoop_acc_1902_itm_1;
  wire [18:0] nl_MultLoop_acc_1902_itm_1;
  reg [17:0] MultLoop_acc_1914_itm_1;
  wire [20:0] nl_MultLoop_acc_1914_itm_1;
  reg [17:0] MultLoop_acc_1920_itm_1;
  wire [20:0] nl_MultLoop_acc_1920_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1;
  reg [17:0] MultLoop_acc_2120_itm_1;
  wire [20:0] nl_MultLoop_acc_2120_itm_1;
  reg [17:0] MultLoop_acc_2119_itm_1;
  wire [20:0] nl_MultLoop_acc_2119_itm_1;
  reg [17:0] MultLoop_acc_2118_itm_1;
  wire [19:0] nl_MultLoop_acc_2118_itm_1;
  reg [15:0] MultLoop_acc_2091_itm_1;
  wire [17:0] nl_MultLoop_acc_2091_itm_1;
  reg [15:0] MultLoop_acc_2090_itm_1;
  wire [17:0] nl_MultLoop_acc_2090_itm_1;
  reg [16:0] MultLoop_acc_2105_itm_1;
  wire [18:0] nl_MultLoop_acc_2105_itm_1;
  reg [16:0] MultLoop_acc_2104_itm_1;
  wire [18:0] nl_MultLoop_acc_2104_itm_1;
  reg [16:0] MultLoop_acc_2103_itm_1;
  wire [17:0] nl_MultLoop_acc_2103_itm_1;
  reg [17:0] MultLoop_acc_2115_itm_1;
  wire [19:0] nl_MultLoop_acc_2115_itm_1;
  reg [17:0] MultLoop_acc_2121_itm_1;
  wire [20:0] nl_MultLoop_acc_2121_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_23_7_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1;
  wire [21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_26_10_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1;
  reg [17:0] MultLoop_acc_2470_itm_1;
  wire [20:0] nl_MultLoop_acc_2470_itm_1;
  reg [17:0] MultLoop_acc_2469_itm_1;
  wire [20:0] nl_MultLoop_acc_2469_itm_1;
  reg [16:0] MultLoop_acc_2458_itm_1;
  wire [19:0] nl_MultLoop_acc_2458_itm_1;
  reg [16:0] MultLoop_acc_2457_itm_1;
  wire [18:0] nl_MultLoop_acc_2457_itm_1;
  reg [15:0] MultLoop_acc_2438_itm_1;
  wire [16:0] nl_MultLoop_acc_2438_itm_1;
  reg [15:0] MultLoop_acc_2437_itm_1;
  wire [16:0] nl_MultLoop_acc_2437_itm_1;
  reg [16:0] MultLoop_acc_2455_itm_1;
  wire [19:0] nl_MultLoop_acc_2455_itm_1;
  reg [17:0] MultLoop_acc_2466_itm_1;
  wire [19:0] nl_MultLoop_acc_2466_itm_1;
  reg [16:0] MultLoop_acc_2452_itm_1;
  wire [17:0] nl_MultLoop_acc_2452_itm_1;
  reg [16:0] MultLoop_acc_2451_itm_1;
  wire [17:0] nl_MultLoop_acc_2451_itm_1;
  reg [17:0] MultLoop_acc_2464_itm_1;
  wire [19:0] nl_MultLoop_acc_2464_itm_1;
  reg [17:0] MultLoop_acc_2463_itm_1;
  wire [19:0] nl_MultLoop_acc_2463_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_25_10_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1;
  reg [17:0] MultLoop_acc_2658_itm_1;
  wire [20:0] nl_MultLoop_acc_2658_itm_1;
  reg [17:0] MultLoop_acc_2657_itm_1;
  wire [19:0] nl_MultLoop_acc_2657_itm_1;
  reg [17:0] MultLoop_acc_2656_itm_1;
  wire [19:0] nl_MultLoop_acc_2656_itm_1;
  reg [15:0] MultLoop_acc_2631_itm_1;
  wire [17:0] nl_MultLoop_acc_2631_itm_1;
  reg [15:0] MultLoop_acc_2630_itm_1;
  wire [16:0] nl_MultLoop_acc_2630_itm_1;
  reg [16:0] MultLoop_acc_2643_itm_1;
  wire [18:0] nl_MultLoop_acc_2643_itm_1;
  reg [16:0] MultLoop_acc_2642_itm_1;
  wire [18:0] nl_MultLoop_acc_2642_itm_1;
  reg [16:0] MultLoop_acc_2641_itm_1;
  wire [19:0] nl_MultLoop_acc_2641_itm_1;
  reg [17:0] MultLoop_acc_2653_itm_1;
  wire [19:0] nl_MultLoop_acc_2653_itm_1;
  reg [17:0] MultLoop_acc_2659_itm_1;
  wire [20:0] nl_MultLoop_acc_2659_itm_1;
  reg [17:0] MultLoop_acc_2773_itm_1;
  wire [19:0] nl_MultLoop_acc_2773_itm_1;
  reg [15:0] MultLoop_acc_2750_itm_1;
  wire [17:0] nl_MultLoop_acc_2750_itm_1;
  reg [15:0] MultLoop_acc_2749_itm_1;
  wire [17:0] nl_MultLoop_acc_2749_itm_1;
  reg [15:0] MultLoop_acc_2748_itm_1;
  wire [17:0] nl_MultLoop_acc_2748_itm_1;
  reg [15:0] MultLoop_acc_2747_itm_1;
  wire [16:0] nl_MultLoop_acc_2747_itm_1;
  reg [16:0] MultLoop_acc_2761_itm_1;
  wire [18:0] nl_MultLoop_acc_2761_itm_1;
  reg [16:0] MultLoop_acc_2760_itm_1;
  wire [18:0] nl_MultLoop_acc_2760_itm_1;
  reg [17:0] MultLoop_acc_2770_itm_1;
  wire [19:0] nl_MultLoop_acc_2770_itm_1;
  reg [17:0] MultLoop_acc_2775_itm_1;
  wire [20:0] nl_MultLoop_acc_2775_itm_1;
  reg [17:0] MultLoop_acc_2774_itm_1;
  wire [20:0] nl_MultLoop_acc_2774_itm_1;
  reg [17:0] MultLoop_acc_2888_itm_1;
  wire [19:0] nl_MultLoop_acc_2888_itm_1;
  reg [17:0] MultLoop_acc_2887_itm_1;
  wire [18:0] nl_MultLoop_acc_2887_itm_1;
  reg [17:0] MultLoop_acc_2886_itm_1;
  wire [18:0] nl_MultLoop_acc_2886_itm_1;
  reg [15:0] MultLoop_acc_2871_itm_1;
  wire [18:0] nl_MultLoop_acc_2871_itm_1;
  reg [15:0] MultLoop_acc_2870_itm_1;
  wire [16:0] nl_MultLoop_acc_2870_itm_1;
  reg [16:0] MultLoop_acc_2884_itm_1;
  wire [18:0] nl_MultLoop_acc_2884_itm_1;
  reg [16:0] MultLoop_acc_2883_itm_1;
  wire [18:0] nl_MultLoop_acc_2883_itm_1;
  reg [17:0] MultLoop_acc_2893_itm_1;
  wire [20:0] nl_MultLoop_acc_2893_itm_1;
  reg [17:0] MultLoop_acc_2898_itm_1;
  wire [20:0] nl_MultLoop_acc_2898_itm_1;
  reg [17:0] MultLoop_acc_2897_itm_1;
  wire [20:0] nl_MultLoop_acc_2897_itm_1;
  reg [17:0] MultLoop_acc_3018_itm_1;
  wire [19:0] nl_MultLoop_acc_3018_itm_1;
  reg [17:0] MultLoop_acc_3008_itm_1;
  wire [18:0] nl_MultLoop_acc_3008_itm_1;
  reg [14:0] MultLoop_acc_2984_itm_1;
  wire [15:0] nl_MultLoop_acc_2984_itm_1;
  reg [14:0] MultLoop_acc_2983_itm_1;
  wire [15:0] nl_MultLoop_acc_2983_itm_1;
  reg [15:0] MultLoop_acc_2993_itm_1;
  wire [17:0] nl_MultLoop_acc_2993_itm_1;
  reg [16:0] MultLoop_acc_3006_itm_1;
  wire [18:0] nl_MultLoop_acc_3006_itm_1;
  reg [16:0] MultLoop_acc_3005_itm_1;
  wire [18:0] nl_MultLoop_acc_3005_itm_1;
  reg [16:0] MultLoop_acc_3004_itm_1;
  wire [18:0] nl_MultLoop_acc_3004_itm_1;
  reg [16:0] MultLoop_acc_3003_itm_1;
  wire [18:0] nl_MultLoop_acc_3003_itm_1;
  reg [17:0] MultLoop_acc_3020_itm_1;
  wire [20:0] nl_MultLoop_acc_3020_itm_1;
  reg [17:0] MultLoop_acc_3012_itm_1;
  wire [19:0] nl_MultLoop_acc_3012_itm_1;
  reg [17:0] MultLoop_acc_3011_itm_1;
  wire [20:0] nl_MultLoop_acc_3011_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_acc_1215_22_6_itm_1;
  reg [14:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1;
  reg [14:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1;
  wire [15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1;
  wire [21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1;
  wire [20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1;
  reg [17:0] MultLoop_acc_3264_itm_1;
  wire [21:0] nl_MultLoop_acc_3264_itm_1;
  reg [17:0] MultLoop_acc_3258_itm_1;
  wire [19:0] nl_MultLoop_acc_3258_itm_1;
  reg [15:0] MultLoop_acc_3233_itm_1;
  wire [18:0] nl_MultLoop_acc_3233_itm_1;
  reg [15:0] MultLoop_acc_3232_itm_1;
  wire [16:0] nl_MultLoop_acc_3232_itm_1;
  reg [16:0] MultLoop_acc_3245_itm_1;
  wire [18:0] nl_MultLoop_acc_3245_itm_1;
  reg [17:0] MultLoop_acc_3256_itm_1;
  wire [20:0] nl_MultLoop_acc_3256_itm_1;
  reg [17:0] MultLoop_acc_3255_itm_1;
  wire [19:0] nl_MultLoop_acc_3255_itm_1;
  reg [17:0] MultLoop_acc_3254_itm_1;
  wire [19:0] nl_MultLoop_acc_3254_itm_1;
  reg [16:0] MultLoop_acc_3238_itm_1;
  wire [17:0] nl_MultLoop_acc_3238_itm_1;
  reg [16:0] MultLoop_acc_3237_itm_1;
  wire [17:0] nl_MultLoop_acc_3237_itm_1;
  reg [17:0] MultLoop_acc_3378_itm_1;
  wire [19:0] nl_MultLoop_acc_3378_itm_1;
  reg [17:0] MultLoop_acc_3368_itm_1;
  wire [20:0] nl_MultLoop_acc_3368_itm_1;
  reg [16:0] MultLoop_acc_3367_itm_1;
  wire [18:0] nl_MultLoop_acc_3367_itm_1;
  reg [16:0] MultLoop_acc_3366_itm_1;
  wire [18:0] nl_MultLoop_acc_3366_itm_1;
  reg [16:0] MultLoop_acc_3365_itm_1;
  wire [18:0] nl_MultLoop_acc_3365_itm_1;
  reg [17:0] MultLoop_acc_3375_itm_1;
  wire [19:0] nl_MultLoop_acc_3375_itm_1;
  reg [16:0] MultLoop_acc_3362_itm_1;
  wire [17:0] nl_MultLoop_acc_3362_itm_1;
  reg [16:0] MultLoop_acc_3361_itm_1;
  wire [17:0] nl_MultLoop_acc_3361_itm_1;
  reg [17:0] MultLoop_acc_3373_itm_1;
  wire [19:0] nl_MultLoop_acc_3373_itm_1;
  reg [17:0] MultLoop_acc_3379_itm_1;
  wire [20:0] nl_MultLoop_acc_3379_itm_1;
  reg [17:0] MultLoop_acc_3495_itm_1;
  wire [20:0] nl_MultLoop_acc_3495_itm_1;
  reg [17:0] MultLoop_acc_3494_itm_1;
  wire [19:0] nl_MultLoop_acc_3494_itm_1;
  reg [15:0] MultLoop_acc_3469_itm_1;
  wire [17:0] nl_MultLoop_acc_3469_itm_1;
  reg [15:0] MultLoop_acc_3468_itm_1;
  wire [16:0] nl_MultLoop_acc_3468_itm_1;
  reg [16:0] MultLoop_acc_3482_itm_1;
  wire [18:0] nl_MultLoop_acc_3482_itm_1;
  reg [16:0] MultLoop_acc_3481_itm_1;
  wire [18:0] nl_MultLoop_acc_3481_itm_1;
  reg [16:0] MultLoop_acc_3480_itm_1;
  wire [18:0] nl_MultLoop_acc_3480_itm_1;
  reg [16:0] MultLoop_acc_3479_itm_1;
  wire [18:0] nl_MultLoop_acc_3479_itm_1;
  reg [16:0] MultLoop_acc_3478_itm_1;
  wire [17:0] nl_MultLoop_acc_3478_itm_1;
  reg [17:0] MultLoop_acc_3490_itm_1;
  wire [19:0] nl_MultLoop_acc_3490_itm_1;
  reg [17:0] MultLoop_acc_3496_itm_1;
  wire [20:0] nl_MultLoop_acc_3496_itm_1;
  reg [17:0] MultLoop_acc_3614_itm_1;
  wire [20:0] nl_MultLoop_acc_3614_itm_1;
  reg [17:0] MultLoop_acc_3598_itm_1;
  wire [18:0] nl_MultLoop_acc_3598_itm_1;
  reg [15:0] MultLoop_acc_3584_itm_1;
  wire [17:0] nl_MultLoop_acc_3584_itm_1;
  reg [15:0] MultLoop_acc_3583_itm_1;
  wire [17:0] nl_MultLoop_acc_3583_itm_1;
  reg [16:0] MultLoop_acc_3596_itm_1;
  wire [19:0] nl_MultLoop_acc_3596_itm_1;
  reg [16:0] MultLoop_acc_3595_itm_1;
  wire [18:0] nl_MultLoop_acc_3595_itm_1;
  reg [16:0] MultLoop_acc_3594_itm_1;
  wire [18:0] nl_MultLoop_acc_3594_itm_1;
  reg [16:0] MultLoop_acc_3593_itm_1;
  wire [17:0] nl_MultLoop_acc_3593_itm_1;
  reg [17:0] MultLoop_acc_3605_itm_1;
  wire [19:0] nl_MultLoop_acc_3605_itm_1;
  reg [17:0] MultLoop_acc_3611_itm_1;
  wire [20:0] nl_MultLoop_acc_3611_itm_1;
  reg [17:0] MultLoop_acc_3720_itm_1;
  wire [19:0] nl_MultLoop_acc_3720_itm_1;
  reg [17:0] MultLoop_acc_3719_itm_1;
  wire [18:0] nl_MultLoop_acc_3719_itm_1;
  reg [17:0] MultLoop_acc_3718_itm_1;
  wire [18:0] nl_MultLoop_acc_3718_itm_1;
  reg [16:0] MultLoop_acc_3716_itm_1;
  wire [19:0] nl_MultLoop_acc_3716_itm_1;
  reg [16:0] MultLoop_acc_3715_itm_1;
  wire [18:0] nl_MultLoop_acc_3715_itm_1;
  reg [17:0] MultLoop_acc_3725_itm_1;
  wire [20:0] nl_MultLoop_acc_3725_itm_1;
  reg [17:0] MultLoop_acc_3724_itm_1;
  wire [19:0] nl_MultLoop_acc_3724_itm_1;
  reg [16:0] MultLoop_acc_3710_itm_1;
  wire [17:0] nl_MultLoop_acc_3710_itm_1;
  reg [16:0] MultLoop_acc_3709_itm_1;
  wire [17:0] nl_MultLoop_acc_3709_itm_1;
  reg [17:0] MultLoop_acc_3722_itm_1;
  wire [19:0] nl_MultLoop_acc_3722_itm_1;
  reg [16:0] MultLoop_acc_3706_itm_1;
  wire [17:0] nl_MultLoop_acc_3706_itm_1;
  reg [16:0] MultLoop_acc_3705_itm_1;
  wire [17:0] nl_MultLoop_acc_3705_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1;
  reg [15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1;
  wire [16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1;
  wire [18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1;
  reg [17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1;
  wire [21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1;
  reg [17:0] MultLoop_acc_3913_itm_1;
  wire [21:0] nl_MultLoop_acc_3913_itm_1;
  reg [15:0] MultLoop_acc_3881_itm_1;
  wire [17:0] nl_MultLoop_acc_3881_itm_1;
  reg [15:0] MultLoop_acc_3880_itm_1;
  wire [16:0] nl_MultLoop_acc_3880_itm_1;
  reg [16:0] MultLoop_acc_3896_itm_1;
  wire [18:0] nl_MultLoop_acc_3896_itm_1;
  reg [16:0] MultLoop_acc_3895_itm_1;
  wire [18:0] nl_MultLoop_acc_3895_itm_1;
  reg [16:0] MultLoop_acc_3894_itm_1;
  wire [18:0] nl_MultLoop_acc_3894_itm_1;
  reg [17:0] MultLoop_acc_3911_itm_1;
  wire [20:0] nl_MultLoop_acc_3911_itm_1;
  reg [17:0] MultLoop_acc_3910_itm_1;
  wire [20:0] nl_MultLoop_acc_3910_itm_1;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0;
  wire [19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0;
  reg [16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0;
  wire [17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0;
  reg [16:0] MultLoop_acc_3717_itm_1_16_0;
  wire [18:0] nl_MultLoop_acc_3717_itm_1_16_0;
  wire [17:0] MultLoop_acc_2133_cse_1;
  wire [18:0] nl_MultLoop_acc_2133_cse_1;
  wire [17:0] MultLoop_acc_2535_cse_1;
  wire [18:0] nl_MultLoop_acc_2535_cse_1;
  wire [10:0] MultLoop_acc_4229_cse_1;
  wire [11:0] nl_MultLoop_acc_4229_cse_1;
  wire [18:0] MultLoop_acc_2591_cse_1;
  wire [19:0] nl_MultLoop_acc_2591_cse_1;
  wire [21:0] MultLoop_acc_3099_cse_1;
  wire [22:0] nl_MultLoop_acc_3099_cse_1;
  wire [17:0] MultLoop_acc_1946_cse_1;
  wire [18:0] nl_MultLoop_acc_1946_cse_1;
  wire [12:0] MultLoop_acc_3961_cse_1;
  wire [13:0] nl_MultLoop_acc_3961_cse_1;
  wire [12:0] Result_acc_192_cse_1;
  wire [13:0] nl_Result_acc_192_cse_1;
  wire [18:0] MultLoop_acc_3661_cse_1;
  wire [19:0] nl_MultLoop_acc_3661_cse_1;
  wire [20:0] MultLoop_acc_2387_cse_1;
  wire [21:0] nl_MultLoop_acc_2387_cse_1;
  wire [18:0] MultLoop_acc_2220_cse_1;
  wire [19:0] nl_MultLoop_acc_2220_cse_1;
  wire [20:0] MultLoop_acc_1722_cse_1;
  wire [21:0] nl_MultLoop_acc_1722_cse_1;
  wire [10:0] MultLoop_acc_4212_cse_1;
  wire [11:0] nl_MultLoop_acc_4212_cse_1;
  wire [18:0] MultLoop_acc_1611_cse_1;
  wire [19:0] nl_MultLoop_acc_1611_cse_1;
  wire [10:0] MultLoop_acc_4167_cse_1;
  wire [11:0] nl_MultLoop_acc_4167_cse_1;
  wire [18:0] MultLoop_acc_2584_cse_1;
  wire [19:0] nl_MultLoop_acc_2584_cse_1;
  wire [19:0] MultLoop_acc_3636_cse_1;
  wire [20:0] nl_MultLoop_acc_3636_cse_1;
  wire [18:0] MultLoop_acc_2057_cse_1;
  wire [19:0] nl_MultLoop_acc_2057_cse_1;
  wire [19:0] MultLoop_acc_3182_cse_1;
  wire [20:0] nl_MultLoop_acc_3182_cse_1;
  wire [17:0] MultLoop_acc_2307_cse_1;
  wire [18:0] nl_MultLoop_acc_2307_cse_1;
  wire [17:0] MultLoop_acc_2685_cse_1;
  wire [18:0] nl_MultLoop_acc_2685_cse_1;
  wire [20:0] MultLoop_acc_1949_cse_1;
  wire [21:0] nl_MultLoop_acc_1949_cse_1;
  wire [10:0] Result_acc_214_cse_1;
  wire [11:0] nl_Result_acc_214_cse_1;
  wire [11:0] MultLoop_acc_4083_cse_1;
  wire [12:0] nl_MultLoop_acc_4083_cse_1;
  wire [12:0] MultLoop_acc_3946_cse_1;
  wire [13:0] nl_MultLoop_acc_3946_cse_1;
  wire [10:0] Result_acc_178_cse_1;
  wire [11:0] nl_Result_acc_178_cse_1;
  wire [11:0] MultLoop_acc_4233_cse_1;
  wire [12:0] nl_MultLoop_acc_4233_cse_1;
  wire [20:0] MultLoop_acc_1618_cse_1;
  wire [21:0] nl_MultLoop_acc_1618_cse_1;
  wire [18:0] MultLoop_acc_2424_cse_1;
  wire [19:0] nl_MultLoop_acc_2424_cse_1;
  wire [17:0] MultLoop_acc_2079_cse_1;
  wire [18:0] nl_MultLoop_acc_2079_cse_1;
  wire [17:0] MultLoop_acc_2568_cse_1;
  wire [18:0] nl_MultLoop_acc_2568_cse_1;
  wire [19:0] MultLoop_acc_2520_cse_1;
  wire [20:0] nl_MultLoop_acc_2520_cse_1;
  wire [20:0] MultLoop_acc_1720_cse_1;
  wire [21:0] nl_MultLoop_acc_1720_cse_1;
  wire [17:0] MultLoop_acc_2375_cse_1;
  wire [18:0] nl_MultLoop_acc_2375_cse_1;
  wire [17:0] MultLoop_acc_3063_cse_1;
  wire [18:0] nl_MultLoop_acc_3063_cse_1;
  wire [18:0] MultLoop_acc_3187_cse_1;
  wire [19:0] nl_MultLoop_acc_3187_cse_1;
  wire [10:0] MultLoop_acc_3974_cse_1;
  wire [11:0] nl_MultLoop_acc_3974_cse_1;
  wire [20:0] MultLoop_acc_2390_cse_1;
  wire [21:0] nl_MultLoop_acc_2390_cse_1;
  wire [12:0] Result_acc_190_cse_1;
  wire [13:0] nl_Result_acc_190_cse_1;
  wire [18:0] MultLoop_acc_1822_cse_1;
  wire [19:0] nl_MultLoop_acc_1822_cse_1;
  wire [10:0] MultLoop_acc_4122_cse_1;
  wire [11:0] nl_MultLoop_acc_4122_cse_1;
  wire [11:0] MultLoop_acc_3941_cse_1;
  wire [12:0] nl_MultLoop_acc_3941_cse_1;
  wire [10:0] MultLoop_acc_4011_cse_1;
  wire [11:0] nl_MultLoop_acc_4011_cse_1;
  wire [20:0] MultLoop_acc_2385_cse_1;
  wire [21:0] nl_MultLoop_acc_2385_cse_1;
  wire [17:0] Result_acc_143_cse_1;
  wire [18:0] nl_Result_acc_143_cse_1;
  wire [18:0] MultLoop_acc_2566_cse_1;
  wire [19:0] nl_MultLoop_acc_2566_cse_1;
  wire [20:0] MultLoop_acc_1743_cse_1;
  wire [21:0] nl_MultLoop_acc_1743_cse_1;
  wire [18:0] Result_acc_111_cse_1;
  wire [19:0] nl_Result_acc_111_cse_1;
  wire [17:0] MultLoop_acc_2574_cse_1;
  wire [18:0] nl_MultLoop_acc_2574_cse_1;
  wire [20:0] MultLoop_acc_1480_cse_1;
  wire [21:0] nl_MultLoop_acc_1480_cse_1;
  wire [17:0] Result_acc_152_cse_1;
  wire [18:0] nl_Result_acc_152_cse_1;
  wire [18:0] MultLoop_acc_2073_cse_1;
  wire [19:0] nl_MultLoop_acc_2073_cse_1;
  wire [18:0] MultLoop_acc_2522_cse_1;
  wire [19:0] nl_MultLoop_acc_2522_cse_1;
  wire [18:0] MultLoop_acc_2967_cse_1;
  wire [19:0] nl_MultLoop_acc_2967_cse_1;
  wire [18:0] MultLoop_acc_2412_cse_1;
  wire [19:0] nl_MultLoop_acc_2412_cse_1;
  wire [20:0] MultLoop_acc_1485_cse_1;
  wire [21:0] nl_MultLoop_acc_1485_cse_1;
  wire [19:0] MultLoop_acc_788_cse_1;
  wire [20:0] nl_MultLoop_acc_788_cse_1;
  wire [19:0] MultLoop_acc_2923_cse_1;
  wire [20:0] nl_MultLoop_acc_2923_cse_1;
  wire [11:0] MultLoop_acc_4162_cse_1;
  wire [12:0] nl_MultLoop_acc_4162_cse_1;
  wire [17:0] MultLoop_acc_1636_cse_1;
  wire [18:0] nl_MultLoop_acc_1636_cse_1;
  wire [10:0] MultLoop_acc_4146_cse_1;
  wire [11:0] nl_MultLoop_acc_4146_cse_1;
  wire [18:0] MultLoop_acc_1962_cse_1;
  wire [19:0] nl_MultLoop_acc_1962_cse_1;
  wire [10:0] Result_acc_206_cse_1;
  wire [11:0] nl_Result_acc_206_cse_1;
  wire [18:0] MultLoop_acc_1708_cse_1;
  wire [19:0] nl_MultLoop_acc_1708_cse_1;
  wire [17:0] MultLoop_acc_2604_cse_1;
  wire [18:0] nl_MultLoop_acc_2604_cse_1;
  wire [13:0] MultLoop_acc_4032_cse_1;
  wire [14:0] nl_MultLoop_acc_4032_cse_1;
  wire [21:0] MultLoop_acc_2592_cse_1;
  wire [22:0] nl_MultLoop_acc_2592_cse_1;
  wire [10:0] MultLoop_acc_3976_cse_1;
  wire [11:0] nl_MultLoop_acc_3976_cse_1;
  wire [20:0] Result_acc_129_cse_1;
  wire [21:0] nl_Result_acc_129_cse_1;
  wire [13:0] MultLoop_acc_4094_cse_1;
  wire [14:0] nl_MultLoop_acc_4094_cse_1;
  wire [18:0] MultLoop_acc_1503_cse_1;
  wire [19:0] nl_MultLoop_acc_1503_cse_1;
  wire [10:0] MultLoop_acc_4186_cse_1;
  wire [11:0] nl_MultLoop_acc_4186_cse_1;
  wire [21:0] MultLoop_acc_2781_cse_1;
  wire [22:0] nl_MultLoop_acc_2781_cse_1;
  wire [19:0] MultLoop_acc_1940_cse_1;
  wire [20:0] nl_MultLoop_acc_1940_cse_1;
  wire [18:0] MultLoop_acc_2337_cse_1;
  wire [19:0] nl_MultLoop_acc_2337_cse_1;
  wire [18:0] MultLoop_acc_2525_cse_1;
  wire [19:0] nl_MultLoop_acc_2525_cse_1;
  wire [11:0] Result_acc_216_cse_1;
  wire [12:0] nl_Result_acc_216_cse_1;
  wire [10:0] MultLoop_acc_4015_cse_1;
  wire [11:0] nl_MultLoop_acc_4015_cse_1;
  wire [12:0] MultLoop_acc_4076_cse_1;
  wire [13:0] nl_MultLoop_acc_4076_cse_1;
  wire [10:0] MultLoop_acc_4191_cse_1;
  wire [11:0] nl_MultLoop_acc_4191_cse_1;
  wire [10:0] MultLoop_acc_4153_cse_1;
  wire [11:0] nl_MultLoop_acc_4153_cse_1;
  wire [12:0] MultLoop_acc_4021_cse_1;
  wire [13:0] nl_MultLoop_acc_4021_cse_1;
  wire [18:0] MultLoop_acc_2500_cse_1;
  wire [19:0] nl_MultLoop_acc_2500_cse_1;
  wire [21:0] MultLoop_acc_1603_cse_1;
  wire [22:0] nl_MultLoop_acc_1603_cse_1;
  wire [18:0] Result_acc_127_cse_1;
  wire [19:0] nl_Result_acc_127_cse_1;
  wire [11:0] MultLoop_acc_3955_cse_1;
  wire [12:0] nl_MultLoop_acc_3955_cse_1;
  wire [10:0] MultLoop_acc_4084_cse_1;
  wire [11:0] nl_MultLoop_acc_4084_cse_1;
  wire [18:0] MultLoop_acc_1741_cse_1;
  wire [19:0] nl_MultLoop_acc_1741_cse_1;
  wire [18:0] MultLoop_acc_1531_cse_1;
  wire [19:0] nl_MultLoop_acc_1531_cse_1;
  wire [11:0] Result_acc_187_cse_1;
  wire [12:0] nl_Result_acc_187_cse_1;
  wire [17:0] MultLoop_acc_2403_cse_1;
  wire [18:0] nl_MultLoop_acc_2403_cse_1;
  wire [20:0] MultLoop_acc_2030_cse_1;
  wire [21:0] nl_MultLoop_acc_2030_cse_1;
  wire [12:0] MultLoop_acc_3916_cse_1;
  wire [13:0] nl_MultLoop_acc_3916_cse_1;
  wire [10:0] MultLoop_acc_4150_cse_1;
  wire [11:0] nl_MultLoop_acc_4150_cse_1;
  wire [10:0] MultLoop_acc_4030_cse_1;
  wire [11:0] nl_MultLoop_acc_4030_cse_1;
  wire [10:0] MultLoop_acc_3987_cse_1;
  wire [11:0] nl_MultLoop_acc_3987_cse_1;
  wire [17:0] MultLoop_acc_2259_cse_1;
  wire [18:0] nl_MultLoop_acc_2259_cse_1;
  wire [11:0] MultLoop_acc_3925_cse_1;
  wire [12:0] nl_MultLoop_acc_3925_cse_1;
  wire [18:0] Result_acc_163_cse_1;
  wire [19:0] nl_Result_acc_163_cse_1;
  wire [17:0] MultLoop_acc_2035_cse_1;
  wire [18:0] nl_MultLoop_acc_2035_cse_1;
  wire [11:0] Result_acc_183_cse_1;
  wire [12:0] nl_Result_acc_183_cse_1;
  wire [12:0] MultLoop_acc_4075_cse_1;
  wire [13:0] nl_MultLoop_acc_4075_cse_1;
  wire [19:0] MultLoop_acc_1043_cse_1;
  wire [20:0] nl_MultLoop_acc_1043_cse_1;
  wire [10:0] MultLoop_acc_3989_cse_1;
  wire [11:0] nl_MultLoop_acc_3989_cse_1;
  wire [20:0] MultLoop_acc_1735_cse_1;
  wire [21:0] nl_MultLoop_acc_1735_cse_1;
  wire [20:0] MultLoop_acc_1957_cse_1;
  wire [21:0] nl_MultLoop_acc_1957_cse_1;
  wire [19:0] MultLoop_acc_1723_cse_1;
  wire [20:0] nl_MultLoop_acc_1723_cse_1;
  wire [18:0] MultLoop_acc_1727_cse_1;
  wire [19:0] nl_MultLoop_acc_1727_cse_1;
  wire [11:0] MultLoop_acc_4036_cse_1;
  wire [12:0] nl_MultLoop_acc_4036_cse_1;
  wire [17:0] MultLoop_acc_1626_cse_1;
  wire [18:0] nl_MultLoop_acc_1626_cse_1;
  wire [17:0] MultLoop_acc_1844_cse_1;
  wire [18:0] nl_MultLoop_acc_1844_cse_1;
  wire [20:0] MultLoop_acc_1702_cse_1;
  wire [21:0] nl_MultLoop_acc_1702_cse_1;
  wire [20:0] MultLoop_acc_1520_cse_1;
  wire [21:0] nl_MultLoop_acc_1520_cse_1;
  wire [20:0] MultLoop_acc_4688;
  wire [21:0] nl_MultLoop_acc_4688;
  wire [22:0] MultLoop_acc_4690;
  wire [23:0] nl_MultLoop_acc_4690;
  wire [19:0] MultLoop_acc_4692;
  wire [20:0] nl_MultLoop_acc_4692;
  wire [17:0] MultLoop_asn_1479;
  wire [18:0] nl_MultLoop_asn_1479;
  wire [13:0] MultLoop_MultLoop_conc_674_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_674_18_5;
  wire [12:0] MultLoop_MultLoop_conc_676_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_676_18_6;
  wire [11:0] MultLoop_MultLoop_conc_678_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_678_18_7;
  wire [10:0] MultLoop_MultLoop_conc_680_16_6;
  wire [11:0] nl_MultLoop_MultLoop_conc_680_16_6;
  wire [10:0] MultLoop_MultLoop_conc_682_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_682_18_8;
  wire [12:0] MultLoop_MultLoop_conc_686_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_686_18_6;
  wire [11:0] MultLoop_MultLoop_conc_688_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_688_18_7;
  wire [12:0] MultLoop_MultLoop_conc_690_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_690_18_6;
  wire [11:0] MultLoop_MultLoop_conc_692_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_692_18_7;
  wire [12:0] MultLoop_MultLoop_conc_694_15_3;
  wire [13:0] nl_MultLoop_MultLoop_conc_694_15_3;
  wire [11:0] MultLoop_MultLoop_conc_696_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_696_18_7;
  wire [11:0] MultLoop_MultLoop_conc_698_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_698_18_7;
  wire [11:0] MultLoop_MultLoop_conc_700_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_700_18_7;
  wire [12:0] MultLoop_MultLoop_conc_702_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_702_18_6;
  wire [12:0] MultLoop_MultLoop_conc_704_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_704_18_6;
  wire [12:0] MultLoop_MultLoop_conc_706_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_706_16_4;
  wire [12:0] MultLoop_MultLoop_conc_708_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_708_18_6;
  wire [13:0] MultLoop_MultLoop_conc_714_15_2;
  wire [14:0] nl_MultLoop_MultLoop_conc_714_15_2;
  wire [11:0] MultLoop_MultLoop_conc_716_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_716_18_7;
  wire [10:0] MultLoop_MultLoop_conc_718_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_718_18_8;
  wire [11:0] MultLoop_MultLoop_conc_720_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_720_18_7;
  wire [10:0] MultLoop_MultLoop_conc_722_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_722_18_8;
  wire [12:0] MultLoop_MultLoop_conc_724_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_724_18_6;
  wire [11:0] MultLoop_MultLoop_conc_726_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_726_18_7;
  wire [10:0] MultLoop_MultLoop_conc_728_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_728_18_8;
  wire [11:0] MultLoop_MultLoop_conc_730_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_730_18_7;
  wire [12:0] MultLoop_MultLoop_conc_732_14_2;
  wire [13:0] nl_MultLoop_MultLoop_conc_732_14_2;
  wire [11:0] MultLoop_MultLoop_conc_734_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_734_18_7;
  wire [11:0] MultLoop_MultLoop_conc_736_16_5;
  wire [12:0] nl_MultLoop_MultLoop_conc_736_16_5;
  wire [14:0] MultLoop_MultLoop_conc_738_18_4;
  wire [15:0] nl_MultLoop_MultLoop_conc_738_18_4;
  wire [12:0] MultLoop_MultLoop_conc_740_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_740_16_4;
  wire [12:0] MultLoop_MultLoop_conc_742_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_742_18_6;
  wire [10:0] MultLoop_MultLoop_conc_746_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_746_18_8;
  wire [11:0] MultLoop_MultLoop_conc_750_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_750_18_7;
  wire [12:0] MultLoop_MultLoop_conc_752_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_752_18_6;
  wire [12:0] MultLoop_MultLoop_conc_754_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_754_18_6;
  wire [10:0] MultLoop_MultLoop_conc_756_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_756_18_8;
  wire [12:0] MultLoop_MultLoop_conc_758_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_758_18_6;
  wire [13:0] MultLoop_MultLoop_conc_760_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_760_18_5;
  wire [11:0] MultLoop_MultLoop_conc_766_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_766_18_7;
  wire [13:0] MultLoop_MultLoop_conc_768_15_2;
  wire [14:0] nl_MultLoop_MultLoop_conc_768_15_2;
  wire [10:0] MultLoop_MultLoop_conc_770_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_770_18_8;
  wire [14:0] MultLoop_MultLoop_conc_772_16_2;
  wire [15:0] nl_MultLoop_MultLoop_conc_772_16_2;
  wire [12:0] MultLoop_MultLoop_conc_774_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_774_16_4;
  wire [11:0] MultLoop_MultLoop_conc_776_15_4;
  wire [12:0] nl_MultLoop_MultLoop_conc_776_15_4;
  wire [10:0] MultLoop_MultLoop_conc_778_16_6;
  wire [11:0] nl_MultLoop_MultLoop_conc_778_16_6;
  wire [10:0] MultLoop_MultLoop_conc_780_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_780_18_8;
  wire [10:0] MultLoop_MultLoop_conc_782_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_782_18_8;
  wire [10:0] MultLoop_MultLoop_conc_784_16_6;
  wire [11:0] nl_MultLoop_MultLoop_conc_784_16_6;
  wire [11:0] MultLoop_MultLoop_conc_786_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_786_18_7;
  wire [13:0] MultLoop_MultLoop_conc_788_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_788_18_5;
  wire [12:0] MultLoop_MultLoop_conc_790_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_790_16_4;
  wire [12:0] MultLoop_MultLoop_conc_792_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_792_18_6;
  wire [11:0] MultLoop_MultLoop_conc_794_16_5;
  wire [12:0] nl_MultLoop_MultLoop_conc_794_16_5;
  wire [10:0] MultLoop_MultLoop_conc_796_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_796_18_8;
  wire [12:0] MultLoop_MultLoop_conc_798_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_798_16_4;
  wire [11:0] MultLoop_MultLoop_conc_800_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_800_18_7;
  wire [10:0] MultLoop_MultLoop_conc_802_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_802_18_8;
  wire [11:0] MultLoop_MultLoop_conc_804_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_804_18_7;
  wire [13:0] MultLoop_MultLoop_conc_806_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_806_18_5;
  wire [13:0] MultLoop_MultLoop_conc_810_15_2;
  wire [14:0] nl_MultLoop_MultLoop_conc_810_15_2;
  wire [10:0] MultLoop_MultLoop_conc_814_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_814_18_8;
  wire [11:0] MultLoop_MultLoop_conc_816_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_816_18_7;
  wire [11:0] MultLoop_MultLoop_conc_818_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_818_18_7;
  wire [10:0] MultLoop_MultLoop_conc_820_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_820_18_8;
  wire [11:0] MultLoop_MultLoop_conc_822_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_822_18_7;
  wire [12:0] MultLoop_MultLoop_conc_824_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_824_18_6;
  wire [13:0] MultLoop_MultLoop_conc_826_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_826_18_5;
  wire [11:0] MultLoop_MultLoop_conc_828_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_828_18_7;
  wire [12:0] MultLoop_MultLoop_conc_830_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_830_18_6;
  wire [11:0] MultLoop_MultLoop_conc_832_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_832_18_7;
  wire [13:0] MultLoop_MultLoop_conc_834_18_5;
  wire [14:0] nl_MultLoop_MultLoop_conc_834_18_5;
  wire [10:0] MultLoop_MultLoop_conc_836_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_836_18_8;
  wire [14:0] MultLoop_MultLoop_conc_838_18_4;
  wire [15:0] nl_MultLoop_MultLoop_conc_838_18_4;
  wire [11:0] MultLoop_MultLoop_conc_840_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_840_18_7;
  wire [12:0] MultLoop_MultLoop_conc_842_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_842_18_6;
  wire [11:0] MultLoop_MultLoop_conc_844_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_844_18_7;
  wire [10:0] MultLoop_MultLoop_conc_846_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_846_18_8;
  wire [11:0] MultLoop_MultLoop_conc_848_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_848_18_7;
  wire [12:0] MultLoop_MultLoop_conc_850_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_850_18_6;
  wire [12:0] MultLoop_MultLoop_conc_852_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_852_18_6;
  wire [10:0] MultLoop_MultLoop_conc_854_18_8;
  wire [11:0] nl_MultLoop_MultLoop_conc_854_18_8;
  wire [11:0] MultLoop_MultLoop_conc_856_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_856_18_7;
  wire [11:0] MultLoop_MultLoop_conc_858_18_7;
  wire [12:0] nl_MultLoop_MultLoop_conc_858_18_7;
  wire [12:0] MultLoop_MultLoop_conc_860_16_4;
  wire [13:0] nl_MultLoop_MultLoop_conc_860_16_4;
  wire [12:0] MultLoop_MultLoop_conc_862_18_6;
  wire [13:0] nl_MultLoop_MultLoop_conc_862_18_6;
  wire [11:0] MultLoop_acc_4133_itm;
  wire [12:0] nl_MultLoop_acc_4133_itm;
  wire [15:0] MultLoop_acc_3683_itm_18_3_1;
  wire [15:0] MultLoop_acc_3532_itm_20_5_1;
  wire [14:0] MultLoop_acc_3281_itm_20_6;
  wire [16:0] MultLoop_acc_1943_itm_18_2;
  wire [18:0] MultLoop_acc_1811_itm_20_2_1;
  wire [15:0] MultLoop_acc_4587_itm_18_3;
  wire [15:0] MultLoop_acc_3190_itm_19_4;
  wire [18:0] MultLoop_acc_3338_itm_20_2_1;
  wire [15:0] MultLoop_acc_1753_itm_19_4;
  wire [12:0] MultLoop_acc_25_itm_17_5;
  wire [13:0] MultLoop_acc_3761_itm_19_6;
  wire [14:0] MultLoop_acc_67_itm_17_3;
  wire [16:0] MultLoop_acc_4588_itm_18_2;
  wire [15:0] MultLoop_acc_2317_itm_20_5;
  wire [14:0] MultLoop_acc_1097_itm_18_4;
  wire [15:0] MultLoop_acc_87_itm_19_4;
  wire [16:0] MultLoop_acc_1095_itm_18_2;
  wire [15:0] MultLoop_acc_3918_itm_17_2;
  wire [13:0] MultLoop_acc_447_itm_20_7;
  wire [14:0] MultLoop_acc_119_itm_23_9;
  wire [14:0] MultLoop_acc_123_itm_17_3;
  wire [15:0] MultLoop_acc_4589_itm_19_4;
  wire [17:0] MultLoop_acc_3556_itm_19_2_1;
  wire [15:0] MultLoop_acc_1145_itm_22_7;
  wire [18:0] MultLoop_acc_2409_itm_20_2_1;
  wire [14:0] MultLoop_acc_1128_itm_21_7;
  wire [14:0] MultLoop_acc_181_itm_22_8;
  wire [15:0] MultLoop_acc_3920_itm_17_2;
  wire [15:0] MultLoop_acc_2026_itm_21_6;
  wire [15:0] MultLoop_acc_149_itm_23_8;
  wire [18:0] MultLoop_acc_3213_itm_21_3_1;
  wire [15:0] MultLoop_acc_2252_itm_20_5;
  wire [15:0] MultLoop_acc_1154_itm_21_6;
  wire [15:0] MultLoop_acc_2040_itm_18_3;
  wire [15:0] MultLoop_acc_434_itm_22_7;
  wire [16:0] MultLoop_acc_2807_itm_18_2;
  wire [15:0] MultLoop_acc_1543_itm_21_6;
  wire [15:0] MultLoop_acc_1152_itm_18_3;
  wire [15:0] MultLoop_acc_1848_itm_21_6;
  wire [16:0] MultLoop_acc_1541_itm_18_2;
  wire [15:0] MultLoop_acc_3062_itm_19_4;
  wire [18:0] MultLoop_acc_1715_itm_20_2_1;
  wire [16:0] MultLoop_acc_1476_itm_18_2;
  wire [14:0] MultLoop_acc_307_itm_21_7;
  wire [15:0] MultLoop_acc_334_itm_20_5;
  wire [15:0] MultLoop_acc_2145_itm_20_5;
  wire [12:0] MultLoop_acc_335_itm_21_9;
  wire [16:0] MultLoop_acc_4594_itm_18_2;
  wire [13:0] MultLoop_acc_2836_itm_19_6;
  wire [14:0] MultLoop_acc_343_itm_19_5;
  wire [14:0] MultLoop_acc_340_itm_17_3;
  wire [15:0] MultLoop_acc_2289_itm_20_5;
  wire [14:0] MultLoop_acc_355_itm_20_6;
  wire [14:0] MultLoop_acc_1204_itm_19_5;
  wire [15:0] MultLoop_acc_1200_itm_19_4;
  wire [15:0] MultLoop_acc_2802_itm_19_4;
  wire [13:0] MultLoop_acc_410_itm_20_7;
  wire [14:0] MultLoop_acc_408_itm_23_9;
  wire [15:0] MultLoop_acc_2906_itm_19_4;
  wire [15:0] MultLoop_acc_400_itm_22_7;
  wire [16:0] MultLoop_acc_1227_itm_21_5;
  wire [15:0] MultLoop_acc_4590_itm_20_5;
  wire [14:0] MultLoop_acc_471_itm_21_7;
  wire [16:0] MultLoop_acc_1237_itm_20_4;
  wire [18:0] MultLoop_acc_2669_itm_20_2_1;
  wire [18:0] MultLoop_acc_1866_itm_20_2_1;
  wire [15:0] MultLoop_acc_3930_itm_17_2;
  wire [12:0] MultLoop_acc_506_itm_17_5;
  wire [15:0] MultLoop_acc_2340_itm_19_4;
  wire [14:0] MultLoop_acc_528_itm_24_10;
  wire [15:0] MultLoop_acc_541_itm_23_8;
  wire [15:0] MultLoop_acc_1275_itm_20_5;
  wire [15:0] MultLoop_acc_579_itm_19_4;
  wire [15:0] MultLoop_acc_570_itm_21_6;
  wire [15:0] MultLoop_acc_1730_itm_22_7;
  wire [18:0] MultLoop_acc_1816_itm_20_2_1;
  wire [15:0] MultLoop_acc_713_itm_23_8;
  wire [13:0] MultLoop_acc_785_itm_17_4;
  wire [15:0] MultLoop_acc_4663_itm_19_4;
  wire [15:0] MultLoop_acc_826_itm_25_10;
  wire [15:0] MultLoop_acc_1479_itm_18_3;
  wire [15:0] MultLoop_acc_4592_itm_18_3;
  wire [15:0] MultLoop_acc_4593_itm_18_3;
  wire [15:0] MultLoop_acc_1350_itm_22_7;
  wire [15:0] MultLoop_acc_807_itm_21_6;
  wire [18:0] MultLoop_acc_1512_itm_20_2_1;
  wire [18:0] Result_acc_102_itm_20_2_1;
  wire [16:0] MultLoop_acc_1993_itm_18_2;
  wire [15:0] MultLoop_acc_856_itm_22_7;
  wire [15:0] Result_acc_154_itm_19_4;
  wire [16:0] MultLoop_acc_4591_itm_18_2;
  wire [13:0] MultLoop_acc_150_itm_17_4;
  wire [14:0] MultLoop_acc_1191_itm_21_7;
  wire [15:0] MultLoop_acc_1211_itm_23_8;
  wire [13:0] MultLoop_acc_1243_itm_19_6;
  wire [15:0] MultLoop_acc_1315_itm_19_4;
  wire [15:0] MultLoop_acc_1324_itm_22_7;

  wire[17:0] MultLoop_acc_1591_nl;
  wire[19:0] nl_MultLoop_acc_1591_nl;
  wire[17:0] MultLoop_acc_1587_nl;
  wire[19:0] nl_MultLoop_acc_1587_nl;
  wire[17:0] MultLoop_acc_3912_nl;
  wire[20:0] nl_MultLoop_acc_3912_nl;
  wire[17:0] MultLoop_acc_1686_nl;
  wire[19:0] nl_MultLoop_acc_1686_nl;
  wire[17:0] MultLoop_acc_1682_nl;
  wire[19:0] nl_MultLoop_acc_1682_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl;
  wire[17:0] MultLoop_acc_1799_nl;
  wire[20:0] nl_MultLoop_acc_1799_nl;
  wire[17:0] MultLoop_acc_3731_nl;
  wire[19:0] nl_MultLoop_acc_3731_nl;
  wire[17:0] MultLoop_acc_3729_nl;
  wire[19:0] nl_MultLoop_acc_3729_nl;
  wire[17:0] MultLoop_acc_3727_nl;
  wire[18:0] nl_MultLoop_acc_3727_nl;
  wire[17:0] MultLoop_acc_3613_nl;
  wire[19:0] nl_MultLoop_acc_3613_nl;
  wire[17:0] MultLoop_acc_3608_nl;
  wire[19:0] nl_MultLoop_acc_3608_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl;
  wire[17:0] MultLoop_acc_3498_nl;
  wire[20:0] nl_MultLoop_acc_3498_nl;
  wire[17:0] MultLoop_acc_2123_nl;
  wire[19:0] nl_MultLoop_acc_2123_nl;
  wire[17:0] MultLoop_acc_3381_nl;
  wire[19:0] nl_MultLoop_acc_3381_nl;
  wire[17:0] MultLoop_acc_3377_nl;
  wire[18:0] nl_MultLoop_acc_3377_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl;
  wire[17:0] MultLoop_acc_3263_nl;
  wire[19:0] nl_MultLoop_acc_3263_nl;
  wire[17:0] MultLoop_acc_3261_nl;
  wire[19:0] nl_MultLoop_acc_3261_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl;
  wire[16:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl;
  wire[17:0] MultLoop_acc_2473_nl;
  wire[20:0] nl_MultLoop_acc_2473_nl;
  wire[17:0] MultLoop_acc_3021_nl;
  wire[19:0] nl_MultLoop_acc_3021_nl;
  wire[17:0] MultLoop_acc_3017_nl;
  wire[19:0] nl_MultLoop_acc_3017_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl;
  wire[20:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl;
  wire[17:0] MultLoop_acc_2899_nl;
  wire[19:0] nl_MultLoop_acc_2899_nl;
  wire[17:0] MultLoop_acc_2895_nl;
  wire[19:0] nl_MultLoop_acc_2895_nl;
  wire[17:0] MultLoop_acc_2661_nl;
  wire[19:0] nl_MultLoop_acc_2661_nl;
  wire[17:0] MultLoop_acc_2777_nl;
  wire[20:0] nl_MultLoop_acc_2777_nl;
  wire[17:0] MultLoop_acc_2776_nl;
  wire[19:0] nl_MultLoop_acc_2776_nl;
  wire[26:0] Result_acc_17_nl;
  wire[27:0] nl_Result_acc_17_nl;
  wire[24:0] Result_acc_77_nl;
  wire[25:0] nl_Result_acc_77_nl;
  wire[17:0] Result_acc_146_nl;
  wire[18:0] nl_Result_acc_146_nl;
  wire[10:0] Result_acc_181_nl;
  wire[11:0] nl_Result_acc_181_nl;
  wire[21:0] Result_acc_59_nl;
  wire[22:0] nl_Result_acc_59_nl;
  wire[18:0] Result_acc_142_nl;
  wire[19:0] nl_Result_acc_142_nl;
  wire[21:0] Result_acc_75_nl;
  wire[22:0] nl_Result_acc_75_nl;
  wire[21:0] Result_acc_23_nl;
  wire[22:0] nl_Result_acc_23_nl;
  wire[21:0] Result_acc_55_nl;
  wire[22:0] nl_Result_acc_55_nl;
  wire[15:0] Result_acc_179_nl;
  wire[16:0] nl_Result_acc_179_nl;
  wire[20:0] Result_acc_57_nl;
  wire[21:0] nl_Result_acc_57_nl;
  wire[22:0] Result_acc_78_nl;
  wire[23:0] nl_Result_acc_78_nl;
  wire[19:0] Result_acc_149_nl;
  wire[21:0] nl_Result_acc_149_nl;
  wire[22:0] Result_acc_79_nl;
  wire[23:0] nl_Result_acc_79_nl;
  wire[17:0] Result_acc_151_nl;
  wire[18:0] nl_Result_acc_151_nl;
  wire[23:0] Result_acc_29_nl;
  wire[25:0] nl_Result_acc_29_nl;
  wire[13:0] Result_acc_184_nl;
  wire[14:0] nl_Result_acc_184_nl;
  wire[18:0] Result_acc_63_nl;
  wire[19:0] nl_Result_acc_63_nl;
  wire[19:0] Result_acc_217_nl;
  wire[20:0] nl_Result_acc_217_nl;
  wire[20:0] Result_acc_64_nl;
  wire[21:0] nl_Result_acc_64_nl;
  wire[17:0] Result_acc_88_nl;
  wire[18:0] nl_Result_acc_88_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[18:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl;
  wire[20:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl;
  wire[21:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl;
  wire[23:0] Result_acc_38_nl;
  wire[24:0] nl_Result_acc_38_nl;
  wire[21:0] Result_acc_89_nl;
  wire[22:0] nl_Result_acc_89_nl;
  wire[12:0] MultLoop_acc_1548_nl;
  wire[14:0] nl_MultLoop_acc_1548_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_9_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_10_nl;
  wire[17:0] Result_acc_186_nl;
  wire[18:0] nl_Result_acc_186_nl;
  wire[22:0] Result_acc_92_nl;
  wire[24:0] nl_Result_acc_92_nl;
  wire[11:0] Result_acc_185_nl;
  wire[12:0] nl_Result_acc_185_nl;
  wire[19:0] Result_acc_65_nl;
  wire[20:0] nl_Result_acc_65_nl;
  wire[17:0] Result_acc_93_nl;
  wire[18:0] nl_Result_acc_93_nl;
  wire[21:0] Result_acc_22_nl;
  wire[22:0] nl_Result_acc_22_nl;
  wire[20:0] Result_acc_96_nl;
  wire[22:0] nl_Result_acc_96_nl;
  wire[17:0] Result_acc_189_nl;
  wire[18:0] nl_Result_acc_189_nl;
  wire[21:0] Result_acc_99_nl;
  wire[23:0] nl_Result_acc_99_nl;
  wire[20:0] Result_acc_66_nl;
  wire[21:0] nl_Result_acc_66_nl;
  wire[17:0] Result_acc_101_nl;
  wire[18:0] nl_Result_acc_101_nl;
  wire[20:0] Result_acc_219_nl;
  wire[21:0] nl_Result_acc_219_nl;
  wire[22:0] Result_acc_67_nl;
  wire[23:0] nl_Result_acc_67_nl;
  wire[18:0] Result_acc_103_nl;
  wire[19:0] nl_Result_acc_103_nl;
  wire[21:0] Result_acc_68_nl;
  wire[22:0] nl_Result_acc_68_nl;
  wire[17:0] Result_acc_104_nl;
  wire[18:0] nl_Result_acc_104_nl;
  wire[23:0] Result_acc_70_nl;
  wire[24:0] nl_Result_acc_70_nl;
  wire[21:0] Result_acc_112_nl;
  wire[22:0] nl_Result_acc_112_nl;
  wire[22:0] Result_acc_71_nl;
  wire[23:0] nl_Result_acc_71_nl;
  wire[20:0] Result_acc_114_nl;
  wire[22:0] nl_Result_acc_114_nl;
  wire[19:0] Result_acc_54_nl;
  wire[20:0] nl_Result_acc_54_nl;
  wire[18:0] Result_acc_106_nl;
  wire[19:0] nl_Result_acc_106_nl;
  wire[20:0] Result_acc_69_nl;
  wire[21:0] nl_Result_acc_69_nl;
  wire[17:0] Result_acc_108_nl;
  wire[18:0] nl_Result_acc_108_nl;
  wire[20:0] Result_acc_58_nl;
  wire[21:0] nl_Result_acc_58_nl;
  wire[18:0] Result_acc_110_nl;
  wire[19:0] nl_Result_acc_110_nl;
  wire[12:0] Result_acc_193_nl;
  wire[13:0] nl_Result_acc_193_nl;
  wire[20:0] Result_acc_30_nl;
  wire[21:0] nl_Result_acc_30_nl;
  wire[20:0] Result_acc_62_nl;
  wire[21:0] nl_Result_acc_62_nl;
  wire[17:0] Result_acc_83_nl;
  wire[18:0] nl_Result_acc_83_nl;
  wire[21:0] Result_acc_72_nl;
  wire[22:0] nl_Result_acc_72_nl;
  wire[18:0] Result_acc_120_nl;
  wire[19:0] nl_Result_acc_120_nl;
  wire[17:0] Result_acc_196_nl;
  wire[18:0] nl_Result_acc_196_nl;
  wire[23:0] Result_acc_116_nl;
  wire[24:0] nl_Result_acc_116_nl;
  wire[17:0] Result_acc_26_nl;
  wire[18:0] nl_Result_acc_26_nl;
  wire[17:0] Result_acc_198_nl;
  wire[18:0] nl_Result_acc_198_nl;
  wire[23:0] Result_acc_119_nl;
  wire[24:0] nl_Result_acc_119_nl;
  wire[19:0] Result_acc_118_nl;
  wire[20:0] nl_Result_acc_118_nl;
  wire[17:0] Result_acc_200_nl;
  wire[18:0] nl_Result_acc_200_nl;
  wire[22:0] Result_acc_123_nl;
  wire[23:0] nl_Result_acc_123_nl;
  wire[19:0] Result_acc_122_nl;
  wire[20:0] nl_Result_acc_122_nl;
  wire[21:0] Result_acc_40_nl;
  wire[22:0] nl_Result_acc_40_nl;
  wire[18:0] Result_acc_125_nl;
  wire[19:0] nl_Result_acc_125_nl;
  wire[25:0] Result_acc_43_nl;
  wire[26:0] nl_Result_acc_43_nl;
  wire[23:0] Result_acc_126_nl;
  wire[24:0] nl_Result_acc_126_nl;
  wire[18:0] Result_acc_218_nl;
  wire[19:0] nl_Result_acc_218_nl;
  wire[17:0] Result_acc_203_nl;
  wire[18:0] nl_Result_acc_203_nl;
  wire[21:0] Result_acc_220_nl;
  wire[22:0] nl_Result_acc_220_nl;
  wire[25:0] Result_acc_48_nl;
  wire[27:0] nl_Result_acc_48_nl;
  wire[23:0] Result_acc_74_nl;
  wire[24:0] nl_Result_acc_74_nl;
  wire[19:0] Result_acc_136_nl;
  wire[21:0] nl_Result_acc_136_nl;
  wire[11:0] Result_acc_205_nl;
  wire[12:0] nl_Result_acc_205_nl;
  wire[23:0] Result_acc_51_nl;
  wire[24:0] nl_Result_acc_51_nl;
  wire[21:0] Result_acc_137_nl;
  wire[22:0] nl_Result_acc_137_nl;
  wire[22:0] Result_acc_53_nl;
  wire[23:0] nl_Result_acc_53_nl;
  wire[21:0] Result_acc_140_nl;
  wire[23:0] nl_Result_acc_140_nl;
  wire[17:0] MultLoop_acc_3908_nl;
  wire[19:0] nl_MultLoop_acc_3908_nl;
  wire[23:0] MultLoop_acc_1080_nl;
  wire[24:0] nl_MultLoop_acc_1080_nl;
  wire[20:0] MultLoop_acc_3865_nl;
  wire[21:0] nl_MultLoop_acc_3865_nl;
  wire[17:0] MultLoop_acc_3864_nl;
  wire[18:0] nl_MultLoop_acc_3864_nl;
  wire[22:0] MultLoop_acc_18_nl;
  wire[23:0] nl_MultLoop_acc_18_nl;
  wire[14:0] MultLoop_acc_4565_nl;
  wire[15:0] nl_MultLoop_acc_4565_nl;
  wire[25:0] MultLoop_acc_13_nl;
  wire[26:0] nl_MultLoop_acc_13_nl;
  wire[18:0] MultLoop_acc_4567_nl;
  wire[19:0] nl_MultLoop_acc_4567_nl;
  wire[17:0] MultLoop_acc_15_nl;
  wire[18:0] nl_MultLoop_acc_15_nl;
  wire[17:0] MultLoop_acc_4559_nl;
  wire[18:0] nl_MultLoop_acc_4559_nl;
  wire[22:0] MultLoop_acc_3854_nl;
  wire[23:0] nl_MultLoop_acc_3854_nl;
  wire[23:0] MultLoop_acc_4658_nl;
  wire[24:0] nl_MultLoop_acc_4658_nl;
  wire[18:0] MultLoop_acc_4563_nl;
  wire[19:0] nl_MultLoop_acc_4563_nl;
  wire[25:0] MultLoop_acc_2_nl;
  wire[26:0] nl_MultLoop_acc_2_nl;
  wire[24:0] MultLoop_acc_3863_nl;
  wire[25:0] nl_MultLoop_acc_3863_nl;
  wire[11:0] MultLoop_acc_4564_nl;
  wire[12:0] nl_MultLoop_acc_4564_nl;
  wire[17:0] MultLoop_acc_4561_nl;
  wire[18:0] nl_MultLoop_acc_4561_nl;
  wire[20:0] MultLoop_acc_3856_nl;
  wire[21:0] nl_MultLoop_acc_3856_nl;
  wire[12:0] MultLoop_acc_4560_nl;
  wire[13:0] nl_MultLoop_acc_4560_nl;
  wire[21:0] MultLoop_acc_7_nl;
  wire[22:0] nl_MultLoop_acc_7_nl;
  wire[19:0] MultLoop_acc_3859_nl;
  wire[20:0] nl_MultLoop_acc_3859_nl;
  wire[17:0] MultLoop_acc_3858_nl;
  wire[18:0] nl_MultLoop_acc_3858_nl;
  wire[10:0] MultLoop_acc_4562_nl;
  wire[11:0] nl_MultLoop_acc_4562_nl;
  wire[17:0] MultLoop_acc_38_nl;
  wire[18:0] nl_MultLoop_acc_38_nl;
  wire[17:0] MultLoop_acc_27_nl;
  wire[18:0] nl_MultLoop_acc_27_nl;
  wire[23:0] MultLoop_acc_46_nl;
  wire[24:0] nl_MultLoop_acc_46_nl;
  wire[21:0] MultLoop_acc_3800_nl;
  wire[22:0] nl_MultLoop_acc_3800_nl;
  wire[19:0] MultLoop_acc_3799_nl;
  wire[20:0] nl_MultLoop_acc_3799_nl;
  wire[17:0] MultLoop_acc_45_nl;
  wire[18:0] nl_MultLoop_acc_45_nl;
  wire[20:0] MultLoop_acc_21_nl;
  wire[21:0] nl_MultLoop_acc_21_nl;
  wire[18:0] MultLoop_acc_3803_nl;
  wire[19:0] nl_MultLoop_acc_3803_nl;
  wire[12:0] MultLoop_acc_4568_nl;
  wire[13:0] nl_MultLoop_acc_4568_nl;
  wire[22:0] MultLoop_acc_47_nl;
  wire[23:0] nl_MultLoop_acc_47_nl;
  wire[20:0] MultLoop_acc_3805_nl;
  wire[21:0] nl_MultLoop_acc_3805_nl;
  wire[13:0] MultLoop_acc_4569_nl;
  wire[14:0] nl_MultLoop_acc_4569_nl;
  wire[17:0] MultLoop_acc_4659_nl;
  wire[18:0] nl_MultLoop_acc_4659_nl;
  wire[17:0] MultLoop_acc_4572_nl;
  wire[18:0] nl_MultLoop_acc_4572_nl;
  wire[21:0] MultLoop_acc_3810_nl;
  wire[23:0] nl_MultLoop_acc_3810_nl;
  wire[17:0] MultLoop_acc_4574_nl;
  wire[18:0] nl_MultLoop_acc_4574_nl;
  wire[22:0] MultLoop_acc_3813_nl;
  wire[24:0] nl_MultLoop_acc_3813_nl;
  wire[17:0] MultLoop_acc_33_nl;
  wire[18:0] nl_MultLoop_acc_33_nl;
  wire[20:0] MultLoop_acc_4660_nl;
  wire[21:0] nl_MultLoop_acc_4660_nl;
  wire[19:0] MultLoop_acc_4661_nl;
  wire[20:0] nl_MultLoop_acc_4661_nl;
  wire[17:0] MultLoop_acc_4576_nl;
  wire[18:0] nl_MultLoop_acc_4576_nl;
  wire[21:0] MultLoop_acc_3818_nl;
  wire[22:0] nl_MultLoop_acc_3818_nl;
  wire[21:0] MultLoop_acc_1079_nl;
  wire[22:0] nl_MultLoop_acc_1079_nl;
  wire[19:0] MultLoop_acc_3820_nl;
  wire[20:0] nl_MultLoop_acc_3820_nl;
  wire[22:0] MultLoop_acc_1076_nl;
  wire[23:0] nl_MultLoop_acc_1076_nl;
  wire[19:0] MultLoop_acc_3823_nl;
  wire[21:0] nl_MultLoop_acc_3823_nl;
  wire[24:0] MultLoop_acc_11_nl;
  wire[25:0] nl_MultLoop_acc_11_nl;
  wire[23:0] MultLoop_acc_3825_nl;
  wire[25:0] nl_MultLoop_acc_3825_nl;
  wire[21:0] MultLoop_acc_1075_nl;
  wire[22:0] nl_MultLoop_acc_1075_nl;
  wire[19:0] MultLoop_acc_3827_nl;
  wire[21:0] nl_MultLoop_acc_3827_nl;
  wire[21:0] MultLoop_acc_43_nl;
  wire[22:0] nl_MultLoop_acc_43_nl;
  wire[18:0] MultLoop_acc_3832_nl;
  wire[19:0] nl_MultLoop_acc_3832_nl;
  wire[21:0] MultLoop_acc_40_nl;
  wire[22:0] nl_MultLoop_acc_40_nl;
  wire[19:0] MultLoop_acc_3835_nl;
  wire[20:0] nl_MultLoop_acc_3835_nl;
  wire[17:0] MultLoop_acc_3834_nl;
  wire[18:0] nl_MultLoop_acc_3834_nl;
  wire[12:0] MultLoop_acc_4580_nl;
  wire[13:0] nl_MultLoop_acc_4580_nl;
  wire[20:0] MultLoop_acc_1087_nl;
  wire[21:0] nl_MultLoop_acc_1087_nl;
  wire[20:0] MultLoop_acc_1088_nl;
  wire[21:0] nl_MultLoop_acc_1088_nl;
  wire[17:0] MultLoop_acc_3830_nl;
  wire[18:0] nl_MultLoop_acc_3830_nl;
  wire[17:0] MultLoop_acc_42_nl;
  wire[18:0] nl_MultLoop_acc_42_nl;
  wire[19:0] MultLoop_acc_4582_nl;
  wire[20:0] nl_MultLoop_acc_4582_nl;
  wire[17:0] MultLoop_acc_4581_nl;
  wire[18:0] nl_MultLoop_acc_4581_nl;
  wire[23:0] MultLoop_acc_1078_nl;
  wire[24:0] nl_MultLoop_acc_1078_nl;
  wire[20:0] MultLoop_acc_3847_nl;
  wire[22:0] nl_MultLoop_acc_3847_nl;
  wire[11:0] MultLoop_acc_4586_nl;
  wire[12:0] nl_MultLoop_acc_4586_nl;
  wire[23:0] MultLoop_acc_1077_nl;
  wire[24:0] nl_MultLoop_acc_1077_nl;
  wire[22:0] MultLoop_acc_3850_nl;
  wire[23:0] nl_MultLoop_acc_3850_nl;
  wire[19:0] MultLoop_acc_3849_nl;
  wire[20:0] nl_MultLoop_acc_3849_nl;
  wire[21:0] MultLoop_acc_31_nl;
  wire[22:0] nl_MultLoop_acc_31_nl;
  wire[15:0] MultLoop_acc_4583_nl;
  wire[16:0] nl_MultLoop_acc_4583_nl;
  wire[21:0] MultLoop_acc_1084_nl;
  wire[22:0] nl_MultLoop_acc_1084_nl;
  wire[21:0] MultLoop_acc_1083_nl;
  wire[22:0] nl_MultLoop_acc_1083_nl;
  wire[20:0] MultLoop_acc_3841_nl;
  wire[21:0] nl_MultLoop_acc_3841_nl;
  wire[17:0] MultLoop_acc_4585_nl;
  wire[18:0] nl_MultLoop_acc_4585_nl;
  wire[20:0] MultLoop_acc_3844_nl;
  wire[22:0] nl_MultLoop_acc_3844_nl;
  wire[23:0] MultLoop_acc_17_nl;
  wire[24:0] nl_MultLoop_acc_17_nl;
  wire[25:0] MultLoop_acc_14_nl;
  wire[26:0] nl_MultLoop_acc_14_nl;
  wire[24:0] MultLoop_acc_3852_nl;
  wire[25:0] nl_MultLoop_acc_3852_nl;
  wire[23:0] MultLoop_acc_1443_nl;
  wire[24:0] nl_MultLoop_acc_1443_nl;
  wire[20:0] MultLoop_acc_1640_nl;
  wire[22:0] nl_MultLoop_acc_1640_nl;
  wire[11:0] MultLoop_acc_3940_nl;
  wire[12:0] nl_MultLoop_acc_3940_nl;
  wire[22:0] MultLoop_acc_1435_nl;
  wire[23:0] nl_MultLoop_acc_1435_nl;
  wire[17:0] MultLoop_acc_1642_nl;
  wire[18:0] nl_MultLoop_acc_1642_nl;
  wire[21:0] Result_acc_80_nl;
  wire[22:0] nl_Result_acc_80_nl;
  wire[17:0] Result_acc_171_nl;
  wire[18:0] nl_Result_acc_171_nl;
  wire[13:0] Result_acc_207_nl;
  wire[14:0] nl_Result_acc_207_nl;
  wire[25:0] Result_acc_8_nl;
  wire[27:0] nl_Result_acc_8_nl;
  wire[26:0] Result_acc_11_nl;
  wire[28:0] nl_Result_acc_11_nl;
  wire[25:0] Result_acc_16_nl;
  wire[27:0] nl_Result_acc_16_nl;
  wire[17:0] MultLoop_acc_3943_nl;
  wire[18:0] nl_MultLoop_acc_3943_nl;
  wire[19:0] MultLoop_acc_1596_nl;
  wire[20:0] nl_MultLoop_acc_1596_nl;
  wire[12:0] MultLoop_acc_3942_nl;
  wire[13:0] nl_MultLoop_acc_3942_nl;
  wire[19:0] MultLoop_acc_1439_nl;
  wire[20:0] nl_MultLoop_acc_1439_nl;
  wire[17:0] MultLoop_acc_1597_nl;
  wire[18:0] nl_MultLoop_acc_1597_nl;
  wire[21:0] MultLoop_acc_1059_nl;
  wire[22:0] nl_MultLoop_acc_1059_nl;
  wire[19:0] MultLoop_acc_1600_nl;
  wire[20:0] nl_MultLoop_acc_1600_nl;
  wire[17:0] MultLoop_acc_1599_nl;
  wire[18:0] nl_MultLoop_acc_1599_nl;
  wire[23:0] MultLoop_acc_1049_nl;
  wire[25:0] nl_MultLoop_acc_1049_nl;
  wire[13:0] MultLoop_acc_3945_nl;
  wire[14:0] nl_MultLoop_acc_3945_nl;
  wire[22:0] Result_acc_5_nl;
  wire[23:0] nl_Result_acc_5_nl;
  wire[19:0] Result_acc_153_nl;
  wire[20:0] nl_Result_acc_153_nl;
  wire[19:0] Result_acc_222_nl;
  wire[20:0] nl_Result_acc_222_nl;
  wire[17:0] Result_acc_7_nl;
  wire[18:0] nl_Result_acc_7_nl;
  wire[24:0] MultLoop_acc_1070_nl;
  wire[25:0] nl_MultLoop_acc_1070_nl;
  wire[23:0] MultLoop_acc_1604_nl;
  wire[24:0] nl_MultLoop_acc_1604_nl;
  wire[22:0] MultLoop_acc_1068_nl;
  wire[23:0] nl_MultLoop_acc_1068_nl;
  wire[21:0] MultLoop_acc_1441_nl;
  wire[22:0] nl_MultLoop_acc_1441_nl;
  wire[20:0] MultLoop_acc_1606_nl;
  wire[21:0] nl_MultLoop_acc_1606_nl;
  wire[17:0] MultLoop_acc_1605_nl;
  wire[18:0] nl_MultLoop_acc_1605_nl;
  wire[19:0] Result_acc_9_nl;
  wire[20:0] nl_Result_acc_9_nl;
  wire[18:0] Result_acc_157_nl;
  wire[19:0] nl_Result_acc_157_nl;
  wire[14:0] Result_acc_211_nl;
  wire[15:0] nl_Result_acc_211_nl;
  wire[18:0] MultLoop_acc_1442_nl;
  wire[19:0] nl_MultLoop_acc_1442_nl;
  wire[22:0] MultLoop_acc_1440_nl;
  wire[23:0] nl_MultLoop_acc_1440_nl;
  wire[19:0] MultLoop_acc_1609_nl;
  wire[21:0] nl_MultLoop_acc_1609_nl;
  wire[24:0] MultLoop_acc_1062_nl;
  wire[25:0] nl_MultLoop_acc_1062_nl;
  wire[19:0] MultLoop_acc_1610_nl;
  wire[20:0] nl_MultLoop_acc_1610_nl;
  wire[21:0] MultLoop_acc_1436_nl;
  wire[22:0] nl_MultLoop_acc_1436_nl;
  wire[19:0] MultLoop_acc_1612_nl;
  wire[20:0] nl_MultLoop_acc_1612_nl;
  wire[24:0] MultLoop_acc_1053_nl;
  wire[26:0] nl_MultLoop_acc_1053_nl;
  wire[24:0] MultLoop_acc_1054_nl;
  wire[25:0] nl_MultLoop_acc_1054_nl;
  wire[22:0] MultLoop_acc_1616_nl;
  wire[23:0] nl_MultLoop_acc_1616_nl;
  wire[19:0] MultLoop_acc_1615_nl;
  wire[20:0] nl_MultLoop_acc_1615_nl;
  wire[20:0] MultLoop_acc_1051_nl;
  wire[21:0] nl_MultLoop_acc_1051_nl;
  wire[17:0] MultLoop_acc_3949_nl;
  wire[18:0] nl_MultLoop_acc_3949_nl;
  wire[20:0] MultLoop_acc_4662_nl;
  wire[21:0] nl_MultLoop_acc_4662_nl;
  wire[17:0] Result_acc_213_nl;
  wire[18:0] nl_Result_acc_213_nl;
  wire[22:0] Result_acc_160_nl;
  wire[24:0] nl_Result_acc_160_nl;
  wire[21:0] MultLoop_acc_1067_nl;
  wire[22:0] nl_MultLoop_acc_1067_nl;
  wire[18:0] MultLoop_acc_1621_nl;
  wire[19:0] nl_MultLoop_acc_1621_nl;
  wire[11:0] MultLoop_acc_3950_nl;
  wire[12:0] nl_MultLoop_acc_3950_nl;
  wire[20:0] Result_acc_81_nl;
  wire[21:0] nl_Result_acc_81_nl;
  wire[17:0] Result_acc_161_nl;
  wire[18:0] nl_Result_acc_161_nl;
  wire[19:0] Result_acc_nl;
  wire[20:0] nl_Result_acc_nl;
  wire[10:0] MultLoop_acc_1643_nl;
  wire[11:0] nl_MultLoop_acc_1643_nl;
  wire[17:0] Result_acc_2_nl;
  wire[18:0] nl_Result_acc_2_nl;
  wire[17:0] MultLoop_acc_1073_nl;
  wire[18:0] nl_MultLoop_acc_1073_nl;
  wire[19:0] MultLoop_acc_1434_nl;
  wire[20:0] nl_MultLoop_acc_1434_nl;
  wire[17:0] MultLoop_acc_1627_nl;
  wire[18:0] nl_MultLoop_acc_1627_nl;
  wire[22:0] MultLoop_acc_1052_nl;
  wire[23:0] nl_MultLoop_acc_1052_nl;
  wire[21:0] MultLoop_acc_1630_nl;
  wire[23:0] nl_MultLoop_acc_1630_nl;
  wire[10:0] MultLoop_acc_3952_nl;
  wire[11:0] nl_MultLoop_acc_3952_nl;
  wire[25:0] MultLoop_acc_1065_nl;
  wire[27:0] nl_MultLoop_acc_1065_nl;
  wire[22:0] MultLoop_acc_1438_nl;
  wire[23:0] nl_MultLoop_acc_1438_nl;
  wire[19:0] MultLoop_acc_1625_nl;
  wire[20:0] nl_MultLoop_acc_1625_nl;
  wire[17:0] MultLoop_acc_1624_nl;
  wire[18:0] nl_MultLoop_acc_1624_nl;
  wire[19:0] MultLoop_acc_1437_nl;
  wire[20:0] nl_MultLoop_acc_1437_nl;
  wire[19:0] MultLoop_acc_1050_nl;
  wire[20:0] nl_MultLoop_acc_1050_nl;
  wire[18:0] MultLoop_acc_1632_nl;
  wire[19:0] nl_MultLoop_acc_1632_nl;
  wire[11:0] MultLoop_acc_3953_nl;
  wire[12:0] nl_MultLoop_acc_3953_nl;
  wire[20:0] MultLoop_acc_1432_nl;
  wire[21:0] nl_MultLoop_acc_1432_nl;
  wire[17:0] MultLoop_acc_1634_nl;
  wire[18:0] nl_MultLoop_acc_1634_nl;
  wire[13:0] MultLoop_acc_3954_nl;
  wire[14:0] nl_MultLoop_acc_3954_nl;
  wire[22:0] MultLoop_acc_1046_nl;
  wire[23:0] nl_MultLoop_acc_1046_nl;
  wire[19:0] MultLoop_acc_1637_nl;
  wire[20:0] nl_MultLoop_acc_1637_nl;
  wire[22:0] Result_acc_10_nl;
  wire[23:0] nl_Result_acc_10_nl;
  wire[21:0] Result_acc_164_nl;
  wire[22:0] nl_Result_acc_164_nl;
  wire[19:0] Result_acc_14_nl;
  wire[20:0] nl_Result_acc_14_nl;
  wire[18:0] Result_acc_166_nl;
  wire[19:0] nl_Result_acc_166_nl;
  wire[14:0] Result_acc_215_nl;
  wire[15:0] nl_Result_acc_215_nl;
  wire[22:0] Result_acc_15_nl;
  wire[23:0] nl_Result_acc_15_nl;
  wire[21:0] Result_acc_169_nl;
  wire[23:0] nl_Result_acc_169_nl;
  wire[25:0] MultLoop_acc_74_nl;
  wire[26:0] nl_MultLoop_acc_74_nl;
  wire[21:0] MultLoop_acc_3795_nl;
  wire[22:0] nl_MultLoop_acc_3795_nl;
  wire[19:0] MultLoop_acc_3794_nl;
  wire[20:0] nl_MultLoop_acc_3794_nl;
  wire[22:0] MultLoop_acc_66_nl;
  wire[23:0] nl_MultLoop_acc_66_nl;
  wire[14:0] MultLoop_acc_4529_nl;
  wire[15:0] nl_MultLoop_acc_4529_nl;
  wire[21:0] MultLoop_acc_1089_nl;
  wire[22:0] nl_MultLoop_acc_1089_nl;
  wire[17:0] MultLoop_acc_3798_nl;
  wire[18:0] nl_MultLoop_acc_3798_nl;
  wire[12:0] MultLoop_acc_4530_nl;
  wire[13:0] nl_MultLoop_acc_4530_nl;
  wire[21:0] MultLoop_acc_90_nl;
  wire[22:0] nl_MultLoop_acc_90_nl;
  wire[19:0] MultLoop_acc_3741_nl;
  wire[20:0] nl_MultLoop_acc_3741_nl;
  wire[17:0] MultLoop_acc_3740_nl;
  wire[18:0] nl_MultLoop_acc_3740_nl;
  wire[20:0] MultLoop_acc_84_nl;
  wire[21:0] nl_MultLoop_acc_84_nl;
  wire[18:0] MultLoop_acc_3743_nl;
  wire[19:0] nl_MultLoop_acc_3743_nl;
  wire[13:0] MultLoop_acc_4532_nl;
  wire[14:0] nl_MultLoop_acc_4532_nl;
  wire[20:0] MultLoop_acc_1091_nl;
  wire[21:0] nl_MultLoop_acc_1091_nl;
  wire[18:0] MultLoop_acc_3744_nl;
  wire[19:0] nl_MultLoop_acc_3744_nl;
  wire[17:0] MultLoop_acc_59_nl;
  wire[18:0] nl_MultLoop_acc_59_nl;
  wire[19:0] MultLoop_acc_60_nl;
  wire[20:0] nl_MultLoop_acc_60_nl;
  wire[18:0] MultLoop_acc_3746_nl;
  wire[19:0] nl_MultLoop_acc_3746_nl;
  wire[13:0] MultLoop_acc_4533_nl;
  wire[14:0] nl_MultLoop_acc_4533_nl;
  wire[21:0] MultLoop_acc_1090_nl;
  wire[22:0] nl_MultLoop_acc_1090_nl;
  wire[17:0] MultLoop_acc_4535_nl;
  wire[18:0] nl_MultLoop_acc_4535_nl;
  wire[21:0] MultLoop_acc_3749_nl;
  wire[22:0] nl_MultLoop_acc_3749_nl;
  wire[12:0] MultLoop_acc_4534_nl;
  wire[13:0] nl_MultLoop_acc_4534_nl;
  wire[21:0] MultLoop_acc_1099_nl;
  wire[22:0] nl_MultLoop_acc_1099_nl;
  wire[21:0] MultLoop_acc_52_nl;
  wire[22:0] nl_MultLoop_acc_52_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl;
  wire[13:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl;
  wire[20:0] MultLoop_acc_69_nl;
  wire[21:0] nl_MultLoop_acc_69_nl;
  wire[16:0] MultLoop_acc_4536_nl;
  wire[17:0] nl_MultLoop_acc_4536_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl;
  wire[24:0] MultLoop_acc_85_nl;
  wire[25:0] nl_MultLoop_acc_85_nl;
  wire[21:0] MultLoop_acc_3753_nl;
  wire[22:0] nl_MultLoop_acc_3753_nl;
  wire[19:0] MultLoop_acc_3752_nl;
  wire[20:0] nl_MultLoop_acc_3752_nl;
  wire[12:0] MultLoop_acc_4537_nl;
  wire[13:0] nl_MultLoop_acc_4537_nl;
  wire[22:0] MultLoop_acc_73_nl;
  wire[23:0] nl_MultLoop_acc_73_nl;
  wire[20:0] MultLoop_acc_3755_nl;
  wire[21:0] nl_MultLoop_acc_3755_nl;
  wire[24:0] MultLoop_acc_71_nl;
  wire[25:0] nl_MultLoop_acc_71_nl;
  wire[21:0] MultLoop_acc_3756_nl;
  wire[22:0] nl_MultLoop_acc_3756_nl;
  wire[24:0] MultLoop_acc_65_nl;
  wire[25:0] nl_MultLoop_acc_65_nl;
  wire[21:0] MultLoop_acc_3759_nl;
  wire[22:0] nl_MultLoop_acc_3759_nl;
  wire[19:0] MultLoop_acc_3758_nl;
  wire[20:0] nl_MultLoop_acc_3758_nl;
  wire[12:0] MultLoop_acc_4539_nl;
  wire[13:0] nl_MultLoop_acc_4539_nl;
  wire[18:0] MultLoop_acc_4655_nl;
  wire[19:0] nl_MultLoop_acc_4655_nl;
  wire[14:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl;
  wire[18:0] MultLoop_acc_4656_nl;
  wire[19:0] nl_MultLoop_acc_4656_nl;
  wire[13:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl;
  wire[14:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl;
  wire[21:0] MultLoop_acc_88_nl;
  wire[22:0] nl_MultLoop_acc_88_nl;
  wire[24:0] MultLoop_acc_93_nl;
  wire[25:0] nl_MultLoop_acc_93_nl;
  wire[23:0] MultLoop_acc_3763_nl;
  wire[25:0] nl_MultLoop_acc_3763_nl;
  wire[22:0] MultLoop_acc_92_nl;
  wire[23:0] nl_MultLoop_acc_92_nl;
  wire[21:0] MultLoop_acc_3766_nl;
  wire[23:0] nl_MultLoop_acc_3766_nl;
  wire[11:0] MultLoop_acc_4540_nl;
  wire[12:0] nl_MultLoop_acc_4540_nl;
  wire[17:0] MultLoop_acc_4542_nl;
  wire[18:0] nl_MultLoop_acc_4542_nl;
  wire[22:0] MultLoop_acc_3769_nl;
  wire[24:0] nl_MultLoop_acc_3769_nl;
  wire[19:0] MultLoop_acc_82_nl;
  wire[20:0] nl_MultLoop_acc_82_nl;
  wire[24:0] MultLoop_acc_83_nl;
  wire[26:0] nl_MultLoop_acc_83_nl;
  wire[17:0] MultLoop_acc_4545_nl;
  wire[18:0] nl_MultLoop_acc_4545_nl;
  wire[22:0] MultLoop_acc_3774_nl;
  wire[24:0] nl_MultLoop_acc_3774_nl;
  wire[18:0] MultLoop_acc_4546_nl;
  wire[19:0] nl_MultLoop_acc_4546_nl;
  wire[18:0] MultLoop_acc_4657_nl;
  wire[19:0] nl_MultLoop_acc_4657_nl;
  wire[22:0] MultLoop_acc_72_nl;
  wire[23:0] nl_MultLoop_acc_72_nl;
  wire[20:0] MultLoop_acc_3779_nl;
  wire[21:0] nl_MultLoop_acc_3779_nl;
  wire[21:0] MultLoop_acc_1094_nl;
  wire[22:0] nl_MultLoop_acc_1094_nl;
  wire[17:0] MultLoop_acc_3781_nl;
  wire[18:0] nl_MultLoop_acc_3781_nl;
  wire[13:0] MultLoop_acc_4548_nl;
  wire[14:0] nl_MultLoop_acc_4548_nl;
  wire[17:0] MultLoop_acc_4550_nl;
  wire[18:0] nl_MultLoop_acc_4550_nl;
  wire[19:0] MultLoop_acc_3783_nl;
  wire[20:0] nl_MultLoop_acc_3783_nl;
  wire[17:0] MultLoop_acc_4552_nl;
  wire[18:0] nl_MultLoop_acc_4552_nl;
  wire[23:0] MultLoop_acc_3786_nl;
  wire[24:0] nl_MultLoop_acc_3786_nl;
  wire[20:0] MultLoop_acc_3785_nl;
  wire[21:0] nl_MultLoop_acc_3785_nl;
  wire[10:0] MultLoop_acc_4551_nl;
  wire[11:0] nl_MultLoop_acc_4551_nl;
  wire[24:0] MultLoop_acc_1096_nl;
  wire[25:0] nl_MultLoop_acc_1096_nl;
  wire[17:0] MultLoop_acc_3792_nl;
  wire[18:0] nl_MultLoop_acc_3792_nl;
  wire[17:0] MultLoop_acc_4554_nl;
  wire[18:0] nl_MultLoop_acc_4554_nl;
  wire[21:0] MultLoop_acc_3788_nl;
  wire[22:0] nl_MultLoop_acc_3788_nl;
  wire[23:0] MultLoop_acc_51_nl;
  wire[25:0] nl_MultLoop_acc_51_nl;
  wire[13:0] MultLoop_acc_4555_nl;
  wire[14:0] nl_MultLoop_acc_4555_nl;
  wire[15:0] MultLoop_49_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_49_MultLoop_acc_3_nl;
  wire[17:0] MultLoop_acc_49_nl;
  wire[18:0] nl_MultLoop_acc_49_nl;
  wire[22:0] MultLoop_acc_78_nl;
  wire[23:0] nl_MultLoop_acc_78_nl;
  wire[20:0] MultLoop_acc_70_nl;
  wire[21:0] nl_MultLoop_acc_70_nl;
  wire[21:0] MultLoop_acc_58_nl;
  wire[22:0] nl_MultLoop_acc_58_nl;
  wire[19:0] MultLoop_acc_3738_nl;
  wire[20:0] nl_MultLoop_acc_3738_nl;
  wire[14:0] MultLoop_acc_4556_nl;
  wire[15:0] nl_MultLoop_acc_4556_nl;
  wire[17:0] MultLoop_acc_1795_nl;
  wire[19:0] nl_MultLoop_acc_1795_nl;
  wire[18:0] MultLoop_acc_3958_nl;
  wire[19:0] nl_MultLoop_acc_3958_nl;
  wire[22:0] MultLoop_acc_1749_nl;
  wire[24:0] nl_MultLoop_acc_1749_nl;
  wire[18:0] MultLoop_acc_3959_nl;
  wire[19:0] nl_MultLoop_acc_3959_nl;
  wire[21:0] MultLoop_acc_1750_nl;
  wire[22:0] nl_MultLoop_acc_1750_nl;
  wire[26:0] MultLoop_acc_1004_nl;
  wire[27:0] nl_MultLoop_acc_1004_nl;
  wire[24:0] MultLoop_acc_1752_nl;
  wire[25:0] nl_MultLoop_acc_1752_nl;
  wire[18:0] MultLoop_acc_3960_nl;
  wire[19:0] nl_MultLoop_acc_3960_nl;
  wire[18:0] MultLoop_acc_4596_nl;
  wire[19:0] nl_MultLoop_acc_4596_nl;
  wire[18:0] MultLoop_acc_1430_nl;
  wire[19:0] nl_MultLoop_acc_1430_nl;
  wire[18:0] MultLoop_acc_4595_nl;
  wire[19:0] nl_MultLoop_acc_4595_nl;
  wire[19:0] MultLoop_acc_3957_nl;
  wire[20:0] nl_MultLoop_acc_3957_nl;
  wire[17:0] MultLoop_acc_3956_nl;
  wire[18:0] nl_MultLoop_acc_3956_nl;
  wire[23:0] MultLoop_acc_1422_nl;
  wire[24:0] nl_MultLoop_acc_1422_nl;
  wire[19:0] MultLoop_acc_1747_nl;
  wire[20:0] nl_MultLoop_acc_1747_nl;
  wire[17:0] MultLoop_acc_1746_nl;
  wire[18:0] nl_MultLoop_acc_1746_nl;
  wire[21:0] MultLoop_acc_1042_nl;
  wire[22:0] nl_MultLoop_acc_1042_nl;
  wire[19:0] MultLoop_acc_1696_nl;
  wire[20:0] nl_MultLoop_acc_1696_nl;
  wire[17:0] MultLoop_acc_1695_nl;
  wire[18:0] nl_MultLoop_acc_1695_nl;
  wire[18:0] MultLoop_acc_1431_nl;
  wire[19:0] nl_MultLoop_acc_1431_nl;
  wire[17:0] MultLoop_acc_3963_nl;
  wire[18:0] nl_MultLoop_acc_3963_nl;
  wire[21:0] MultLoop_acc_1698_nl;
  wire[22:0] nl_MultLoop_acc_1698_nl;
  wire[21:0] MultLoop_acc_1002_nl;
  wire[22:0] nl_MultLoop_acc_1002_nl;
  wire[9:0] MultLoop_acc_1756_nl;
  wire[10:0] nl_MultLoop_acc_1756_nl;
  wire[20:0] MultLoop_acc_1423_nl;
  wire[21:0] nl_MultLoop_acc_1423_nl;
  wire[17:0] MultLoop_acc_1701_nl;
  wire[18:0] nl_MultLoop_acc_1701_nl;
  wire[14:0] MultLoop_acc_3964_nl;
  wire[15:0] nl_MultLoop_acc_3964_nl;
  wire[19:0] MultLoop_acc_4597_nl;
  wire[20:0] nl_MultLoop_acc_4597_nl;
  wire[17:0] MultLoop_acc_3966_nl;
  wire[18:0] nl_MultLoop_acc_3966_nl;
  wire[22:0] MultLoop_acc_1706_nl;
  wire[24:0] nl_MultLoop_acc_1706_nl;
  wire[20:0] MultLoop_acc_1429_nl;
  wire[21:0] nl_MultLoop_acc_1429_nl;
  wire[18:0] MultLoop_acc_1707_nl;
  wire[19:0] nl_MultLoop_acc_1707_nl;
  wire[22:0] MultLoop_acc_1427_nl;
  wire[23:0] nl_MultLoop_acc_1427_nl;
  wire[20:0] MultLoop_acc_1709_nl;
  wire[21:0] nl_MultLoop_acc_1709_nl;
  wire[19:0] MultLoop_acc_1418_nl;
  wire[20:0] nl_MultLoop_acc_1418_nl;
  wire[17:0] MultLoop_acc_1703_nl;
  wire[18:0] nl_MultLoop_acc_1703_nl;
  wire[24:0] MultLoop_acc_1027_nl;
  wire[26:0] nl_MultLoop_acc_1027_nl;
  wire[20:0] MultLoop_acc_1426_nl;
  wire[21:0] nl_MultLoop_acc_1426_nl;
  wire[17:0] MultLoop_acc_1712_nl;
  wire[18:0] nl_MultLoop_acc_1712_nl;
  wire[21:0] MultLoop_acc_1424_nl;
  wire[22:0] nl_MultLoop_acc_1424_nl;
  wire[17:0] MultLoop_acc_1714_nl;
  wire[18:0] nl_MultLoop_acc_1714_nl;
  wire[12:0] MultLoop_acc_3968_nl;
  wire[13:0] nl_MultLoop_acc_3968_nl;
  wire[22:0] MultLoop_acc_1022_nl;
  wire[23:0] nl_MultLoop_acc_1022_nl;
  wire[14:0] MultLoop_acc_3969_nl;
  wire[15:0] nl_MultLoop_acc_3969_nl;
  wire[24:0] MultLoop_acc_1020_nl;
  wire[26:0] nl_MultLoop_acc_1020_nl;
  wire[12:0] MultLoop_acc_3970_nl;
  wire[13:0] nl_MultLoop_acc_3970_nl;
  wire[21:0] MultLoop_acc_1419_nl;
  wire[22:0] nl_MultLoop_acc_1419_nl;
  wire[18:0] MultLoop_acc_1719_nl;
  wire[19:0] nl_MultLoop_acc_1719_nl;
  wire[24:0] MultLoop_acc_1003_nl;
  wire[25:0] nl_MultLoop_acc_1003_nl;
  wire[22:0] MultLoop_acc_1721_nl;
  wire[23:0] nl_MultLoop_acc_1721_nl;
  wire[20:0] MultLoop_acc_4598_nl;
  wire[21:0] nl_MultLoop_acc_4598_nl;
  wire[22:0] MultLoop_acc_1038_nl;
  wire[24:0] nl_MultLoop_acc_1038_nl;
  wire[20:0] MultLoop_acc_1013_nl;
  wire[21:0] nl_MultLoop_acc_1013_nl;
  wire[18:0] MultLoop_acc_1693_nl;
  wire[19:0] nl_MultLoop_acc_1693_nl;
  wire[13:0] MultLoop_acc_3972_nl;
  wire[14:0] nl_MultLoop_acc_3972_nl;
  wire[25:0] MultLoop_acc_1037_nl;
  wire[26:0] nl_MultLoop_acc_1037_nl;
  wire[21:0] MultLoop_acc_1724_nl;
  wire[22:0] nl_MultLoop_acc_1724_nl;
  wire[18:0] MultLoop_acc_4599_nl;
  wire[19:0] nl_MultLoop_acc_4599_nl;
  wire[25:0] MultLoop_acc_1030_nl;
  wire[26:0] nl_MultLoop_acc_1030_nl;
  wire[21:0] MultLoop_acc_1726_nl;
  wire[22:0] nl_MultLoop_acc_1726_nl;
  wire[22:0] MultLoop_acc_1425_nl;
  wire[23:0] nl_MultLoop_acc_1425_nl;
  wire[20:0] MultLoop_acc_1728_nl;
  wire[21:0] nl_MultLoop_acc_1728_nl;
  wire[23:0] MultLoop_acc_1024_nl;
  wire[24:0] nl_MultLoop_acc_1024_nl;
  wire[21:0] MultLoop_acc_1729_nl;
  wire[22:0] nl_MultLoop_acc_1729_nl;
  wire[18:0] MultLoop_acc_3975_nl;
  wire[19:0] nl_MultLoop_acc_3975_nl;
  wire[21:0] MultLoop_acc_1736_nl;
  wire[22:0] nl_MultLoop_acc_1736_nl;
  wire[25:0] MultLoop_acc_1000_nl;
  wire[26:0] nl_MultLoop_acc_1000_nl;
  wire[24:0] MultLoop_acc_1738_nl;
  wire[26:0] nl_MultLoop_acc_1738_nl;
  wire[18:0] MultLoop_acc_3973_nl;
  wire[19:0] nl_MultLoop_acc_3973_nl;
  wire[24:0] MultLoop_acc_1011_nl;
  wire[25:0] nl_MultLoop_acc_1011_nl;
  wire[23:0] MultLoop_acc_1731_nl;
  wire[24:0] nl_MultLoop_acc_1731_nl;
  wire[22:0] MultLoop_acc_1008_nl;
  wire[23:0] nl_MultLoop_acc_1008_nl;
  wire[20:0] MultLoop_acc_1734_nl;
  wire[21:0] nl_MultLoop_acc_1734_nl;
  wire[17:0] MultLoop_acc_1733_nl;
  wire[18:0] nl_MultLoop_acc_1733_nl;
  wire[23:0] MultLoop_acc_4600_nl;
  wire[24:0] nl_MultLoop_acc_4600_nl;
  wire[24:0] MultLoop_acc_1001_nl;
  wire[25:0] nl_MultLoop_acc_1001_nl;
  wire[21:0] MultLoop_acc_1740_nl;
  wire[23:0] nl_MultLoop_acc_1740_nl;
  wire[22:0] MultLoop_acc_1417_nl;
  wire[23:0] nl_MultLoop_acc_1417_nl;
  wire[20:0] MultLoop_acc_1742_nl;
  wire[21:0] nl_MultLoop_acc_1742_nl;
  wire[22:0] MultLoop_acc_106_nl;
  wire[24:0] nl_MultLoop_acc_106_nl;
  wire[14:0] MultLoop_acc_4500_nl;
  wire[15:0] nl_MultLoop_acc_4500_nl;
  wire[25:0] MultLoop_acc_107_nl;
  wire[27:0] nl_MultLoop_acc_107_nl;
  wire[11:0] MultLoop_acc_4501_nl;
  wire[12:0] nl_MultLoop_acc_4501_nl;
  wire[25:0] MultLoop_acc_101_nl;
  wire[27:0] nl_MultLoop_acc_101_nl;
  wire[23:0] MultLoop_acc_1120_nl;
  wire[24:0] nl_MultLoop_acc_1120_nl;
  wire[20:0] MultLoop_acc_3677_nl;
  wire[21:0] nl_MultLoop_acc_3677_nl;
  wire[17:0] MultLoop_acc_3676_nl;
  wire[18:0] nl_MultLoop_acc_3676_nl;
  wire[23:0] MultLoop_acc_1117_nl;
  wire[24:0] nl_MultLoop_acc_1117_nl;
  wire[20:0] MultLoop_acc_3680_nl;
  wire[21:0] nl_MultLoop_acc_3680_nl;
  wire[17:0] MultLoop_acc_3679_nl;
  wire[18:0] nl_MultLoop_acc_3679_nl;
  wire[21:0] MultLoop_acc_1104_nl;
  wire[22:0] nl_MultLoop_acc_1104_nl;
  wire[17:0] MultLoop_acc_3682_nl;
  wire[18:0] nl_MultLoop_acc_3682_nl;
  wire[13:0] MultLoop_acc_4505_nl;
  wire[14:0] nl_MultLoop_acc_4505_nl;
  wire[16:0] MultLoop_100_MultLoop_acc_3_nl;
  wire[18:0] nl_MultLoop_100_MultLoop_acc_3_nl;
  wire[20:0] MultLoop_acc_1102_nl;
  wire[21:0] nl_MultLoop_acc_1102_nl;
  wire[17:0] MultLoop_acc_3687_nl;
  wire[18:0] nl_MultLoop_acc_3687_nl;
  wire[11:0] MultLoop_acc_4506_nl;
  wire[12:0] nl_MultLoop_acc_4506_nl;
  wire[20:0] MultLoop_acc_1103_nl;
  wire[21:0] nl_MultLoop_acc_1103_nl;
  wire[18:0] MultLoop_acc_3688_nl;
  wire[19:0] nl_MultLoop_acc_3688_nl;
  wire[19:0] MultLoop_acc_4653_nl;
  wire[20:0] nl_MultLoop_acc_4653_nl;
  wire[13:0] MultLoop_97_MultLoop_acc_3_nl;
  wire[14:0] nl_MultLoop_97_MultLoop_acc_3_nl;
  wire[18:0] MultLoop_acc_4696_nl;
  wire[19:0] nl_MultLoop_acc_4696_nl;
  wire[21:0] MultLoop_acc_100_nl;
  wire[22:0] nl_MultLoop_acc_100_nl;
  wire[15:0] MultLoop_acc_4507_nl;
  wire[16:0] nl_MultLoop_acc_4507_nl;
  wire[14:0] MultLoop_acc_3696_nl;
  wire[16:0] nl_MultLoop_acc_3696_nl;
  wire[20:0] MultLoop_acc_103_nl;
  wire[21:0] nl_MultLoop_acc_103_nl;
  wire[16:0] MultLoop_acc_4508_nl;
  wire[17:0] nl_MultLoop_acc_4508_nl;
  wire[21:0] MultLoop_acc_134_nl;
  wire[22:0] nl_MultLoop_acc_134_nl;
  wire[19:0] MultLoop_acc_3618_nl;
  wire[20:0] nl_MultLoop_acc_3618_nl;
  wire[14:0] MultLoop_acc_4509_nl;
  wire[15:0] nl_MultLoop_acc_4509_nl;
  wire[23:0] MultLoop_acc_130_nl;
  wire[24:0] nl_MultLoop_acc_130_nl;
  wire[22:0] MultLoop_acc_3621_nl;
  wire[23:0] nl_MultLoop_acc_3621_nl;
  wire[21:0] MultLoop_acc_1115_nl;
  wire[22:0] nl_MultLoop_acc_1115_nl;
  wire[18:0] MultLoop_acc_3622_nl;
  wire[19:0] nl_MultLoop_acc_3622_nl;
  wire[21:0] MultLoop_acc_1119_nl;
  wire[22:0] nl_MultLoop_acc_1119_nl;
  wire[20:0] MultLoop_acc_3625_nl;
  wire[21:0] nl_MultLoop_acc_3625_nl;
  wire[17:0] MultLoop_acc_3624_nl;
  wire[18:0] nl_MultLoop_acc_3624_nl;
  wire[17:0] MultLoop_acc_4511_nl;
  wire[18:0] nl_MultLoop_acc_4511_nl;
  wire[22:0] MultLoop_acc_3628_nl;
  wire[24:0] nl_MultLoop_acc_3628_nl;
  wire[11:0] MultLoop_acc_4510_nl;
  wire[12:0] nl_MultLoop_acc_4510_nl;
  wire[23:0] MultLoop_acc_120_nl;
  wire[24:0] nl_MultLoop_acc_120_nl;
  wire[22:0] MultLoop_acc_3623_nl;
  wire[23:0] nl_MultLoop_acc_3623_nl;
  wire[18:0] MultLoop_acc_1105_nl;
  wire[19:0] nl_MultLoop_acc_1105_nl;
  wire[20:0] MultLoop_acc_1112_nl;
  wire[21:0] nl_MultLoop_acc_1112_nl;
  wire[19:0] MultLoop_acc_129_nl;
  wire[20:0] nl_MultLoop_acc_129_nl;
  wire[18:0] MultLoop_acc_3630_nl;
  wire[19:0] nl_MultLoop_acc_3630_nl;
  wire[14:0] MultLoop_acc_4512_nl;
  wire[15:0] nl_MultLoop_acc_4512_nl;
  wire[19:0] MultLoop_acc_1114_nl;
  wire[20:0] nl_MultLoop_acc_1114_nl;
  wire[17:0] MultLoop_acc_3631_nl;
  wire[18:0] nl_MultLoop_acc_3631_nl;
  wire[20:0] MultLoop_acc_118_nl;
  wire[21:0] nl_MultLoop_acc_118_nl;
  wire[18:0] MultLoop_acc_3633_nl;
  wire[19:0] nl_MultLoop_acc_3633_nl;
  wire[18:0] MultLoop_acc_4514_nl;
  wire[19:0] nl_MultLoop_acc_4514_nl;
  wire[21:0] MultLoop_acc_3635_nl;
  wire[22:0] nl_MultLoop_acc_3635_nl;
  wire[24:0] MultLoop_acc_143_nl;
  wire[25:0] nl_MultLoop_acc_143_nl;
  wire[22:0] MultLoop_acc_3637_nl;
  wire[23:0] nl_MultLoop_acc_3637_nl;
  wire[23:0] MultLoop_acc_1118_nl;
  wire[24:0] nl_MultLoop_acc_1118_nl;
  wire[20:0] MultLoop_acc_3640_nl;
  wire[21:0] nl_MultLoop_acc_3640_nl;
  wire[17:0] MultLoop_acc_3639_nl;
  wire[18:0] nl_MultLoop_acc_3639_nl;
  wire[17:0] MultLoop_acc_110_nl;
  wire[18:0] nl_MultLoop_acc_110_nl;
  wire[17:0] MultLoop_acc_4517_nl;
  wire[18:0] nl_MultLoop_acc_4517_nl;
  wire[19:0] MultLoop_acc_4686_nl;
  wire[20:0] nl_MultLoop_acc_4686_nl;
  wire[17:0] MultLoop_acc_4519_nl;
  wire[18:0] nl_MultLoop_acc_4519_nl;
  wire[22:0] MultLoop_acc_3646_nl;
  wire[24:0] nl_MultLoop_acc_3646_nl;
  wire[21:0] MultLoop_acc_132_nl;
  wire[22:0] nl_MultLoop_acc_132_nl;
  wire[18:0] MultLoop_acc_3648_nl;
  wire[19:0] nl_MultLoop_acc_3648_nl;
  wire[12:0] MultLoop_acc_4520_nl;
  wire[13:0] nl_MultLoop_acc_4520_nl;
  wire[19:0] MultLoop_acc_1116_nl;
  wire[20:0] nl_MultLoop_acc_1116_nl;
  wire[17:0] MultLoop_acc_3649_nl;
  wire[18:0] nl_MultLoop_acc_3649_nl;
  wire[25:0] MultLoop_acc_126_nl;
  wire[27:0] nl_MultLoop_acc_126_nl;
  wire[17:0] MultLoop_acc_4523_nl;
  wire[18:0] nl_MultLoop_acc_4523_nl;
  wire[19:0] MultLoop_acc_3654_nl;
  wire[20:0] nl_MultLoop_acc_3654_nl;
  wire[23:0] MultLoop_acc_1110_nl;
  wire[24:0] nl_MultLoop_acc_1110_nl;
  wire[19:0] MultLoop_acc_3657_nl;
  wire[21:0] nl_MultLoop_acc_3657_nl;
  wire[18:0] MultLoop_acc_1111_nl;
  wire[19:0] nl_MultLoop_acc_1111_nl;
  wire[18:0] MultLoop_acc_4525_nl;
  wire[19:0] nl_MultLoop_acc_4525_nl;
  wire[23:0] MultLoop_acc_115_nl;
  wire[24:0] nl_MultLoop_acc_115_nl;
  wire[21:0] MultLoop_acc_3660_nl;
  wire[22:0] nl_MultLoop_acc_3660_nl;
  wire[19:0] MultLoop_acc_3659_nl;
  wire[20:0] nl_MultLoop_acc_3659_nl;
  wire[18:0] MultLoop_acc_4654_nl;
  wire[19:0] nl_MultLoop_acc_4654_nl;
  wire[17:0] MultLoop_acc_4527_nl;
  wire[18:0] nl_MultLoop_acc_4527_nl;
  wire[23:0] MultLoop_acc_3665_nl;
  wire[25:0] nl_MultLoop_acc_3665_nl;
  wire[10:0] MultLoop_acc_4526_nl;
  wire[11:0] nl_MultLoop_acc_4526_nl;
  wire[23:0] MultLoop_acc_1107_nl;
  wire[24:0] nl_MultLoop_acc_1107_nl;
  wire[21:0] MultLoop_acc_3667_nl;
  wire[22:0] nl_MultLoop_acc_3667_nl;
  wire[22:0] MultLoop_acc_965_nl;
  wire[23:0] nl_MultLoop_acc_965_nl;
  wire[19:0] MultLoop_acc_1839_nl;
  wire[20:0] nl_MultLoop_acc_1839_nl;
  wire[17:0] MultLoop_acc_1838_nl;
  wire[18:0] nl_MultLoop_acc_1838_nl;
  wire[22:0] MultLoop_acc_1405_nl;
  wire[23:0] nl_MultLoop_acc_1405_nl;
  wire[17:0] MultLoop_acc_1841_nl;
  wire[18:0] nl_MultLoop_acc_1841_nl;
  wire[11:0] MultLoop_acc_3977_nl;
  wire[12:0] nl_MultLoop_acc_3977_nl;
  wire[25:0] MultLoop_acc_963_nl;
  wire[26:0] nl_MultLoop_acc_963_nl;
  wire[24:0] MultLoop_acc_1843_nl;
  wire[25:0] nl_MultLoop_acc_1843_nl;
  wire[21:0] MultLoop_acc_1403_nl;
  wire[22:0] nl_MultLoop_acc_1403_nl;
  wire[23:0] MultLoop_acc_1404_nl;
  wire[24:0] nl_MultLoop_acc_1404_nl;
  wire[21:0] MultLoop_acc_1846_nl;
  wire[23:0] nl_MultLoop_acc_1846_nl;
  wire[18:0] MultLoop_acc_4664_nl;
  wire[19:0] nl_MultLoop_acc_4664_nl;
  wire[25:0] MultLoop_acc_954_nl;
  wire[27:0] nl_MultLoop_acc_954_nl;
  wire[20:0] MultLoop_acc_3983_nl;
  wire[21:0] nl_MultLoop_acc_3983_nl;
  wire[17:0] MultLoop_acc_3982_nl;
  wire[18:0] nl_MultLoop_acc_3982_nl;
  wire[19:0] MultLoop_acc_1856_nl;
  wire[20:0] nl_MultLoop_acc_1856_nl;
  wire[10:0] MultLoop_acc_3981_nl;
  wire[11:0] nl_MultLoop_acc_3981_nl;
  wire[18:0] MultLoop_acc_4601_nl;
  wire[19:0] nl_MultLoop_acc_4601_nl;
  wire[25:0] MultLoop_acc_984_nl;
  wire[26:0] nl_MultLoop_acc_984_nl;
  wire[21:0] MultLoop_acc_1861_nl;
  wire[22:0] nl_MultLoop_acc_1861_nl;
  wire[19:0] MultLoop_acc_1860_nl;
  wire[20:0] nl_MultLoop_acc_1860_nl;
  wire[11:0] MultLoop_acc_3984_nl;
  wire[12:0] nl_MultLoop_acc_3984_nl;
  wire[17:0] MultLoop_acc_3980_nl;
  wire[18:0] nl_MultLoop_acc_3980_nl;
  wire[22:0] MultLoop_acc_1854_nl;
  wire[23:0] nl_MultLoop_acc_1854_nl;
  wire[19:0] MultLoop_acc_1853_nl;
  wire[20:0] nl_MultLoop_acc_1853_nl;
  wire[19:0] MultLoop_acc_953_nl;
  wire[20:0] nl_MultLoop_acc_953_nl;
  wire[25:0] MultLoop_acc_982_nl;
  wire[26:0] nl_MultLoop_acc_982_nl;
  wire[22:0] MultLoop_acc_1864_nl;
  wire[23:0] nl_MultLoop_acc_1864_nl;
  wire[19:0] MultLoop_acc_1863_nl;
  wire[20:0] nl_MultLoop_acc_1863_nl;
  wire[23:0] MultLoop_acc_4665_nl;
  wire[24:0] nl_MultLoop_acc_4665_nl;
  wire[22:0] MultLoop_acc_1410_nl;
  wire[23:0] nl_MultLoop_acc_1410_nl;
  wire[19:0] MultLoop_acc_1869_nl;
  wire[21:0] nl_MultLoop_acc_1869_nl;
  wire[25:0] MultLoop_acc_974_nl;
  wire[27:0] nl_MultLoop_acc_974_nl;
  wire[16:0] MultLoop_acc_1904_nl;
  wire[19:0] nl_MultLoop_acc_1904_nl;
  wire[24:0] MultLoop_acc_951_nl;
  wire[25:0] nl_MultLoop_acc_951_nl;
  wire[12:0] MultLoop_acc_3991_nl;
  wire[13:0] nl_MultLoop_acc_3991_nl;
  wire[22:0] MultLoop_acc_991_nl;
  wire[23:0] nl_MultLoop_acc_991_nl;
  wire[17:0] MultLoop_acc_970_nl;
  wire[18:0] nl_MultLoop_acc_970_nl;
  wire[20:0] MultLoop_acc_1409_nl;
  wire[21:0] nl_MultLoop_acc_1409_nl;
  wire[17:0] MultLoop_acc_1807_nl;
  wire[18:0] nl_MultLoop_acc_1807_nl;
  wire[22:0] MultLoop_acc_968_nl;
  wire[23:0] nl_MultLoop_acc_968_nl;
  wire[19:0] MultLoop_acc_1808_nl;
  wire[20:0] nl_MultLoop_acc_1808_nl;
  wire[24:0] MultLoop_acc_1406_nl;
  wire[25:0] nl_MultLoop_acc_1406_nl;
  wire[21:0] MultLoop_acc_1875_nl;
  wire[23:0] nl_MultLoop_acc_1875_nl;
  wire[24:0] MultLoop_acc_1402_nl;
  wire[25:0] nl_MultLoop_acc_1402_nl;
  wire[19:0] MultLoop_acc_1878_nl;
  wire[21:0] nl_MultLoop_acc_1878_nl;
  wire[10:0] MultLoop_acc_3990_nl;
  wire[11:0] nl_MultLoop_acc_3990_nl;
  wire[24:0] MultLoop_acc_988_nl;
  wire[25:0] nl_MultLoop_acc_988_nl;
  wire[22:0] MultLoop_acc_1809_nl;
  wire[23:0] nl_MultLoop_acc_1809_nl;
  wire[22:0] MultLoop_acc_990_nl;
  wire[24:0] nl_MultLoop_acc_990_nl;
  wire[14:0] MultLoop_acc_3994_nl;
  wire[15:0] nl_MultLoop_acc_3994_nl;
  wire[20:0] MultLoop_acc_4602_nl;
  wire[21:0] nl_MultLoop_acc_4602_nl;
  wire[21:0] MultLoop_acc_976_nl;
  wire[22:0] nl_MultLoop_acc_976_nl;
  wire[15:0] MultLoop_acc_3995_nl;
  wire[16:0] nl_MultLoop_acc_3995_nl;
  wire[17:0] MultLoop_acc_3997_nl;
  wire[18:0] nl_MultLoop_acc_3997_nl;
  wire[22:0] MultLoop_acc_1814_nl;
  wire[23:0] nl_MultLoop_acc_1814_nl;
  wire[11:0] MultLoop_acc_3996_nl;
  wire[12:0] nl_MultLoop_acc_3996_nl;
  wire[22:0] MultLoop_acc_4666_nl;
  wire[23:0] nl_MultLoop_acc_4666_nl;
  wire[21:0] MultLoop_acc_994_nl;
  wire[22:0] nl_MultLoop_acc_994_nl;
  wire[20:0] MultLoop_acc_1820_nl;
  wire[22:0] nl_MultLoop_acc_1820_nl;
  wire[10:0] MultLoop_acc_3999_nl;
  wire[11:0] nl_MultLoop_acc_3999_nl;
  wire[22:0] MultLoop_acc_1416_nl;
  wire[23:0] nl_MultLoop_acc_1416_nl;
  wire[19:0] MultLoop_acc_1823_nl;
  wire[20:0] nl_MultLoop_acc_1823_nl;
  wire[17:0] MultLoop_acc_4002_nl;
  wire[18:0] nl_MultLoop_acc_4002_nl;
  wire[22:0] MultLoop_acc_1825_nl;
  wire[23:0] nl_MultLoop_acc_1825_nl;
  wire[14:0] MultLoop_961_MultLoop_acc_3_nl;
  wire[15:0] nl_MultLoop_961_MultLoop_acc_3_nl;
  wire[19:0] MultLoop_acc_950_nl;
  wire[20:0] nl_MultLoop_acc_950_nl;
  wire[17:0] MultLoop_acc_1817_nl;
  wire[18:0] nl_MultLoop_acc_1817_nl;
  wire[22:0] MultLoop_acc_985_nl;
  wire[23:0] nl_MultLoop_acc_985_nl;
  wire[25:0] MultLoop_acc_972_nl;
  wire[26:0] nl_MultLoop_acc_972_nl;
  wire[23:0] MultLoop_acc_1833_nl;
  wire[24:0] nl_MultLoop_acc_1833_nl;
  wire[23:0] MultLoop_acc_1415_nl;
  wire[24:0] nl_MultLoop_acc_1415_nl;
  wire[22:0] MultLoop_acc_1828_nl;
  wire[24:0] nl_MultLoop_acc_1828_nl;
  wire[17:0] MultLoop_acc_1826_nl;
  wire[18:0] nl_MultLoop_acc_1826_nl;
  wire[21:0] MultLoop_acc_1412_nl;
  wire[22:0] nl_MultLoop_acc_1412_nl;
  wire[17:0] MultLoop_acc_1830_nl;
  wire[18:0] nl_MultLoop_acc_1830_nl;
  wire[13:0] MultLoop_acc_4003_nl;
  wire[14:0] nl_MultLoop_acc_4003_nl;
  wire[21:0] MultLoop_acc_1408_nl;
  wire[22:0] nl_MultLoop_acc_1408_nl;
  wire[18:0] MultLoop_acc_1831_nl;
  wire[19:0] nl_MultLoop_acc_1831_nl;
  wire[20:0] MultLoop_acc_1407_nl;
  wire[21:0] nl_MultLoop_acc_1407_nl;
  wire[17:0] MultLoop_acc_1834_nl;
  wire[18:0] nl_MultLoop_acc_1834_nl;
  wire[25:0] MultLoop_acc_964_nl;
  wire[26:0] nl_MultLoop_acc_964_nl;
  wire[23:0] MultLoop_acc_1836_nl;
  wire[25:0] nl_MultLoop_acc_1836_nl;
  wire[17:0] MultLoop_acc_3609_nl;
  wire[19:0] nl_MultLoop_acc_3609_nl;
  wire[20:0] MultLoop_acc_1137_nl;
  wire[21:0] nl_MultLoop_acc_1137_nl;
  wire[18:0] MultLoop_acc_3560_nl;
  wire[19:0] nl_MultLoop_acc_3560_nl;
  wire[18:0] MultLoop_acc_4473_nl;
  wire[19:0] nl_MultLoop_acc_4473_nl;
  wire[19:0] MultLoop_acc_4695_nl;
  wire[20:0] nl_MultLoop_acc_4695_nl;
  wire[23:0] MultLoop_acc_173_nl;
  wire[24:0] nl_MultLoop_acc_173_nl;
  wire[22:0] MultLoop_acc_3563_nl;
  wire[23:0] nl_MultLoop_acc_3563_nl;
  wire[24:0] MultLoop_acc_1132_nl;
  wire[25:0] nl_MultLoop_acc_1132_nl;
  wire[22:0] MultLoop_acc_3565_nl;
  wire[23:0] nl_MultLoop_acc_3565_nl;
  wire[20:0] MultLoop_acc_1122_nl;
  wire[21:0] nl_MultLoop_acc_1122_nl;
  wire[18:0] MultLoop_acc_3552_nl;
  wire[19:0] nl_MultLoop_acc_3552_nl;
  wire[21:0] MultLoop_acc_1140_nl;
  wire[22:0] nl_MultLoop_acc_1140_nl;
  wire[18:0] MultLoop_acc_3557_nl;
  wire[19:0] nl_MultLoop_acc_3557_nl;
  wire[22:0] MultLoop_acc_1138_nl;
  wire[23:0] nl_MultLoop_acc_1138_nl;
  wire[19:0] MultLoop_acc_3559_nl;
  wire[20:0] nl_MultLoop_acc_3559_nl;
  wire[17:0] MultLoop_acc_3558_nl;
  wire[18:0] nl_MultLoop_acc_3558_nl;
  wire[21:0] MultLoop_acc_1123_nl;
  wire[22:0] nl_MultLoop_acc_1123_nl;
  wire[17:0] MultLoop_acc_3554_nl;
  wire[18:0] nl_MultLoop_acc_3554_nl;
  wire[12:0] MultLoop_acc_4472_nl;
  wire[13:0] nl_MultLoop_acc_4472_nl;
  wire[20:0] MultLoop_acc_4651_nl;
  wire[21:0] nl_MultLoop_acc_4651_nl;
  wire[22:0] MultLoop_acc_1125_nl;
  wire[23:0] nl_MultLoop_acc_1125_nl;
  wire[19:0] MultLoop_acc_3567_nl;
  wire[20:0] nl_MultLoop_acc_3567_nl;
  wire[18:0] MultLoop_acc_4474_nl;
  wire[19:0] nl_MultLoop_acc_4474_nl;
  wire[17:0] MultLoop_acc_188_nl;
  wire[18:0] nl_MultLoop_acc_188_nl;
  wire[17:0] MultLoop_acc_4476_nl;
  wire[18:0] nl_MultLoop_acc_4476_nl;
  wire[21:0] MultLoop_acc_3504_nl;
  wire[22:0] nl_MultLoop_acc_3504_nl;
  wire[18:0] MultLoop_acc_1133_nl;
  wire[19:0] nl_MultLoop_acc_1133_nl;
  wire[20:0] MultLoop_acc_1131_nl;
  wire[21:0] nl_MultLoop_acc_1131_nl;
  wire[17:0] MultLoop_acc_3506_nl;
  wire[18:0] nl_MultLoop_acc_3506_nl;
  wire[19:0] MultLoop_acc_1127_nl;
  wire[20:0] nl_MultLoop_acc_1127_nl;
  wire[17:0] MultLoop_acc_3507_nl;
  wire[18:0] nl_MultLoop_acc_3507_nl;
  wire[17:0] MultLoop_acc_4479_nl;
  wire[18:0] nl_MultLoop_acc_4479_nl;
  wire[21:0] MultLoop_acc_3509_nl;
  wire[22:0] nl_MultLoop_acc_3509_nl;
  wire[12:0] MultLoop_acc_4478_nl;
  wire[13:0] nl_MultLoop_acc_4478_nl;
  wire[22:0] MultLoop_acc_153_nl;
  wire[23:0] nl_MultLoop_acc_153_nl;
  wire[14:0] MultLoop_acc_4480_nl;
  wire[15:0] nl_MultLoop_acc_4480_nl;
  wire[22:0] MultLoop_acc_1141_nl;
  wire[23:0] nl_MultLoop_acc_1141_nl;
  wire[23:0] MultLoop_acc_183_nl;
  wire[24:0] nl_MultLoop_acc_183_nl;
  wire[12:0] MultLoop_acc_3571_nl;
  wire[13:0] nl_MultLoop_acc_3571_nl;
  wire[20:0] MultLoop_acc_166_nl;
  wire[21:0] nl_MultLoop_acc_166_nl;
  wire[16:0] MultLoop_acc_4481_nl;
  wire[17:0] nl_MultLoop_acc_4481_nl;
  wire[9:0] MultLoop_acc_4482_nl;
  wire[10:0] nl_MultLoop_acc_4482_nl;
  wire[17:0] MultLoop_acc_175_nl;
  wire[18:0] nl_MultLoop_acc_175_nl;
  wire[19:0] MultLoop_acc_4685_nl;
  wire[20:0] nl_MultLoop_acc_4685_nl;
  wire[19:0] MultLoop_acc_1126_nl;
  wire[20:0] nl_MultLoop_acc_1126_nl;
  wire[17:0] MultLoop_acc_3514_nl;
  wire[18:0] nl_MultLoop_acc_3514_nl;
  wire[14:0] MultLoop_acc_3577_nl;
  wire[15:0] nl_MultLoop_acc_3577_nl;
  wire[19:0] MultLoop_acc_4652_nl;
  wire[20:0] nl_MultLoop_acc_4652_nl;
  wire[17:0] MultLoop_acc_4485_nl;
  wire[18:0] nl_MultLoop_acc_4485_nl;
  wire[22:0] MultLoop_acc_3517_nl;
  wire[24:0] nl_MultLoop_acc_3517_nl;
  wire[25:0] MultLoop_acc_192_nl;
  wire[26:0] nl_MultLoop_acc_192_nl;
  wire[21:0] MultLoop_acc_3519_nl;
  wire[22:0] nl_MultLoop_acc_3519_nl;
  wire[17:0] MultLoop_acc_4487_nl;
  wire[18:0] nl_MultLoop_acc_4487_nl;
  wire[24:0] MultLoop_acc_3523_nl;
  wire[26:0] nl_MultLoop_acc_3523_nl;
  wire[17:0] MultLoop_acc_4489_nl;
  wire[18:0] nl_MultLoop_acc_4489_nl;
  wire[23:0] MultLoop_acc_3526_nl;
  wire[24:0] nl_MultLoop_acc_3526_nl;
  wire[20:0] MultLoop_acc_3525_nl;
  wire[21:0] nl_MultLoop_acc_3525_nl;
  wire[17:0] MultLoop_acc_4491_nl;
  wire[18:0] nl_MultLoop_acc_4491_nl;
  wire[22:0] MultLoop_acc_3530_nl;
  wire[23:0] nl_MultLoop_acc_3530_nl;
  wire[19:0] MultLoop_acc_3529_nl;
  wire[20:0] nl_MultLoop_acc_3529_nl;
  wire[17:0] MultLoop_acc_3528_nl;
  wire[18:0] nl_MultLoop_acc_3528_nl;
  wire[18:0] MultLoop_acc_4693_nl;
  wire[19:0] nl_MultLoop_acc_4693_nl;
  wire[22:0] MultLoop_acc_1135_nl;
  wire[23:0] nl_MultLoop_acc_1135_nl;
  wire[20:0] MultLoop_acc_3535_nl;
  wire[21:0] nl_MultLoop_acc_3535_nl;
  wire[17:0] MultLoop_acc_3534_nl;
  wire[18:0] nl_MultLoop_acc_3534_nl;
  wire[17:0] MultLoop_acc_4496_nl;
  wire[18:0] nl_MultLoop_acc_4496_nl;
  wire[22:0] MultLoop_acc_3546_nl;
  wire[23:0] nl_MultLoop_acc_3546_nl;
  wire[17:0] MultLoop_acc_4498_nl;
  wire[18:0] nl_MultLoop_acc_4498_nl;
  wire[19:0] MultLoop_acc_3548_nl;
  wire[20:0] nl_MultLoop_acc_3548_nl;
  wire[19:0] MultLoop_acc_1134_nl;
  wire[20:0] nl_MultLoop_acc_1134_nl;
  wire[17:0] MultLoop_acc_3536_nl;
  wire[18:0] nl_MultLoop_acc_3536_nl;
  wire[22:0] MultLoop_acc_174_nl;
  wire[23:0] nl_MultLoop_acc_174_nl;
  wire[21:0] MultLoop_acc_3539_nl;
  wire[22:0] nl_MultLoop_acc_3539_nl;
  wire[21:0] MultLoop_acc_1129_nl;
  wire[22:0] nl_MultLoop_acc_1129_nl;
  wire[20:0] MultLoop_acc_3541_nl;
  wire[21:0] nl_MultLoop_acc_3541_nl;
  wire[17:0] MultLoop_acc_3540_nl;
  wire[18:0] nl_MultLoop_acc_3540_nl;
  wire[23:0] MultLoop_acc_1130_nl;
  wire[24:0] nl_MultLoop_acc_1130_nl;
  wire[20:0] MultLoop_acc_3544_nl;
  wire[21:0] nl_MultLoop_acc_3544_nl;
  wire[17:0] MultLoop_acc_3543_nl;
  wire[18:0] nl_MultLoop_acc_3543_nl;
  wire[22:0] MultLoop_acc_154_nl;
  wire[23:0] nl_MultLoop_acc_154_nl;
  wire[20:0] MultLoop_acc_3550_nl;
  wire[21:0] nl_MultLoop_acc_3550_nl;
  wire[20:0] MultLoop_acc_1124_nl;
  wire[21:0] nl_MultLoop_acc_1124_nl;
  wire[23:0] MultLoop_acc_1401_nl;
  wire[24:0] nl_MultLoop_acc_1401_nl;
  wire[20:0] MultLoop_acc_1992_nl;
  wire[22:0] nl_MultLoop_acc_1992_nl;
  wire[18:0] MultLoop_acc_4603_nl;
  wire[19:0] nl_MultLoop_acc_4603_nl;
  wire[19:0] MultLoop_acc_1385_nl;
  wire[20:0] nl_MultLoop_acc_1385_nl;
  wire[17:0] MultLoop_acc_1983_nl;
  wire[18:0] nl_MultLoop_acc_1983_nl;
  wire[17:0] MultLoop_acc_4005_nl;
  wire[18:0] nl_MultLoop_acc_4005_nl;
  wire[23:0] MultLoop_acc_1986_nl;
  wire[25:0] nl_MultLoop_acc_1986_nl;
  wire[10:0] MultLoop_acc_4004_nl;
  wire[11:0] nl_MultLoop_acc_4004_nl;
  wire[19:0] MultLoop_acc_4007_nl;
  wire[20:0] nl_MultLoop_acc_4007_nl;
  wire[17:0] MultLoop_acc_4006_nl;
  wire[18:0] nl_MultLoop_acc_4006_nl;
  wire[17:0] MultLoop_acc_4010_nl;
  wire[18:0] nl_MultLoop_acc_4010_nl;
  wire[20:0] MultLoop_acc_1929_nl;
  wire[21:0] nl_MultLoop_acc_1929_nl;
  wire[12:0] MultLoop_acc_4009_nl;
  wire[13:0] nl_MultLoop_acc_4009_nl;
  wire[19:0] MultLoop_acc_927_nl;
  wire[20:0] nl_MultLoop_acc_927_nl;
  wire[18:0] MultLoop_acc_1927_nl;
  wire[19:0] nl_MultLoop_acc_1927_nl;
  wire[26:0] MultLoop_acc_933_nl;
  wire[28:0] nl_MultLoop_acc_933_nl;
  wire[10:0] MultLoop_acc_4012_nl;
  wire[11:0] nl_MultLoop_acc_4012_nl;
  wire[23:0] MultLoop_acc_920_nl;
  wire[25:0] nl_MultLoop_acc_920_nl;
  wire[13:0] MultLoop_acc_4013_nl;
  wire[14:0] nl_MultLoop_acc_4013_nl;
  wire[22:0] MultLoop_acc_1386_nl;
  wire[23:0] nl_MultLoop_acc_1386_nl;
  wire[19:0] MultLoop_acc_1999_nl;
  wire[20:0] nl_MultLoop_acc_1999_nl;
  wire[26:0] MultLoop_acc_910_nl;
  wire[28:0] nl_MultLoop_acc_910_nl;
  wire[16:0] MultLoop_914_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_914_MultLoop_acc_3_nl;
  wire[14:0] MultLoop_acc_2007_nl;
  wire[15:0] nl_MultLoop_acc_2007_nl;
  wire[24:0] MultLoop_acc_903_nl;
  wire[25:0] nl_MultLoop_acc_903_nl;
  wire[22:0] MultLoop_acc_2004_nl;
  wire[23:0] nl_MultLoop_acc_2004_nl;
  wire[19:0] MultLoop_acc_2003_nl;
  wire[20:0] nl_MultLoop_acc_2003_nl;
  wire[20:0] MultLoop_acc_902_nl;
  wire[21:0] nl_MultLoop_acc_902_nl;
  wire[17:0] MultLoop_acc_2006_nl;
  wire[18:0] nl_MultLoop_acc_2006_nl;
  wire[22:0] MultLoop_acc_934_nl;
  wire[23:0] nl_MultLoop_acc_934_nl;
  wire[14:0] MultLoop_acc_4016_nl;
  wire[15:0] nl_MultLoop_acc_4016_nl;
  wire[20:0] MultLoop_acc_1392_nl;
  wire[21:0] nl_MultLoop_acc_1392_nl;
  wire[18:0] MultLoop_acc_1931_nl;
  wire[19:0] nl_MultLoop_acc_1931_nl;
  wire[23:0] MultLoop_acc_921_nl;
  wire[25:0] nl_MultLoop_acc_921_nl;
  wire[13:0] MultLoop_acc_4017_nl;
  wire[14:0] nl_MultLoop_acc_4017_nl;
  wire[20:0] MultLoop_acc_917_nl;
  wire[21:0] nl_MultLoop_acc_917_nl;
  wire[16:0] MultLoop_acc_4018_nl;
  wire[17:0] nl_MultLoop_acc_4018_nl;
  wire[18:0] MultLoop_acc_4604_nl;
  wire[19:0] nl_MultLoop_acc_4604_nl;
  wire[17:0] MultLoop_acc_4020_nl;
  wire[18:0] nl_MultLoop_acc_4020_nl;
  wire[22:0] MultLoop_acc_1937_nl;
  wire[23:0] nl_MultLoop_acc_1937_nl;
  wire[19:0] MultLoop_acc_1936_nl;
  wire[20:0] nl_MultLoop_acc_1936_nl;
  wire[19:0] MultLoop_acc_908_nl;
  wire[20:0] nl_MultLoop_acc_908_nl;
  wire[18:0] MultLoop_acc_1939_nl;
  wire[19:0] nl_MultLoop_acc_1939_nl;
  wire[22:0] MultLoop_acc_937_nl;
  wire[24:0] nl_MultLoop_acc_937_nl;
  wire[14:0] MultLoop_acc_4022_nl;
  wire[15:0] nl_MultLoop_acc_4022_nl;
  wire[18:0] MultLoop_acc_4605_nl;
  wire[19:0] nl_MultLoop_acc_4605_nl;
  wire[14:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl;
  wire[18:0] MultLoop_acc_1384_nl;
  wire[19:0] nl_MultLoop_acc_1384_nl;
  wire[13:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl;
  wire[18:0] MultLoop_acc_1400_nl;
  wire[19:0] nl_MultLoop_acc_1400_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[13:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl;
  wire[17:0] MultLoop_acc_945_nl;
  wire[18:0] nl_MultLoop_acc_945_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_8_nl;
  wire[17:0] MultLoop_acc_918_nl;
  wire[18:0] nl_MultLoop_acc_918_nl;
  wire[19:0] MultLoop_acc_1398_nl;
  wire[20:0] nl_MultLoop_acc_1398_nl;
  wire[17:0] MultLoop_acc_1945_nl;
  wire[18:0] nl_MultLoop_acc_1945_nl;
  wire[21:0] MultLoop_acc_1399_nl;
  wire[22:0] nl_MultLoop_acc_1399_nl;
  wire[20:0] MultLoop_acc_1947_nl;
  wire[21:0] nl_MultLoop_acc_1947_nl;
  wire[21:0] MultLoop_acc_1387_nl;
  wire[22:0] nl_MultLoop_acc_1387_nl;
  wire[18:0] MultLoop_acc_1944_nl;
  wire[19:0] nl_MultLoop_acc_1944_nl;
  wire[17:0] MultLoop_acc_4024_nl;
  wire[18:0] nl_MultLoop_acc_4024_nl;
  wire[23:0] MultLoop_acc_1951_nl;
  wire[25:0] nl_MultLoop_acc_1951_nl;
  wire[24:0] MultLoop_acc_942_nl;
  wire[26:0] nl_MultLoop_acc_942_nl;
  wire[19:0] MultLoop_acc_1952_nl;
  wire[20:0] nl_MultLoop_acc_1952_nl;
  wire[22:0] MultLoop_acc_1397_nl;
  wire[23:0] nl_MultLoop_acc_1397_nl;
  wire[20:0] MultLoop_acc_1955_nl;
  wire[21:0] nl_MultLoop_acc_1955_nl;
  wire[17:0] MultLoop_acc_1954_nl;
  wire[18:0] nl_MultLoop_acc_1954_nl;
  wire[24:0] MultLoop_acc_936_nl;
  wire[26:0] nl_MultLoop_acc_936_nl;
  wire[25:0] MultLoop_acc_931_nl;
  wire[26:0] nl_MultLoop_acc_931_nl;
  wire[17:0] MultLoop_acc_4028_nl;
  wire[18:0] nl_MultLoop_acc_4028_nl;
  wire[19:0] MultLoop_acc_1961_nl;
  wire[20:0] nl_MultLoop_acc_1961_nl;
  wire[18:0] MultLoop_acc_4606_nl;
  wire[19:0] nl_MultLoop_acc_4606_nl;
  wire[22:0] MultLoop_acc_928_nl;
  wire[23:0] nl_MultLoop_acc_928_nl;
  wire[19:0] MultLoop_acc_1965_nl;
  wire[20:0] nl_MultLoop_acc_1965_nl;
  wire[17:0] MultLoop_acc_1964_nl;
  wire[18:0] nl_MultLoop_acc_1964_nl;
  wire[11:0] MultLoop_acc_4029_nl;
  wire[12:0] nl_MultLoop_acc_4029_nl;
  wire[19:0] MultLoop_acc_1391_nl;
  wire[20:0] nl_MultLoop_acc_1391_nl;
  wire[17:0] MultLoop_acc_1977_nl;
  wire[18:0] nl_MultLoop_acc_1977_nl;
  wire[21:0] MultLoop_acc_1390_nl;
  wire[22:0] nl_MultLoop_acc_1390_nl;
  wire[20:0] MultLoop_acc_1979_nl;
  wire[21:0] nl_MultLoop_acc_1979_nl;
  wire[17:0] MultLoop_acc_4031_nl;
  wire[18:0] nl_MultLoop_acc_4031_nl;
  wire[22:0] MultLoop_acc_1969_nl;
  wire[23:0] nl_MultLoop_acc_1969_nl;
  wire[19:0] MultLoop_acc_1968_nl;
  wire[20:0] nl_MultLoop_acc_1968_nl;
  wire[17:0] MultLoop_acc_1967_nl;
  wire[18:0] nl_MultLoop_acc_1967_nl;
  wire[19:0] MultLoop_acc_923_nl;
  wire[20:0] nl_MultLoop_acc_923_nl;
  wire[18:0] MultLoop_acc_1971_nl;
  wire[19:0] nl_MultLoop_acc_1971_nl;
  wire[17:0] MultLoop_acc_4034_nl;
  wire[18:0] nl_MultLoop_acc_4034_nl;
  wire[23:0] MultLoop_acc_1974_nl;
  wire[24:0] nl_MultLoop_acc_1974_nl;
  wire[20:0] MultLoop_acc_1973_nl;
  wire[21:0] nl_MultLoop_acc_1973_nl;
  wire[25:0] MultLoop_acc_922_nl;
  wire[27:0] nl_MultLoop_acc_922_nl;
  wire[20:0] MultLoop_acc_1388_nl;
  wire[21:0] nl_MultLoop_acc_1388_nl;
  wire[17:0] MultLoop_acc_1980_nl;
  wire[18:0] nl_MultLoop_acc_1980_nl;
  wire[22:0] MultLoop_acc_911_nl;
  wire[23:0] nl_MultLoop_acc_911_nl;
  wire[18:0] MultLoop_acc_1982_nl;
  wire[19:0] nl_MultLoop_acc_1982_nl;
  wire[15:0] MultLoop_acc_3470_nl;
  wire[17:0] nl_MultLoop_acc_3470_nl;
  wire[12:0] MultLoop_acc_3456_nl;
  wire[13:0] nl_MultLoop_acc_3456_nl;
  wire[20:0] MultLoop_acc_1142_nl;
  wire[21:0] nl_MultLoop_acc_1142_nl;
  wire[17:0] MultLoop_acc_3386_nl;
  wire[18:0] nl_MultLoop_acc_3386_nl;
  wire[14:0] MultLoop_acc_4442_nl;
  wire[15:0] nl_MultLoop_acc_4442_nl;
  wire[24:0] MultLoop_acc_1158_nl;
  wire[25:0] nl_MultLoop_acc_1158_nl;
  wire[19:0] MultLoop_acc_3444_nl;
  wire[21:0] nl_MultLoop_acc_3444_nl;
  wire[10:0] MultLoop_acc_4443_nl;
  wire[11:0] nl_MultLoop_acc_4443_nl;
  wire[24:0] MultLoop_acc_1155_nl;
  wire[25:0] nl_MultLoop_acc_1155_nl;
  wire[19:0] MultLoop_acc_3446_nl;
  wire[20:0] nl_MultLoop_acc_3446_nl;
  wire[22:0] MultLoop_acc_197_nl;
  wire[23:0] nl_MultLoop_acc_197_nl;
  wire[19:0] MultLoop_acc_3439_nl;
  wire[20:0] nl_MultLoop_acc_3439_nl;
  wire[18:0] MultLoop_acc_4441_nl;
  wire[19:0] nl_MultLoop_acc_4441_nl;
  wire[23:0] MultLoop_acc_1148_nl;
  wire[24:0] nl_MultLoop_acc_1148_nl;
  wire[21:0] MultLoop_acc_3449_nl;
  wire[22:0] nl_MultLoop_acc_3449_nl;
  wire[17:0] MultLoop_acc_3448_nl;
  wire[18:0] nl_MultLoop_acc_3448_nl;
  wire[26:0] MultLoop_acc_212_nl;
  wire[28:0] nl_MultLoop_acc_212_nl;
  wire[10:0] MultLoop_acc_4445_nl;
  wire[11:0] nl_MultLoop_acc_4445_nl;
  wire[26:0] MultLoop_acc_204_nl;
  wire[28:0] nl_MultLoop_acc_204_nl;
  wire[24:0] MultLoop_acc_200_nl;
  wire[25:0] nl_MultLoop_acc_200_nl;
  wire[17:0] MultLoop_acc_4684_nl;
  wire[18:0] nl_MultLoop_acc_4684_nl;
  wire[20:0] MultLoop_acc_1146_nl;
  wire[21:0] nl_MultLoop_acc_1146_nl;
  wire[13:0] MultLoop_193_MultLoop_acc_3_nl;
  wire[14:0] nl_MultLoop_193_MultLoop_acc_3_nl;
  wire[21:0] MultLoop_acc_193_nl;
  wire[22:0] nl_MultLoop_acc_193_nl;
  wire[18:0] MultLoop_acc_3389_nl;
  wire[19:0] nl_MultLoop_acc_3389_nl;
  wire[12:0] MultLoop_acc_4448_nl;
  wire[13:0] nl_MultLoop_acc_4448_nl;
  wire[17:0] MultLoop_acc_4451_nl;
  wire[18:0] nl_MultLoop_acc_4451_nl;
  wire[21:0] MultLoop_acc_3393_nl;
  wire[22:0] nl_MultLoop_acc_3393_nl;
  wire[21:0] MultLoop_acc_232_nl;
  wire[22:0] nl_MultLoop_acc_232_nl;
  wire[20:0] MultLoop_acc_3394_nl;
  wire[21:0] nl_MultLoop_acc_3394_nl;
  wire[18:0] MultLoop_acc_4648_nl;
  wire[19:0] nl_MultLoop_acc_4648_nl;
  wire[23:0] MultLoop_acc_230_nl;
  wire[25:0] nl_MultLoop_acc_230_nl;
  wire[13:0] MultLoop_acc_4452_nl;
  wire[14:0] nl_MultLoop_acc_4452_nl;
  wire[21:0] MultLoop_acc_229_nl;
  wire[22:0] nl_MultLoop_acc_229_nl;
  wire[19:0] MultLoop_acc_3399_nl;
  wire[20:0] nl_MultLoop_acc_3399_nl;
  wire[17:0] MultLoop_acc_226_nl;
  wire[18:0] nl_MultLoop_acc_226_nl;
  wire[21:0] MultLoop_acc_1151_nl;
  wire[22:0] nl_MultLoop_acc_1151_nl;
  wire[17:0] MultLoop_acc_3401_nl;
  wire[18:0] nl_MultLoop_acc_3401_nl;
  wire[20:0] MultLoop_acc_217_nl;
  wire[21:0] nl_MultLoop_acc_217_nl;
  wire[18:0] MultLoop_acc_3403_nl;
  wire[19:0] nl_MultLoop_acc_3403_nl;
  wire[11:0] MultLoop_acc_4455_nl;
  wire[12:0] nl_MultLoop_acc_4455_nl;
  wire[21:0] MultLoop_acc_1150_nl;
  wire[22:0] nl_MultLoop_acc_1150_nl;
  wire[18:0] MultLoop_acc_3404_nl;
  wire[19:0] nl_MultLoop_acc_3404_nl;
  wire[20:0] MultLoop_acc_216_nl;
  wire[21:0] nl_MultLoop_acc_216_nl;
  wire[18:0] MultLoop_acc_3406_nl;
  wire[19:0] nl_MultLoop_acc_3406_nl;
  wire[13:0] MultLoop_acc_4456_nl;
  wire[14:0] nl_MultLoop_acc_4456_nl;
  wire[17:0] MultLoop_acc_4458_nl;
  wire[18:0] nl_MultLoop_acc_4458_nl;
  wire[22:0] MultLoop_acc_3408_nl;
  wire[23:0] nl_MultLoop_acc_3408_nl;
  wire[23:0] MultLoop_acc_208_nl;
  wire[24:0] nl_MultLoop_acc_208_nl;
  wire[13:0] MultLoop_acc_4459_nl;
  wire[14:0] nl_MultLoop_acc_4459_nl;
  wire[24:0] MultLoop_acc_201_nl;
  wire[26:0] nl_MultLoop_acc_201_nl;
  wire[12:0] MultLoop_acc_4460_nl;
  wire[13:0] nl_MultLoop_acc_4460_nl;
  wire[18:0] MultLoop_acc_4649_nl;
  wire[19:0] nl_MultLoop_acc_4649_nl;
  wire[21:0] MultLoop_acc_1143_nl;
  wire[22:0] nl_MultLoop_acc_1143_nl;
  wire[18:0] MultLoop_acc_3413_nl;
  wire[19:0] nl_MultLoop_acc_3413_nl;
  wire[25:0] MultLoop_acc_238_nl;
  wire[27:0] nl_MultLoop_acc_238_nl;
  wire[17:0] MultLoop_acc_4463_nl;
  wire[18:0] nl_MultLoop_acc_4463_nl;
  wire[22:0] MultLoop_acc_3419_nl;
  wire[24:0] nl_MultLoop_acc_3419_nl;
  wire[23:0] MultLoop_acc_1157_nl;
  wire[24:0] nl_MultLoop_acc_1157_nl;
  wire[20:0] MultLoop_acc_3421_nl;
  wire[22:0] nl_MultLoop_acc_3421_nl;
  wire[18:0] MultLoop_acc_1153_nl;
  wire[19:0] nl_MultLoop_acc_1153_nl;
  wire[20:0] MultLoop_acc_220_nl;
  wire[21:0] nl_MultLoop_acc_220_nl;
  wire[18:0] MultLoop_acc_3423_nl;
  wire[19:0] nl_MultLoop_acc_3423_nl;
  wire[11:0] MultLoop_acc_4464_nl;
  wire[12:0] nl_MultLoop_acc_4464_nl;
  wire[21:0] MultLoop_acc_1147_nl;
  wire[22:0] nl_MultLoop_acc_1147_nl;
  wire[17:0] MultLoop_acc_3432_nl;
  wire[18:0] nl_MultLoop_acc_3432_nl;
  wire[13:0] MultLoop_acc_4469_nl;
  wire[14:0] nl_MultLoop_acc_4469_nl;
  wire[17:0] MultLoop_acc_4471_nl;
  wire[18:0] nl_MultLoop_acc_4471_nl;
  wire[22:0] MultLoop_acc_3436_nl;
  wire[23:0] nl_MultLoop_acc_3436_nl;
  wire[19:0] MultLoop_acc_3435_nl;
  wire[20:0] nl_MultLoop_acc_3435_nl;
  wire[17:0] MultLoop_acc_3434_nl;
  wire[18:0] nl_MultLoop_acc_3434_nl;
  wire[24:0] MultLoop_acc_221_nl;
  wire[25:0] nl_MultLoop_acc_221_nl;
  wire[21:0] MultLoop_acc_218_nl;
  wire[22:0] nl_MultLoop_acc_218_nl;
  wire[19:0] MultLoop_acc_3427_nl;
  wire[20:0] nl_MultLoop_acc_3427_nl;
  wire[17:0] MultLoop_acc_3426_nl;
  wire[18:0] nl_MultLoop_acc_3426_nl;
  wire[11:0] MultLoop_acc_4466_nl;
  wire[12:0] nl_MultLoop_acc_4466_nl;
  wire[18:0] MultLoop_acc_1149_nl;
  wire[19:0] nl_MultLoop_acc_1149_nl;
  wire[17:0] MultLoop_acc_4468_nl;
  wire[18:0] nl_MultLoop_acc_4468_nl;
  wire[23:0] MultLoop_acc_3430_nl;
  wire[24:0] nl_MultLoop_acc_3430_nl;
  wire[20:0] MultLoop_acc_3429_nl;
  wire[21:0] nl_MultLoop_acc_3429_nl;
  wire[10:0] MultLoop_acc_4467_nl;
  wire[11:0] nl_MultLoop_acc_4467_nl;
  wire[19:0] MultLoop_acc_4650_nl;
  wire[20:0] nl_MultLoop_acc_4650_nl;
  wire[22:0] MultLoop_acc_203_nl;
  wire[23:0] nl_MultLoop_acc_203_nl;
  wire[21:0] MultLoop_acc_3438_nl;
  wire[22:0] nl_MultLoop_acc_3438_nl;
  wire[19:0] MultLoop_acc_1368_nl;
  wire[20:0] nl_MultLoop_acc_1368_nl;
  wire[17:0] MultLoop_acc_2063_nl;
  wire[18:0] nl_MultLoop_acc_2063_nl;
  wire[23:0] MultLoop_acc_1366_nl;
  wire[24:0] nl_MultLoop_acc_1366_nl;
  wire[20:0] MultLoop_acc_2066_nl;
  wire[22:0] nl_MultLoop_acc_2066_nl;
  wire[11:0] MultLoop_acc_4040_nl;
  wire[12:0] nl_MultLoop_acc_4040_nl;
  wire[19:0] MultLoop_acc_1369_nl;
  wire[20:0] nl_MultLoop_acc_1369_nl;
  wire[17:0] MultLoop_acc_2056_nl;
  wire[18:0] nl_MultLoop_acc_2056_nl;
  wire[23:0] MultLoop_acc_1370_nl;
  wire[24:0] nl_MultLoop_acc_1370_nl;
  wire[21:0] MultLoop_acc_2058_nl;
  wire[22:0] nl_MultLoop_acc_2058_nl;
  wire[17:0] MultLoop_acc_4038_nl;
  wire[18:0] nl_MultLoop_acc_4038_nl;
  wire[23:0] MultLoop_acc_2060_nl;
  wire[24:0] nl_MultLoop_acc_2060_nl;
  wire[22:0] MultLoop_acc_1367_nl;
  wire[23:0] nl_MultLoop_acc_1367_nl;
  wire[17:0] MultLoop_acc_2062_nl;
  wire[18:0] nl_MultLoop_acc_2062_nl;
  wire[20:0] MultLoop_acc_1363_nl;
  wire[21:0] nl_MultLoop_acc_1363_nl;
  wire[17:0] MultLoop_acc_2067_nl;
  wire[18:0] nl_MultLoop_acc_2067_nl;
  wire[15:0] MultLoop_866_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_866_MultLoop_acc_3_nl;
  wire[14:0] MultLoop_acc_2068_nl;
  wire[15:0] nl_MultLoop_acc_2068_nl;
  wire[18:0] MultLoop_acc_855_nl;
  wire[19:0] nl_MultLoop_acc_855_nl;
  wire[18:0] MultLoop_acc_4607_nl;
  wire[19:0] nl_MultLoop_acc_4607_nl;
  wire[18:0] MultLoop_acc_4044_nl;
  wire[19:0] nl_MultLoop_acc_4044_nl;
  wire[24:0] MultLoop_acc_2075_nl;
  wire[25:0] nl_MultLoop_acc_2075_nl;
  wire[20:0] MultLoop_acc_2074_nl;
  wire[21:0] nl_MultLoop_acc_2074_nl;
  wire[17:0] MultLoop_acc_4042_nl;
  wire[18:0] nl_MultLoop_acc_4042_nl;
  wire[20:0] MultLoop_acc_2070_nl;
  wire[21:0] nl_MultLoop_acc_2070_nl;
  wire[23:0] MultLoop_acc_1362_nl;
  wire[24:0] nl_MultLoop_acc_1362_nl;
  wire[18:0] MultLoop_acc_4045_nl;
  wire[19:0] nl_MultLoop_acc_4045_nl;
  wire[24:0] MultLoop_acc_2077_nl;
  wire[25:0] nl_MultLoop_acc_2077_nl;
  wire[19:0] MultLoop_acc_2076_nl;
  wire[20:0] nl_MultLoop_acc_2076_nl;
  wire[24:0] MultLoop_acc_874_nl;
  wire[25:0] nl_MultLoop_acc_874_nl;
  wire[21:0] MultLoop_acc_2078_nl;
  wire[22:0] nl_MultLoop_acc_2078_nl;
  wire[22:0] MultLoop_acc_1365_nl;
  wire[23:0] nl_MultLoop_acc_1365_nl;
  wire[19:0] MultLoop_acc_2080_nl;
  wire[20:0] nl_MultLoop_acc_2080_nl;
  wire[18:0] MultLoop_acc_4608_nl;
  wire[19:0] nl_MultLoop_acc_4608_nl;
  wire[21:0] MultLoop_acc_892_nl;
  wire[22:0] nl_MultLoop_acc_892_nl;
  wire[15:0] MultLoop_acc_4046_nl;
  wire[16:0] nl_MultLoop_acc_4046_nl;
  wire[19:0] MultLoop_acc_4667_nl;
  wire[20:0] nl_MultLoop_acc_4667_nl;
  wire[17:0] MultLoop_acc_4048_nl;
  wire[18:0] nl_MultLoop_acc_4048_nl;
  wire[21:0] MultLoop_acc_2012_nl;
  wire[22:0] nl_MultLoop_acc_2012_nl;
  wire[19:0] MultLoop_acc_877_nl;
  wire[20:0] nl_MultLoop_acc_877_nl;
  wire[18:0] MultLoop_acc_2014_nl;
  wire[19:0] nl_MultLoop_acc_2014_nl;
  wire[19:0] MultLoop_acc_4609_nl;
  wire[20:0] nl_MultLoop_acc_4609_nl;
  wire[12:0] MultLoop_acc_2082_nl;
  wire[13:0] nl_MultLoop_acc_2082_nl;
  wire[22:0] MultLoop_acc_888_nl;
  wire[23:0] nl_MultLoop_acc_888_nl;
  wire[14:0] MultLoop_acc_4050_nl;
  wire[15:0] nl_MultLoop_acc_4050_nl;
  wire[19:0] MultLoop_acc_1374_nl;
  wire[20:0] nl_MultLoop_acc_1374_nl;
  wire[17:0] MultLoop_acc_2016_nl;
  wire[18:0] nl_MultLoop_acc_2016_nl;
  wire[18:0] MultLoop_acc_4610_nl;
  wire[19:0] nl_MultLoop_acc_4610_nl;
  wire[21:0] MultLoop_acc_1373_nl;
  wire[22:0] nl_MultLoop_acc_1373_nl;
  wire[20:0] MultLoop_acc_2019_nl;
  wire[21:0] nl_MultLoop_acc_2019_nl;
  wire[17:0] MultLoop_acc_2018_nl;
  wire[18:0] nl_MultLoop_acc_2018_nl;
  wire[22:0] MultLoop_acc_1371_nl;
  wire[23:0] nl_MultLoop_acc_1371_nl;
  wire[17:0] MultLoop_acc_2021_nl;
  wire[18:0] nl_MultLoop_acc_2021_nl;
  wire[12:0] MultLoop_acc_4051_nl;
  wire[13:0] nl_MultLoop_acc_4051_nl;
  wire[17:0] MultLoop_acc_4053_nl;
  wire[18:0] nl_MultLoop_acc_4053_nl;
  wire[23:0] MultLoop_acc_2024_nl;
  wire[24:0] nl_MultLoop_acc_2024_nl;
  wire[19:0] MultLoop_acc_2023_nl;
  wire[20:0] nl_MultLoop_acc_2023_nl;
  wire[18:0] MultLoop_acc_4611_nl;
  wire[19:0] nl_MultLoop_acc_4611_nl;
  wire[17:0] MultLoop_acc_4055_nl;
  wire[18:0] nl_MultLoop_acc_4055_nl;
  wire[22:0] MultLoop_acc_2028_nl;
  wire[23:0] nl_MultLoop_acc_2028_nl;
  wire[24:0] MultLoop_acc_897_nl;
  wire[26:0] nl_MultLoop_acc_897_nl;
  wire[20:0] MultLoop_acc_1383_nl;
  wire[21:0] nl_MultLoop_acc_1383_nl;
  wire[17:0] MultLoop_acc_2032_nl;
  wire[18:0] nl_MultLoop_acc_2032_nl;
  wire[18:0] MultLoop_acc_4057_nl;
  wire[19:0] nl_MultLoop_acc_4057_nl;
  wire[18:0] MultLoop_acc_4612_nl;
  wire[19:0] nl_MultLoop_acc_4612_nl;
  wire[23:0] MultLoop_acc_1382_nl;
  wire[24:0] nl_MultLoop_acc_1382_nl;
  wire[21:0] MultLoop_acc_2037_nl;
  wire[22:0] nl_MultLoop_acc_2037_nl;
  wire[19:0] MultLoop_acc_2036_nl;
  wire[20:0] nl_MultLoop_acc_2036_nl;
  wire[20:0] MultLoop_acc_1380_nl;
  wire[21:0] nl_MultLoop_acc_1380_nl;
  wire[17:0] MultLoop_acc_2039_nl;
  wire[18:0] nl_MultLoop_acc_2039_nl;
  wire[23:0] MultLoop_acc_1372_nl;
  wire[24:0] nl_MultLoop_acc_1372_nl;
  wire[22:0] MultLoop_acc_2047_nl;
  wire[23:0] nl_MultLoop_acc_2047_nl;
  wire[19:0] MultLoop_acc_2046_nl;
  wire[21:0] nl_MultLoop_acc_2046_nl;
  wire[17:0] MultLoop_acc_4062_nl;
  wire[18:0] nl_MultLoop_acc_4062_nl;
  wire[22:0] MultLoop_acc_2050_nl;
  wire[24:0] nl_MultLoop_acc_2050_nl;
  wire[18:0] MultLoop_acc_4613_nl;
  wire[19:0] nl_MultLoop_acc_4613_nl;
  wire[22:0] MultLoop_acc_1376_nl;
  wire[23:0] nl_MultLoop_acc_1376_nl;
  wire[17:0] MultLoop_acc_2042_nl;
  wire[18:0] nl_MultLoop_acc_2042_nl;
  wire[12:0] MultLoop_acc_4059_nl;
  wire[13:0] nl_MultLoop_acc_4059_nl;
  wire[20:0] MultLoop_acc_878_nl;
  wire[21:0] nl_MultLoop_acc_878_nl;
  wire[18:0] MultLoop_acc_2044_nl;
  wire[19:0] nl_MultLoop_acc_2044_nl;
  wire[25:0] MultLoop_acc_871_nl;
  wire[26:0] nl_MultLoop_acc_871_nl;
  wire[22:0] MultLoop_acc_2053_nl;
  wire[23:0] nl_MultLoop_acc_2053_nl;
  wire[20:0] MultLoop_acc_2052_nl;
  wire[21:0] nl_MultLoop_acc_2052_nl;
  wire[11:0] MultLoop_acc_4063_nl;
  wire[12:0] nl_MultLoop_acc_4063_nl;
  wire[25:0] MultLoop_acc_870_nl;
  wire[26:0] nl_MultLoop_acc_870_nl;
  wire[24:0] MultLoop_acc_2055_nl;
  wire[26:0] nl_MultLoop_acc_2055_nl;
  wire[21:0] MultLoop_acc_1167_nl;
  wire[22:0] nl_MultLoop_acc_1167_nl;
  wire[17:0] MultLoop_acc_3328_nl;
  wire[18:0] nl_MultLoop_acc_3328_nl;
  wire[13:0] MultLoop_acc_4415_nl;
  wire[14:0] nl_MultLoop_acc_4415_nl;
  wire[20:0] MultLoop_acc_1166_nl;
  wire[21:0] nl_MultLoop_acc_1166_nl;
  wire[18:0] MultLoop_acc_3329_nl;
  wire[19:0] nl_MultLoop_acc_3329_nl;
  wire[25:0] MultLoop_acc_256_nl;
  wire[27:0] nl_MultLoop_acc_256_nl;
  wire[26:0] MultLoop_acc_254_nl;
  wire[28:0] nl_MultLoop_acc_254_nl;
  wire[10:0] MultLoop_acc_4417_nl;
  wire[11:0] nl_MultLoop_acc_4417_nl;
  wire[16:0] MultLoop_248_MultLoop_acc_3_nl;
  wire[18:0] nl_MultLoop_248_MultLoop_acc_3_nl;
  wire[15:0] MultLoop_244_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_244_MultLoop_acc_3_nl;
  wire[14:0] MultLoop_acc_3341_nl;
  wire[16:0] nl_MultLoop_acc_3341_nl;
  wire[17:0] MultLoop_acc_243_nl;
  wire[18:0] nl_MultLoop_acc_243_nl;
  wire[12:0] MultLoop_241_MultLoop_acc_3_nl;
  wire[13:0] nl_MultLoop_241_MultLoop_acc_3_nl;
  wire[17:0] MultLoop_acc_240_nl;
  wire[18:0] nl_MultLoop_acc_240_nl;
  wire[17:0] MultLoop_acc_242_nl;
  wire[18:0] nl_MultLoop_acc_242_nl;
  wire[18:0] MultLoop_acc_4419_nl;
  wire[19:0] nl_MultLoop_acc_4419_nl;
  wire[19:0] MultLoop_acc_4645_nl;
  wire[20:0] nl_MultLoop_acc_4645_nl;
  wire[21:0] MultLoop_acc_1159_nl;
  wire[22:0] nl_MultLoop_acc_1159_nl;
  wire[18:0] MultLoop_acc_3342_nl;
  wire[19:0] nl_MultLoop_acc_3342_nl;
  wire[14:0] MultLoop_acc_3344_nl;
  wire[15:0] nl_MultLoop_acc_3344_nl;
  wire[24:0] MultLoop_acc_247_nl;
  wire[26:0] nl_MultLoop_acc_247_nl;
  wire[12:0] MultLoop_acc_3343_nl;
  wire[13:0] nl_MultLoop_acc_3343_nl;
  wire[13:0] MultLoop_acc_3348_nl;
  wire[14:0] nl_MultLoop_acc_3348_nl;
  wire[20:0] MultLoop_acc_269_nl;
  wire[21:0] nl_MultLoop_acc_269_nl;
  wire[16:0] MultLoop_acc_4420_nl;
  wire[17:0] nl_MultLoop_acc_4420_nl;
  wire[12:0] MultLoop_acc_3346_nl;
  wire[13:0] nl_MultLoop_acc_3346_nl;
  wire[21:0] MultLoop_acc_250_nl;
  wire[22:0] nl_MultLoop_acc_250_nl;
  wire[15:0] MultLoop_acc_4421_nl;
  wire[16:0] nl_MultLoop_acc_4421_nl;
  wire[21:0] MultLoop_acc_282_nl;
  wire[22:0] nl_MultLoop_acc_282_nl;
  wire[20:0] MultLoop_acc_3267_nl;
  wire[21:0] nl_MultLoop_acc_3267_nl;
  wire[20:0] MultLoop_acc_1163_nl;
  wire[21:0] nl_MultLoop_acc_1163_nl;
  wire[19:0] MultLoop_acc_271_nl;
  wire[20:0] nl_MultLoop_acc_271_nl;
  wire[18:0] MultLoop_acc_3271_nl;
  wire[19:0] nl_MultLoop_acc_3271_nl;
  wire[21:0] MultLoop_acc_1174_nl;
  wire[22:0] nl_MultLoop_acc_1174_nl;
  wire[20:0] MultLoop_acc_3274_nl;
  wire[21:0] nl_MultLoop_acc_3274_nl;
  wire[19:0] MultLoop_acc_1173_nl;
  wire[20:0] nl_MultLoop_acc_1173_nl;
  wire[17:0] MultLoop_acc_3275_nl;
  wire[18:0] nl_MultLoop_acc_3275_nl;
  wire[22:0] MultLoop_acc_1172_nl;
  wire[23:0] nl_MultLoop_acc_1172_nl;
  wire[20:0] MultLoop_acc_3277_nl;
  wire[21:0] nl_MultLoop_acc_3277_nl;
  wire[24:0] MultLoop_acc_275_nl;
  wire[25:0] nl_MultLoop_acc_275_nl;
  wire[22:0] MultLoop_acc_3279_nl;
  wire[23:0] nl_MultLoop_acc_3279_nl;
  wire[20:0] MultLoop_acc_4646_nl;
  wire[21:0] nl_MultLoop_acc_4646_nl;
  wire[18:0] MultLoop_acc_4647_nl;
  wire[19:0] nl_MultLoop_acc_4647_nl;
  wire[21:0] MultLoop_acc_270_nl;
  wire[22:0] nl_MultLoop_acc_270_nl;
  wire[20:0] MultLoop_acc_3282_nl;
  wire[21:0] nl_MultLoop_acc_3282_nl;
  wire[22:0] MultLoop_acc_1169_nl;
  wire[23:0] nl_MultLoop_acc_1169_nl;
  wire[20:0] MultLoop_acc_3284_nl;
  wire[21:0] nl_MultLoop_acc_3284_nl;
  wire[17:0] MultLoop_acc_4424_nl;
  wire[18:0] nl_MultLoop_acc_4424_nl;
  wire[21:0] MultLoop_acc_3290_nl;
  wire[22:0] nl_MultLoop_acc_3290_nl;
  wire[19:0] MultLoop_acc_3289_nl;
  wire[21:0] nl_MultLoop_acc_3289_nl;
  wire[18:0] MultLoop_acc_1164_nl;
  wire[19:0] nl_MultLoop_acc_1164_nl;
  wire[23:0] MultLoop_acc_249_nl;
  wire[24:0] nl_MultLoop_acc_249_nl;
  wire[22:0] MultLoop_acc_3286_nl;
  wire[24:0] nl_MultLoop_acc_3286_nl;
  wire[25:0] MultLoop_acc_284_nl;
  wire[27:0] nl_MultLoop_acc_284_nl;
  wire[23:0] MultLoop_acc_281_nl;
  wire[24:0] nl_MultLoop_acc_281_nl;
  wire[21:0] MultLoop_acc_3293_nl;
  wire[22:0] nl_MultLoop_acc_3293_nl;
  wire[17:0] MultLoop_acc_4427_nl;
  wire[18:0] nl_MultLoop_acc_4427_nl;
  wire[24:0] MultLoop_acc_3296_nl;
  wire[25:0] nl_MultLoop_acc_3296_nl;
  wire[19:0] MultLoop_acc_3295_nl;
  wire[20:0] nl_MultLoop_acc_3295_nl;
  wire[24:0] MultLoop_acc_280_nl;
  wire[26:0] nl_MultLoop_acc_280_nl;
  wire[17:0] MultLoop_acc_4430_nl;
  wire[18:0] nl_MultLoop_acc_4430_nl;
  wire[21:0] MultLoop_acc_3301_nl;
  wire[22:0] nl_MultLoop_acc_3301_nl;
  wire[17:0] MultLoop_acc_3300_nl;
  wire[18:0] nl_MultLoop_acc_3300_nl;
  wire[10:0] MultLoop_acc_4429_nl;
  wire[11:0] nl_MultLoop_acc_4429_nl;
  wire[17:0] MultLoop_acc_4432_nl;
  wire[18:0] nl_MultLoop_acc_4432_nl;
  wire[23:0] MultLoop_acc_3304_nl;
  wire[24:0] nl_MultLoop_acc_3304_nl;
  wire[19:0] MultLoop_acc_3303_nl;
  wire[20:0] nl_MultLoop_acc_3303_nl;
  wire[10:0] MultLoop_acc_4431_nl;
  wire[11:0] nl_MultLoop_acc_4431_nl;
  wire[25:0] MultLoop_acc_268_nl;
  wire[26:0] nl_MultLoop_acc_268_nl;
  wire[17:0] MultLoop_acc_4434_nl;
  wire[18:0] nl_MultLoop_acc_4434_nl;
  wire[23:0] MultLoop_acc_3308_nl;
  wire[25:0] nl_MultLoop_acc_3308_nl;
  wire[10:0] MultLoop_acc_4433_nl;
  wire[11:0] nl_MultLoop_acc_4433_nl;
  wire[20:0] MultLoop_acc_1165_nl;
  wire[21:0] nl_MultLoop_acc_1165_nl;
  wire[18:0] MultLoop_acc_3309_nl;
  wire[19:0] nl_MultLoop_acc_3309_nl;
  wire[22:0] MultLoop_acc_259_nl;
  wire[23:0] nl_MultLoop_acc_259_nl;
  wire[20:0] MultLoop_acc_3312_nl;
  wire[21:0] nl_MultLoop_acc_3312_nl;
  wire[17:0] MultLoop_acc_3311_nl;
  wire[18:0] nl_MultLoop_acc_3311_nl;
  wire[11:0] MultLoop_acc_4435_nl;
  wire[12:0] nl_MultLoop_acc_4435_nl;
  wire[17:0] MultLoop_acc_4437_nl;
  wire[18:0] nl_MultLoop_acc_4437_nl;
  wire[23:0] MultLoop_acc_3315_nl;
  wire[24:0] nl_MultLoop_acc_3315_nl;
  wire[19:0] MultLoop_acc_3314_nl;
  wire[20:0] nl_MultLoop_acc_3314_nl;
  wire[11:0] MultLoop_acc_4436_nl;
  wire[12:0] nl_MultLoop_acc_4436_nl;
  wire[25:0] MultLoop_acc_255_nl;
  wire[26:0] nl_MultLoop_acc_255_nl;
  wire[22:0] MultLoop_acc_3316_nl;
  wire[23:0] nl_MultLoop_acc_3316_nl;
  wire[22:0] MultLoop_acc_1170_nl;
  wire[23:0] nl_MultLoop_acc_1170_nl;
  wire[18:0] MultLoop_acc_3323_nl;
  wire[19:0] nl_MultLoop_acc_3323_nl;
  wire[23:0] MultLoop_acc_1168_nl;
  wire[24:0] nl_MultLoop_acc_1168_nl;
  wire[19:0] MultLoop_acc_3326_nl;
  wire[21:0] nl_MultLoop_acc_3326_nl;
  wire[10:0] MultLoop_acc_4440_nl;
  wire[11:0] nl_MultLoop_acc_4440_nl;
  wire[22:0] MultLoop_acc_252_nl;
  wire[23:0] nl_MultLoop_acc_252_nl;
  wire[20:0] MultLoop_acc_3318_nl;
  wire[21:0] nl_MultLoop_acc_3318_nl;
  wire[13:0] MultLoop_acc_4438_nl;
  wire[14:0] nl_MultLoop_acc_4438_nl;
  wire[23:0] MultLoop_acc_1162_nl;
  wire[24:0] nl_MultLoop_acc_1162_nl;
  wire[17:0] MultLoop_acc_3320_nl;
  wire[18:0] nl_MultLoop_acc_3320_nl;
  wire[19:0] MultLoop_acc_1161_nl;
  wire[20:0] nl_MultLoop_acc_1161_nl;
  wire[17:0] MultLoop_acc_3321_nl;
  wire[18:0] nl_MultLoop_acc_3321_nl;
  wire[21:0] MultLoop_acc_4694_nl;
  wire[22:0] nl_MultLoop_acc_4694_nl;
  wire[22:0] MultLoop_acc_4668_nl;
  wire[23:0] nl_MultLoop_acc_4668_nl;
  wire[23:0] MultLoop_acc_1356_nl;
  wire[24:0] nl_MultLoop_acc_1356_nl;
  wire[20:0] MultLoop_acc_2178_nl;
  wire[21:0] nl_MultLoop_acc_2178_nl;
  wire[17:0] MultLoop_acc_2177_nl;
  wire[18:0] nl_MultLoop_acc_2177_nl;
  wire[11:0] MultLoop_acc_4066_nl;
  wire[12:0] nl_MultLoop_acc_4066_nl;
  wire[24:0] MultLoop_acc_1352_nl;
  wire[25:0] nl_MultLoop_acc_1352_nl;
  wire[21:0] MultLoop_acc_2182_nl;
  wire[23:0] nl_MultLoop_acc_2182_nl;
  wire[18:0] MultLoop_acc_4064_nl;
  wire[19:0] nl_MultLoop_acc_4064_nl;
  wire[22:0] MultLoop_acc_2173_nl;
  wire[23:0] nl_MultLoop_acc_2173_nl;
  wire[14:0] MultLoop_acc_806_nl;
  wire[15:0] nl_MultLoop_acc_806_nl;
  wire[25:0] MultLoop_acc_828_nl;
  wire[27:0] nl_MultLoop_acc_828_nl;
  wire[23:0] MultLoop_acc_821_nl;
  wire[25:0] nl_MultLoop_acc_821_nl;
  wire[13:0] MultLoop_acc_4069_nl;
  wire[14:0] nl_MultLoop_acc_4069_nl;
  wire[23:0] MultLoop_acc_815_nl;
  wire[25:0] nl_MultLoop_acc_815_nl;
  wire[13:0] MultLoop_acc_4070_nl;
  wire[14:0] nl_MultLoop_acc_4070_nl;
  wire[13:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl;
  wire[19:0] MultLoop_acc_852_nl;
  wire[20:0] nl_MultLoop_acc_852_nl;
  wire[18:0] MultLoop_acc_2129_nl;
  wire[19:0] nl_MultLoop_acc_2129_nl;
  wire[14:0] MultLoop_acc_4071_nl;
  wire[15:0] nl_MultLoop_acc_4071_nl;
  wire[21:0] MultLoop_acc_810_nl;
  wire[22:0] nl_MultLoop_acc_810_nl;
  wire[20:0] MultLoop_acc_2127_nl;
  wire[21:0] nl_MultLoop_acc_2127_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_7_nl;
  wire[18:0] MultLoop_acc_1361_nl;
  wire[19:0] nl_MultLoop_acc_1361_nl;
  wire[23:0] MultLoop_acc_848_nl;
  wire[25:0] nl_MultLoop_acc_848_nl;
  wire[22:0] MultLoop_acc_838_nl;
  wire[23:0] nl_MultLoop_acc_838_nl;
  wire[14:0] MultLoop_acc_4073_nl;
  wire[15:0] nl_MultLoop_acc_4073_nl;
  wire[19:0] MultLoop_acc_1355_nl;
  wire[20:0] nl_MultLoop_acc_1355_nl;
  wire[18:0] MultLoop_acc_1353_nl;
  wire[19:0] nl_MultLoop_acc_1353_nl;
  wire[20:0] MultLoop_acc_851_nl;
  wire[21:0] nl_MultLoop_acc_851_nl;
  wire[23:0] MultLoop_acc_824_nl;
  wire[25:0] nl_MultLoop_acc_824_nl;
  wire[13:0] MultLoop_acc_4074_nl;
  wire[14:0] nl_MultLoop_acc_4074_nl;
  wire[20:0] MultLoop_acc_822_nl;
  wire[21:0] nl_MultLoop_acc_822_nl;
  wire[18:0] MultLoop_acc_2137_nl;
  wire[19:0] nl_MultLoop_acc_2137_nl;
  wire[20:0] MultLoop_acc_847_nl;
  wire[21:0] nl_MultLoop_acc_847_nl;
  wire[18:0] MultLoop_acc_2139_nl;
  wire[19:0] nl_MultLoop_acc_2139_nl;
  wire[17:0] MultLoop_acc_4078_nl;
  wire[18:0] nl_MultLoop_acc_4078_nl;
  wire[20:0] MultLoop_acc_2141_nl;
  wire[21:0] nl_MultLoop_acc_2141_nl;
  wire[17:0] MultLoop_acc_4080_nl;
  wire[18:0] nl_MultLoop_acc_4080_nl;
  wire[21:0] MultLoop_acc_2144_nl;
  wire[23:0] nl_MultLoop_acc_2144_nl;
  wire[18:0] MultLoop_acc_4614_nl;
  wire[19:0] nl_MultLoop_acc_4614_nl;
  wire[18:0] MultLoop_acc_1348_nl;
  wire[19:0] nl_MultLoop_acc_1348_nl;
  wire[21:0] MultLoop_acc_1347_nl;
  wire[22:0] nl_MultLoop_acc_1347_nl;
  wire[19:0] MultLoop_acc_2147_nl;
  wire[21:0] nl_MultLoop_acc_2147_nl;
  wire[21:0] MultLoop_acc_814_nl;
  wire[22:0] nl_MultLoop_acc_814_nl;
  wire[15:0] MultLoop_acc_4081_nl;
  wire[16:0] nl_MultLoop_acc_4081_nl;
  wire[21:0] MultLoop_acc_1345_nl;
  wire[22:0] nl_MultLoop_acc_1345_nl;
  wire[17:0] MultLoop_acc_2149_nl;
  wire[18:0] nl_MultLoop_acc_2149_nl;
  wire[20:0] MultLoop_acc_808_nl;
  wire[21:0] nl_MultLoop_acc_808_nl;
  wire[16:0] MultLoop_acc_4082_nl;
  wire[17:0] nl_MultLoop_acc_4082_nl;
  wire[18:0] MultLoop_acc_4615_nl;
  wire[19:0] nl_MultLoop_acc_4615_nl;
  wire[21:0] MultLoop_acc_849_nl;
  wire[22:0] nl_MultLoop_acc_849_nl;
  wire[20:0] MultLoop_acc_2154_nl;
  wire[22:0] nl_MultLoop_acc_2154_nl;
  wire[23:0] MultLoop_acc_846_nl;
  wire[24:0] nl_MultLoop_acc_846_nl;
  wire[21:0] MultLoop_acc_2156_nl;
  wire[22:0] nl_MultLoop_acc_2156_nl;
  wire[19:0] MultLoop_acc_2155_nl;
  wire[20:0] nl_MultLoop_acc_2155_nl;
  wire[22:0] MultLoop_acc_840_nl;
  wire[23:0] nl_MultLoop_acc_840_nl;
  wire[18:0] MultLoop_acc_2158_nl;
  wire[19:0] nl_MultLoop_acc_2158_nl;
  wire[22:0] MultLoop_acc_1357_nl;
  wire[23:0] nl_MultLoop_acc_1357_nl;
  wire[19:0] MultLoop_acc_2161_nl;
  wire[21:0] nl_MultLoop_acc_2161_nl;
  wire[22:0] MultLoop_acc_823_nl;
  wire[23:0] nl_MultLoop_acc_823_nl;
  wire[19:0] MultLoop_acc_2171_nl;
  wire[20:0] nl_MultLoop_acc_2171_nl;
  wire[17:0] MultLoop_acc_2170_nl;
  wire[18:0] nl_MultLoop_acc_2170_nl;
  wire[25:0] MultLoop_acc_835_nl;
  wire[27:0] nl_MultLoop_acc_835_nl;
  wire[11:0] MultLoop_acc_4086_nl;
  wire[12:0] nl_MultLoop_acc_4086_nl;
  wire[22:0] MultLoop_acc_1354_nl;
  wire[23:0] nl_MultLoop_acc_1354_nl;
  wire[17:0] MultLoop_acc_2165_nl;
  wire[18:0] nl_MultLoop_acc_2165_nl;
  wire[22:0] MultLoop_acc_1351_nl;
  wire[23:0] nl_MultLoop_acc_1351_nl;
  wire[19:0] MultLoop_acc_2168_nl;
  wire[21:0] nl_MultLoop_acc_2168_nl;
  wire[11:0] MultLoop_acc_4088_nl;
  wire[12:0] nl_MultLoop_acc_4088_nl;
  wire[18:0] MultLoop_acc_1349_nl;
  wire[19:0] nl_MultLoop_acc_1349_nl;
  wire[19:0] MultLoop_acc_4616_nl;
  wire[20:0] nl_MultLoop_acc_4616_nl;
  wire[18:0] MultLoop_acc_1346_nl;
  wire[19:0] nl_MultLoop_acc_1346_nl;
  wire[17:0] MultLoop_acc_3259_nl;
  wire[19:0] nl_MultLoop_acc_3259_nl;
  wire[24:0] MultLoop_acc_317_nl;
  wire[25:0] nl_MultLoop_acc_317_nl;
  wire[22:0] MultLoop_acc_3207_nl;
  wire[23:0] nl_MultLoop_acc_3207_nl;
  wire[18:0] MultLoop_acc_4401_nl;
  wire[19:0] nl_MultLoop_acc_4401_nl;
  wire[23:0] MultLoop_acc_3210_nl;
  wire[24:0] nl_MultLoop_acc_3210_nl;
  wire[21:0] MultLoop_acc_3209_nl;
  wire[22:0] nl_MultLoop_acc_3209_nl;
  wire[18:0] MultLoop_acc_4402_nl;
  wire[19:0] nl_MultLoop_acc_4402_nl;
  wire[18:0] MultLoop_acc_4639_nl;
  wire[19:0] nl_MultLoop_acc_4639_nl;
  wire[19:0] MultLoop_acc_4403_nl;
  wire[20:0] nl_MultLoop_acc_4403_nl;
  wire[22:0] MultLoop_acc_4640_nl;
  wire[23:0] nl_MultLoop_acc_4640_nl;
  wire[20:0] MultLoop_acc_1180_nl;
  wire[21:0] nl_MultLoop_acc_1180_nl;
  wire[17:0] MultLoop_acc_3200_nl;
  wire[18:0] nl_MultLoop_acc_3200_nl;
  wire[12:0] MultLoop_acc_4399_nl;
  wire[13:0] nl_MultLoop_acc_4399_nl;
  wire[23:0] MultLoop_acc_1193_nl;
  wire[24:0] nl_MultLoop_acc_1193_nl;
  wire[20:0] MultLoop_acc_3205_nl;
  wire[21:0] nl_MultLoop_acc_3205_nl;
  wire[17:0] MultLoop_acc_3204_nl;
  wire[18:0] nl_MultLoop_acc_3204_nl;
  wire[17:0] MultLoop_acc_324_nl;
  wire[18:0] nl_MultLoop_acc_324_nl;
  wire[22:0] MultLoop_acc_1178_nl;
  wire[23:0] nl_MultLoop_acc_1178_nl;
  wire[17:0] MultLoop_acc_3202_nl;
  wire[18:0] nl_MultLoop_acc_3202_nl;
  wire[12:0] MultLoop_acc_4400_nl;
  wire[13:0] nl_MultLoop_acc_4400_nl;
  wire[20:0] MultLoop_acc_1176_nl;
  wire[21:0] nl_MultLoop_acc_1176_nl;
  wire[17:0] MultLoop_acc_3203_nl;
  wire[18:0] nl_MultLoop_acc_3203_nl;
  wire[18:0] MultLoop_acc_4641_nl;
  wire[19:0] nl_MultLoop_acc_4641_nl;
  wire[18:0] MultLoop_acc_4404_nl;
  wire[19:0] nl_MultLoop_acc_4404_nl;
  wire[21:0] MultLoop_acc_3217_nl;
  wire[23:0] nl_MultLoop_acc_3217_nl;
  wire[18:0] MultLoop_acc_4405_nl;
  wire[19:0] nl_MultLoop_acc_4405_nl;
  wire[19:0] MultLoop_acc_4642_nl;
  wire[20:0] nl_MultLoop_acc_4642_nl;
  wire[21:0] MultLoop_acc_1175_nl;
  wire[22:0] nl_MultLoop_acc_1175_nl;
  wire[20:0] MultLoop_acc_3221_nl;
  wire[21:0] nl_MultLoop_acc_3221_nl;
  wire[17:0] MultLoop_acc_3220_nl;
  wire[18:0] nl_MultLoop_acc_3220_nl;
  wire[22:0] MultLoop_acc_322_nl;
  wire[23:0] nl_MultLoop_acc_322_nl;
  wire[20:0] MultLoop_acc_3161_nl;
  wire[21:0] nl_MultLoop_acc_3161_nl;
  wire[22:0] MultLoop_acc_308_nl;
  wire[23:0] nl_MultLoop_acc_308_nl;
  wire[19:0] MultLoop_acc_1179_nl;
  wire[20:0] nl_MultLoop_acc_1179_nl;
  wire[17:0] MultLoop_acc_3162_nl;
  wire[18:0] nl_MultLoop_acc_3162_nl;
  wire[17:0] MultLoop_acc_310_nl;
  wire[18:0] nl_MultLoop_acc_310_nl;
  wire[7:0] MultLoop_acc_288_nl;
  wire[8:0] nl_MultLoop_acc_288_nl;
  wire[17:0] MultLoop_acc_4408_nl;
  wire[18:0] nl_MultLoop_acc_4408_nl;
  wire[19:0] MultLoop_acc_3164_nl;
  wire[20:0] nl_MultLoop_acc_3164_nl;
  wire[21:0] MultLoop_acc_1192_nl;
  wire[22:0] nl_MultLoop_acc_1192_nl;
  wire[19:0] MultLoop_acc_3166_nl;
  wire[20:0] nl_MultLoop_acc_3166_nl;
  wire[17:0] MultLoop_acc_321_nl;
  wire[18:0] nl_MultLoop_acc_321_nl;
  wire[24:0] MultLoop_acc_316_nl;
  wire[25:0] nl_MultLoop_acc_316_nl;
  wire[22:0] MultLoop_acc_3168_nl;
  wire[23:0] nl_MultLoop_acc_3168_nl;
  wire[19:0] MultLoop_acc_3167_nl;
  wire[20:0] nl_MultLoop_acc_3167_nl;
  wire[18:0] MultLoop_acc_4643_nl;
  wire[19:0] nl_MultLoop_acc_4643_nl;
  wire[22:0] MultLoop_acc_1194_nl;
  wire[23:0] nl_MultLoop_acc_1194_nl;
  wire[20:0] MultLoop_acc_3174_nl;
  wire[22:0] nl_MultLoop_acc_3174_nl;
  wire[21:0] MultLoop_acc_290_nl;
  wire[22:0] nl_MultLoop_acc_290_nl;
  wire[15:0] MultLoop_acc_4409_nl;
  wire[16:0] nl_MultLoop_acc_4409_nl;
  wire[17:0] MultLoop_acc_4411_nl;
  wire[18:0] nl_MultLoop_acc_4411_nl;
  wire[19:0] MultLoop_acc_3159_nl;
  wire[20:0] nl_MultLoop_acc_3159_nl;
  wire[12:0] MultLoop_acc_4410_nl;
  wire[13:0] nl_MultLoop_acc_4410_nl;
  wire[20:0] MultLoop_acc_4681_nl;
  wire[21:0] nl_MultLoop_acc_4681_nl;
  wire[24:0] MultLoop_acc_299_nl;
  wire[25:0] nl_MultLoop_acc_299_nl;
  wire[20:0] MultLoop_acc_3171_nl;
  wire[21:0] nl_MultLoop_acc_3171_nl;
  wire[24:0] MultLoop_acc_330_nl;
  wire[25:0] nl_MultLoop_acc_330_nl;
  wire[21:0] MultLoop_acc_3175_nl;
  wire[22:0] nl_MultLoop_acc_3175_nl;
  wire[25:0] MultLoop_acc_331_nl;
  wire[26:0] nl_MultLoop_acc_331_nl;
  wire[20:0] MultLoop_acc_3176_nl;
  wire[21:0] nl_MultLoop_acc_3176_nl;
  wire[25:0] MultLoop_acc_325_nl;
  wire[27:0] nl_MultLoop_acc_325_nl;
  wire[18:0] MultLoop_acc_4644_nl;
  wire[19:0] nl_MultLoop_acc_4644_nl;
  wire[23:0] MultLoop_acc_1189_nl;
  wire[24:0] nl_MultLoop_acc_1189_nl;
  wire[21:0] MultLoop_acc_3183_nl;
  wire[22:0] nl_MultLoop_acc_3183_nl;
  wire[22:0] MultLoop_acc_1187_nl;
  wire[23:0] nl_MultLoop_acc_1187_nl;
  wire[20:0] MultLoop_acc_3185_nl;
  wire[21:0] nl_MultLoop_acc_3185_nl;
  wire[17:0] MultLoop_acc_3184_nl;
  wire[18:0] nl_MultLoop_acc_3184_nl;
  wire[21:0] MultLoop_acc_1188_nl;
  wire[22:0] nl_MultLoop_acc_1188_nl;
  wire[23:0] MultLoop_acc_1185_nl;
  wire[24:0] nl_MultLoop_acc_1185_nl;
  wire[19:0] MultLoop_acc_3188_nl;
  wire[20:0] nl_MultLoop_acc_3188_nl;
  wire[18:0] MultLoop_acc_4682_nl;
  wire[19:0] nl_MultLoop_acc_4682_nl;
  wire[18:0] MultLoop_acc_4683_nl;
  wire[19:0] nl_MultLoop_acc_4683_nl;
  wire[25:0] MultLoop_acc_304_nl;
  wire[26:0] nl_MultLoop_acc_304_nl;
  wire[23:0] MultLoop_acc_3194_nl;
  wire[24:0] nl_MultLoop_acc_3194_nl;
  wire[17:0] MultLoop_acc_4414_nl;
  wire[18:0] nl_MultLoop_acc_4414_nl;
  wire[22:0] MultLoop_acc_3198_nl;
  wire[24:0] nl_MultLoop_acc_3198_nl;
  wire[16:0] MultLoop_772_MultLoop_acc_3_nl;
  wire[18:0] nl_MultLoop_772_MultLoop_acc_3_nl;
  wire[15:0] MultLoop_770_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_770_MultLoop_acc_3_nl;
  wire[13:0] MultLoop_acc_2262_nl;
  wire[14:0] nl_MultLoop_acc_2262_nl;
  wire[22:0] MultLoop_acc_760_nl;
  wire[23:0] nl_MultLoop_acc_760_nl;
  wire[23:0] MultLoop_acc_759_nl;
  wire[24:0] nl_MultLoop_acc_759_nl;
  wire[21:0] MultLoop_acc_2261_nl;
  wire[22:0] nl_MultLoop_acc_2261_nl;
  wire[25:0] MultLoop_acc_762_nl;
  wire[27:0] nl_MultLoop_acc_762_nl;
  wire[20:0] MultLoop_acc_1327_nl;
  wire[21:0] nl_MultLoop_acc_1327_nl;
  wire[25:0] MultLoop_acc_763_nl;
  wire[26:0] nl_MultLoop_acc_763_nl;
  wire[22:0] MultLoop_acc_2268_nl;
  wire[23:0] nl_MultLoop_acc_2268_nl;
  wire[19:0] MultLoop_acc_2267_nl;
  wire[20:0] nl_MultLoop_acc_2267_nl;
  wire[21:0] MultLoop_acc_780_nl;
  wire[22:0] nl_MultLoop_acc_780_nl;
  wire[19:0] MultLoop_acc_2192_nl;
  wire[20:0] nl_MultLoop_acc_2192_nl;
  wire[14:0] MultLoop_acc_4093_nl;
  wire[15:0] nl_MultLoop_acc_4093_nl;
  wire[20:0] MultLoop_acc_770_nl;
  wire[21:0] nl_MultLoop_acc_770_nl;
  wire[16:0] MultLoop_acc_4092_nl;
  wire[17:0] nl_MultLoop_acc_4092_nl;
  wire[18:0] MultLoop_acc_1330_nl;
  wire[19:0] nl_MultLoop_acc_1330_nl;
  wire[17:0] MultLoop_acc_779_nl;
  wire[18:0] nl_MultLoop_acc_779_nl;
  wire[18:0] MultLoop_acc_4617_nl;
  wire[19:0] nl_MultLoop_acc_4617_nl;
  wire[21:0] MultLoop_acc_1344_nl;
  wire[22:0] nl_MultLoop_acc_1344_nl;
  wire[18:0] MultLoop_acc_2194_nl;
  wire[19:0] nl_MultLoop_acc_2194_nl;
  wire[17:0] MultLoop_acc_792_nl;
  wire[18:0] nl_MultLoop_acc_792_nl;
  wire[21:0] MultLoop_acc_1338_nl;
  wire[22:0] nl_MultLoop_acc_1338_nl;
  wire[17:0] MultLoop_acc_2196_nl;
  wire[18:0] nl_MultLoop_acc_2196_nl;
  wire[23:0] MultLoop_acc_783_nl;
  wire[25:0] nl_MultLoop_acc_783_nl;
  wire[13:0] MultLoop_acc_4095_nl;
  wire[14:0] nl_MultLoop_acc_4095_nl;
  wire[24:0] MultLoop_acc_781_nl;
  wire[25:0] nl_MultLoop_acc_781_nl;
  wire[20:0] MultLoop_acc_2199_nl;
  wire[21:0] nl_MultLoop_acc_2199_nl;
  wire[17:0] MultLoop_acc_4098_nl;
  wire[18:0] nl_MultLoop_acc_4098_nl;
  wire[23:0] MultLoop_acc_2206_nl;
  wire[25:0] nl_MultLoop_acc_2206_nl;
  wire[22:0] MultLoop_acc_1334_nl;
  wire[23:0] nl_MultLoop_acc_1334_nl;
  wire[20:0] MultLoop_acc_2202_nl;
  wire[21:0] nl_MultLoop_acc_2202_nl;
  wire[17:0] MultLoop_acc_2201_nl;
  wire[18:0] nl_MultLoop_acc_2201_nl;
  wire[21:0] MultLoop_acc_1332_nl;
  wire[22:0] nl_MultLoop_acc_1332_nl;
  wire[17:0] MultLoop_acc_2203_nl;
  wire[18:0] nl_MultLoop_acc_2203_nl;
  wire[24:0] MultLoop_acc_802_nl;
  wire[25:0] nl_MultLoop_acc_802_nl;
  wire[21:0] MultLoop_acc_2209_nl;
  wire[22:0] nl_MultLoop_acc_2209_nl;
  wire[19:0] MultLoop_acc_2208_nl;
  wire[20:0] nl_MultLoop_acc_2208_nl;
  wire[21:0] MultLoop_acc_801_nl;
  wire[22:0] nl_MultLoop_acc_801_nl;
  wire[20:0] MultLoop_acc_2212_nl;
  wire[22:0] nl_MultLoop_acc_2212_nl;
  wire[24:0] MultLoop_acc_798_nl;
  wire[26:0] nl_MultLoop_acc_798_nl;
  wire[19:0] MultLoop_acc_1343_nl;
  wire[20:0] nl_MultLoop_acc_1343_nl;
  wire[17:0] MultLoop_acc_2216_nl;
  wire[18:0] nl_MultLoop_acc_2216_nl;
  wire[21:0] MultLoop_acc_1341_nl;
  wire[22:0] nl_MultLoop_acc_1341_nl;
  wire[17:0] MultLoop_acc_2218_nl;
  wire[18:0] nl_MultLoop_acc_2218_nl;
  wire[23:0] MultLoop_acc_1342_nl;
  wire[24:0] nl_MultLoop_acc_1342_nl;
  wire[20:0] MultLoop_acc_2221_nl;
  wire[21:0] nl_MultLoop_acc_2221_nl;
  wire[17:0] MultLoop_acc_4105_nl;
  wire[18:0] nl_MultLoop_acc_4105_nl;
  wire[23:0] MultLoop_acc_2224_nl;
  wire[25:0] nl_MultLoop_acc_2224_nl;
  wire[17:0] MultLoop_acc_4107_nl;
  wire[18:0] nl_MultLoop_acc_4107_nl;
  wire[21:0] MultLoop_acc_2227_nl;
  wire[23:0] nl_MultLoop_acc_2227_nl;
  wire[17:0] MultLoop_acc_4109_nl;
  wire[18:0] nl_MultLoop_acc_4109_nl;
  wire[21:0] MultLoop_acc_2230_nl;
  wire[23:0] nl_MultLoop_acc_2230_nl;
  wire[12:0] MultLoop_acc_4108_nl;
  wire[13:0] nl_MultLoop_acc_4108_nl;
  wire[20:0] MultLoop_acc_1337_nl;
  wire[21:0] nl_MultLoop_acc_1337_nl;
  wire[17:0] MultLoop_acc_2232_nl;
  wire[18:0] nl_MultLoop_acc_2232_nl;
  wire[18:0] MultLoop_acc_4618_nl;
  wire[19:0] nl_MultLoop_acc_4618_nl;
  wire[17:0] MultLoop_acc_4112_nl;
  wire[18:0] nl_MultLoop_acc_4112_nl;
  wire[22:0] MultLoop_acc_2237_nl;
  wire[24:0] nl_MultLoop_acc_2237_nl;
  wire[10:0] MultLoop_acc_4111_nl;
  wire[11:0] nl_MultLoop_acc_4111_nl;
  wire[17:0] MultLoop_acc_4114_nl;
  wire[18:0] nl_MultLoop_acc_4114_nl;
  wire[24:0] MultLoop_acc_2240_nl;
  wire[25:0] nl_MultLoop_acc_2240_nl;
  wire[21:0] MultLoop_acc_2239_nl;
  wire[22:0] nl_MultLoop_acc_2239_nl;
  wire[10:0] MultLoop_acc_4113_nl;
  wire[11:0] nl_MultLoop_acc_4113_nl;
  wire[25:0] MultLoop_acc_774_nl;
  wire[26:0] nl_MultLoop_acc_774_nl;
  wire[24:0] MultLoop_acc_2243_nl;
  wire[26:0] nl_MultLoop_acc_2243_nl;
  wire[24:0] MultLoop_acc_1340_nl;
  wire[25:0] nl_MultLoop_acc_1340_nl;
  wire[21:0] MultLoop_acc_2258_nl;
  wire[23:0] nl_MultLoop_acc_2258_nl;
  wire[23:0] MultLoop_acc_1329_nl;
  wire[24:0] nl_MultLoop_acc_1329_nl;
  wire[20:0] MultLoop_acc_2255_nl;
  wire[21:0] nl_MultLoop_acc_2255_nl;
  wire[17:0] MultLoop_acc_2254_nl;
  wire[18:0] nl_MultLoop_acc_2254_nl;
  wire[23:0] MultLoop_acc_1335_nl;
  wire[24:0] nl_MultLoop_acc_1335_nl;
  wire[22:0] MultLoop_acc_2246_nl;
  wire[24:0] nl_MultLoop_acc_2246_nl;
  wire[17:0] MultLoop_acc_2244_nl;
  wire[18:0] nl_MultLoop_acc_2244_nl;
  wire[22:0] MultLoop_acc_1333_nl;
  wire[23:0] nl_MultLoop_acc_1333_nl;
  wire[19:0] MultLoop_acc_2249_nl;
  wire[21:0] nl_MultLoop_acc_2249_nl;
  wire[11:0] MultLoop_acc_4115_nl;
  wire[12:0] nl_MultLoop_acc_4115_nl;
  wire[23:0] MultLoop_acc_1331_nl;
  wire[24:0] nl_MultLoop_acc_1331_nl;
  wire[17:0] MultLoop_acc_2251_nl;
  wire[18:0] nl_MultLoop_acc_2251_nl;
  wire[11:0] MultLoop_acc_4116_nl;
  wire[12:0] nl_MultLoop_acc_4116_nl;
  wire[19:0] MultLoop_acc_4118_nl;
  wire[20:0] nl_MultLoop_acc_4118_nl;
  wire[17:0] MultLoop_acc_4117_nl;
  wire[18:0] nl_MultLoop_acc_4117_nl;
  wire[18:0] MultLoop_acc_1336_nl;
  wire[19:0] nl_MultLoop_acc_1336_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl;
  wire[13:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl;
  wire[17:0] MultLoop_acc_767_nl;
  wire[18:0] nl_MultLoop_acc_767_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_6_nl;
  wire[17:0] MultLoop_acc_800_nl;
  wire[18:0] nl_MultLoop_acc_800_nl;
  wire[21:0] MultLoop_acc_1207_nl;
  wire[22:0] nl_MultLoop_acc_1207_nl;
  wire[20:0] MultLoop_acc_3097_nl;
  wire[21:0] nl_MultLoop_acc_3097_nl;
  wire[17:0] MultLoop_acc_3096_nl;
  wire[18:0] nl_MultLoop_acc_3096_nl;
  wire[22:0] MultLoop_acc_356_nl;
  wire[23:0] nl_MultLoop_acc_356_nl;
  wire[14:0] MultLoop_acc_4371_nl;
  wire[15:0] nl_MultLoop_acc_4371_nl;
  wire[20:0] MultLoop_acc_4636_nl;
  wire[21:0] nl_MultLoop_acc_4636_nl;
  wire[17:0] MultLoop_acc_4373_nl;
  wire[18:0] nl_MultLoop_acc_4373_nl;
  wire[21:0] MultLoop_acc_3101_nl;
  wire[22:0] nl_MultLoop_acc_3101_nl;
  wire[18:0] MultLoop_acc_1210_nl;
  wire[19:0] nl_MultLoop_acc_1210_nl;
  wire[18:0] MultLoop_acc_4637_nl;
  wire[19:0] nl_MultLoop_acc_4637_nl;
  wire[22:0] MultLoop_acc_376_nl;
  wire[23:0] nl_MultLoop_acc_376_nl;
  wire[20:0] MultLoop_acc_3104_nl;
  wire[21:0] nl_MultLoop_acc_3104_nl;
  wire[13:0] MultLoop_acc_4374_nl;
  wire[14:0] nl_MultLoop_acc_4374_nl;
  wire[22:0] MultLoop_acc_1201_nl;
  wire[23:0] nl_MultLoop_acc_1201_nl;
  wire[20:0] MultLoop_acc_3106_nl;
  wire[21:0] nl_MultLoop_acc_3106_nl;
  wire[22:0] MultLoop_acc_358_nl;
  wire[23:0] nl_MultLoop_acc_358_nl;
  wire[20:0] MultLoop_acc_3108_nl;
  wire[21:0] nl_MultLoop_acc_3108_nl;
  wire[13:0] MultLoop_acc_4375_nl;
  wire[14:0] nl_MultLoop_acc_4375_nl;
  wire[21:0] MultLoop_acc_1197_nl;
  wire[22:0] nl_MultLoop_acc_1197_nl;
  wire[20:0] MultLoop_acc_3110_nl;
  wire[21:0] nl_MultLoop_acc_3110_nl;
  wire[17:0] MultLoop_acc_3109_nl;
  wire[18:0] nl_MultLoop_acc_3109_nl;
  wire[21:0] MultLoop_acc_348_nl;
  wire[22:0] nl_MultLoop_acc_348_nl;
  wire[15:0] MultLoop_acc_4376_nl;
  wire[16:0] nl_MultLoop_acc_4376_nl;
  wire[20:0] MultLoop_acc_1196_nl;
  wire[21:0] nl_MultLoop_acc_1196_nl;
  wire[17:0] MultLoop_acc_3112_nl;
  wire[18:0] nl_MultLoop_acc_3112_nl;
  wire[17:0] MultLoop_acc_4378_nl;
  wire[18:0] nl_MultLoop_acc_4378_nl;
  wire[24:0] MultLoop_acc_3115_nl;
  wire[25:0] nl_MultLoop_acc_3115_nl;
  wire[21:0] MultLoop_acc_3114_nl;
  wire[22:0] nl_MultLoop_acc_3114_nl;
  wire[10:0] MultLoop_acc_4377_nl;
  wire[11:0] nl_MultLoop_acc_4377_nl;
  wire[17:0] MultLoop_acc_4380_nl;
  wire[18:0] nl_MultLoop_acc_4380_nl;
  wire[22:0] MultLoop_acc_3119_nl;
  wire[24:0] nl_MultLoop_acc_3119_nl;
  wire[17:0] MultLoop_acc_4382_nl;
  wire[18:0] nl_MultLoop_acc_4382_nl;
  wire[24:0] MultLoop_acc_3122_nl;
  wire[25:0] nl_MultLoop_acc_3122_nl;
  wire[21:0] MultLoop_acc_3121_nl;
  wire[22:0] nl_MultLoop_acc_3121_nl;
  wire[10:0] MultLoop_acc_4381_nl;
  wire[11:0] nl_MultLoop_acc_4381_nl;
  wire[23:0] MultLoop_acc_1205_nl;
  wire[24:0] nl_MultLoop_acc_1205_nl;
  wire[21:0] MultLoop_acc_3124_nl;
  wire[23:0] nl_MultLoop_acc_3124_nl;
  wire[22:0] MultLoop_acc_365_nl;
  wire[23:0] nl_MultLoop_acc_365_nl;
  wire[19:0] MultLoop_acc_3127_nl;
  wire[20:0] nl_MultLoop_acc_3127_nl;
  wire[17:0] MultLoop_acc_3126_nl;
  wire[18:0] nl_MultLoop_acc_3126_nl;
  wire[24:0] MultLoop_acc_366_nl;
  wire[25:0] nl_MultLoop_acc_366_nl;
  wire[21:0] MultLoop_acc_1203_nl;
  wire[22:0] nl_MultLoop_acc_1203_nl;
  wire[19:0] MultLoop_acc_3129_nl;
  wire[20:0] nl_MultLoop_acc_3129_nl;
  wire[24:0] MultLoop_acc_360_nl;
  wire[25:0] nl_MultLoop_acc_360_nl;
  wire[23:0] MultLoop_acc_3131_nl;
  wire[25:0] nl_MultLoop_acc_3131_nl;
  wire[21:0] MultLoop_acc_357_nl;
  wire[22:0] nl_MultLoop_acc_357_nl;
  wire[19:0] MultLoop_acc_3133_nl;
  wire[20:0] nl_MultLoop_acc_3133_nl;
  wire[14:0] MultLoop_acc_4384_nl;
  wire[15:0] nl_MultLoop_acc_4384_nl;
  wire[17:0] MultLoop_acc_4386_nl;
  wire[18:0] nl_MultLoop_acc_4386_nl;
  wire[23:0] MultLoop_acc_3136_nl;
  wire[24:0] nl_MultLoop_acc_3136_nl;
  wire[20:0] MultLoop_acc_3135_nl;
  wire[21:0] nl_MultLoop_acc_3135_nl;
  wire[17:0] MultLoop_acc_352_nl;
  wire[18:0] nl_MultLoop_acc_352_nl;
  wire[18:0] MultLoop_acc_1198_nl;
  wire[19:0] nl_MultLoop_acc_1198_nl;
  wire[18:0] MultLoop_acc_4638_nl;
  wire[19:0] nl_MultLoop_acc_4638_nl;
  wire[25:0] MultLoop_acc_349_nl;
  wire[27:0] nl_MultLoop_acc_349_nl;
  wire[11:0] MultLoop_acc_4387_nl;
  wire[12:0] nl_MultLoop_acc_4387_nl;
  wire[25:0] MultLoop_acc_346_nl;
  wire[27:0] nl_MultLoop_acc_346_nl;
  wire[20:0] MultLoop_acc_344_nl;
  wire[21:0] nl_MultLoop_acc_344_nl;
  wire[18:0] MultLoop_acc_3144_nl;
  wire[19:0] nl_MultLoop_acc_3144_nl;
  wire[25:0] MultLoop_acc_342_nl;
  wire[27:0] nl_MultLoop_acc_342_nl;
  wire[15:0] MultLoop_340_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_340_MultLoop_acc_3_nl;
  wire[14:0] MultLoop_acc_3154_nl;
  wire[15:0] nl_MultLoop_acc_3154_nl;
  wire[13:0] MultLoop_338_MultLoop_acc_3_nl;
  wire[14:0] nl_MultLoop_338_MultLoop_acc_3_nl;
  wire[11:0] MultLoop_acc_4392_nl;
  wire[12:0] nl_MultLoop_acc_4392_nl;
  wire[23:0] MultLoop_acc_337_nl;
  wire[24:0] nl_MultLoop_acc_337_nl;
  wire[13:0] MultLoop_acc_4393_nl;
  wire[14:0] nl_MultLoop_acc_4393_nl;
  wire[23:0] MultLoop_acc_1195_nl;
  wire[24:0] nl_MultLoop_acc_1195_nl;
  wire[21:0] MultLoop_acc_3153_nl;
  wire[22:0] nl_MultLoop_acc_3153_nl;
  wire[13:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl;
  wire[19:0] MultLoop_acc_345_nl;
  wire[20:0] nl_MultLoop_acc_345_nl;
  wire[18:0] MultLoop_acc_3094_nl;
  wire[19:0] nl_MultLoop_acc_3094_nl;
  wire[14:0] MultLoop_acc_4395_nl;
  wire[15:0] nl_MultLoop_acc_4395_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl;
  wire[13:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl;
  wire[20:0] MultLoop_acc_370_nl;
  wire[21:0] nl_MultLoop_acc_370_nl;
  wire[16:0] MultLoop_acc_4396_nl;
  wire[17:0] nl_MultLoop_acc_4396_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl;
  wire[20:0] MultLoop_acc_1209_nl;
  wire[21:0] nl_MultLoop_acc_1209_nl;
  wire[17:0] MultLoop_acc_3095_nl;
  wire[18:0] nl_MultLoop_acc_3095_nl;
  wire[26:0] MultLoop_acc_375_nl;
  wire[27:0] nl_MultLoop_acc_375_nl;
  wire[21:0] MultLoop_acc_1208_nl;
  wire[22:0] nl_MultLoop_acc_1208_nl;
  wire[17:0] MultLoop_acc_3157_nl;
  wire[18:0] nl_MultLoop_acc_3157_nl;
  wire[10:0] MultLoop_acc_4398_nl;
  wire[11:0] nl_MultLoop_acc_4398_nl;
  wire[24:0] MultLoop_acc_1319_nl;
  wire[25:0] nl_MultLoop_acc_1319_nl;
  wire[19:0] MultLoop_acc_2344_nl;
  wire[21:0] nl_MultLoop_acc_2344_nl;
  wire[21:0] MultLoop_acc_1318_nl;
  wire[22:0] nl_MultLoop_acc_1318_nl;
  wire[17:0] MultLoop_acc_2346_nl;
  wire[18:0] nl_MultLoop_acc_2346_nl;
  wire[12:0] MultLoop_acc_4123_nl;
  wire[13:0] nl_MultLoop_acc_4123_nl;
  wire[25:0] MultLoop_acc_724_nl;
  wire[27:0] nl_MultLoop_acc_724_nl;
  wire[13:0] MultLoop_acc_712_nl;
  wire[14:0] nl_MultLoop_acc_712_nl;
  wire[14:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl;
  wire[16:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl;
  wire[24:0] MultLoop_acc_727_nl;
  wire[26:0] nl_MultLoop_acc_727_nl;
  wire[22:0] MultLoop_acc_748_nl;
  wire[24:0] nl_MultLoop_acc_748_nl;
  wire[26:0] MultLoop_acc_720_nl;
  wire[28:0] nl_MultLoop_acc_720_nl;
  wire[10:0] MultLoop_acc_4125_nl;
  wire[11:0] nl_MultLoop_acc_4125_nl;
  wire[13:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl;
  wire[15:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl;
  wire[20:0] MultLoop_acc_716_nl;
  wire[21:0] nl_MultLoop_acc_716_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_5_nl;
  wire[20:0] MultLoop_acc_1326_nl;
  wire[21:0] nl_MultLoop_acc_1326_nl;
  wire[23:0] MultLoop_acc_751_nl;
  wire[25:0] nl_MultLoop_acc_751_nl;
  wire[13:0] MultLoop_acc_4126_nl;
  wire[14:0] nl_MultLoop_acc_4126_nl;
  wire[21:0] MultLoop_acc_743_nl;
  wire[22:0] nl_MultLoop_acc_743_nl;
  wire[19:0] MultLoop_acc_2277_nl;
  wire[20:0] nl_MultLoop_acc_2277_nl;
  wire[17:0] MultLoop_acc_2276_nl;
  wire[18:0] nl_MultLoop_acc_2276_nl;
  wire[12:0] MultLoop_acc_4127_nl;
  wire[13:0] nl_MultLoop_acc_4127_nl;
  wire[20:0] MultLoop_acc_740_nl;
  wire[21:0] nl_MultLoop_acc_740_nl;
  wire[16:0] MultLoop_acc_4128_nl;
  wire[17:0] nl_MultLoop_acc_4128_nl;
  wire[19:0] MultLoop_acc_733_nl;
  wire[20:0] nl_MultLoop_acc_733_nl;
  wire[18:0] MultLoop_acc_2280_nl;
  wire[19:0] nl_MultLoop_acc_2280_nl;
  wire[14:0] MultLoop_acc_4129_nl;
  wire[15:0] nl_MultLoop_acc_4129_nl;
  wire[23:0] MultLoop_acc_728_nl;
  wire[24:0] nl_MultLoop_acc_728_nl;
  wire[17:0] MultLoop_acc_4132_nl;
  wire[18:0] nl_MultLoop_acc_4132_nl;
  wire[19:0] MultLoop_acc_4669_nl;
  wire[20:0] nl_MultLoop_acc_4669_nl;
  wire[17:0] MultLoop_acc_4134_nl;
  wire[18:0] nl_MultLoop_acc_4134_nl;
  wire[22:0] MultLoop_acc_2288_nl;
  wire[23:0] nl_MultLoop_acc_2288_nl;
  wire[19:0] MultLoop_acc_2287_nl;
  wire[20:0] nl_MultLoop_acc_2287_nl;
  wire[23:0] MultLoop_acc_719_nl;
  wire[24:0] nl_MultLoop_acc_719_nl;
  wire[21:0] MultLoop_acc_2285_nl;
  wire[22:0] nl_MultLoop_acc_2285_nl;
  wire[21:0] MultLoop_acc_750_nl;
  wire[22:0] nl_MultLoop_acc_750_nl;
  wire[20:0] MultLoop_acc_2269_nl;
  wire[21:0] nl_MultLoop_acc_2269_nl;
  wire[18:0] MultLoop_acc_4619_nl;
  wire[19:0] nl_MultLoop_acc_4619_nl;
  wire[17:0] MultLoop_acc_4136_nl;
  wire[18:0] nl_MultLoop_acc_4136_nl;
  wire[22:0] MultLoop_acc_2292_nl;
  wire[23:0] nl_MultLoop_acc_2292_nl;
  wire[19:0] MultLoop_acc_2291_nl;
  wire[20:0] nl_MultLoop_acc_2291_nl;
  wire[22:0] MultLoop_acc_1323_nl;
  wire[23:0] nl_MultLoop_acc_1323_nl;
  wire[20:0] MultLoop_acc_2294_nl;
  wire[21:0] nl_MultLoop_acc_2294_nl;
  wire[23:0] MultLoop_acc_735_nl;
  wire[24:0] nl_MultLoop_acc_735_nl;
  wire[19:0] MultLoop_acc_757_nl;
  wire[20:0] nl_MultLoop_acc_757_nl;
  wire[18:0] MultLoop_acc_2303_nl;
  wire[19:0] nl_MultLoop_acc_2303_nl;
  wire[13:0] MultLoop_acc_4139_nl;
  wire[14:0] nl_MultLoop_acc_4139_nl;
  wire[20:0] MultLoop_acc_1320_nl;
  wire[21:0] nl_MultLoop_acc_1320_nl;
  wire[17:0] MultLoop_acc_2297_nl;
  wire[18:0] nl_MultLoop_acc_2297_nl;
  wire[13:0] MultLoop_acc_4138_nl;
  wire[14:0] nl_MultLoop_acc_4138_nl;
  wire[24:0] MultLoop_acc_731_nl;
  wire[25:0] nl_MultLoop_acc_731_nl;
  wire[23:0] MultLoop_acc_2299_nl;
  wire[25:0] nl_MultLoop_acc_2299_nl;
  wire[18:0] MultLoop_acc_4140_nl;
  wire[19:0] nl_MultLoop_acc_4140_nl;
  wire[20:0] MultLoop_acc_2304_nl;
  wire[21:0] nl_MultLoop_acc_2304_nl;
  wire[17:0] MultLoop_acc_4620_nl;
  wire[18:0] nl_MultLoop_acc_4620_nl;
  wire[19:0] MultLoop_acc_1325_nl;
  wire[20:0] nl_MultLoop_acc_1325_nl;
  wire[17:0] MultLoop_acc_4143_nl;
  wire[18:0] nl_MultLoop_acc_4143_nl;
  wire[22:0] MultLoop_acc_2310_nl;
  wire[24:0] nl_MultLoop_acc_2310_nl;
  wire[20:0] MultLoop_acc_747_nl;
  wire[21:0] nl_MultLoop_acc_747_nl;
  wire[16:0] MultLoop_acc_4144_nl;
  wire[17:0] nl_MultLoop_acc_4144_nl;
  wire[22:0] MultLoop_acc_745_nl;
  wire[23:0] nl_MultLoop_acc_745_nl;
  wire[20:0] MultLoop_acc_2314_nl;
  wire[22:0] nl_MultLoop_acc_2314_nl;
  wire[11:0] MultLoop_acc_4145_nl;
  wire[12:0] nl_MultLoop_acc_4145_nl;
  wire[19:0] MultLoop_acc_741_nl;
  wire[20:0] nl_MultLoop_acc_741_nl;
  wire[18:0] MultLoop_acc_2316_nl;
  wire[19:0] nl_MultLoop_acc_2316_nl;
  wire[18:0] MultLoop_acc_4621_nl;
  wire[19:0] nl_MultLoop_acc_4621_nl;
  wire[18:0] MultLoop_acc_1322_nl;
  wire[19:0] nl_MultLoop_acc_1322_nl;
  wire[17:0] MultLoop_acc_4148_nl;
  wire[18:0] nl_MultLoop_acc_4148_nl;
  wire[23:0] MultLoop_acc_2320_nl;
  wire[24:0] nl_MultLoop_acc_2320_nl;
  wire[19:0] MultLoop_acc_2319_nl;
  wire[20:0] nl_MultLoop_acc_2319_nl;
  wire[23:0] MultLoop_acc_734_nl;
  wire[25:0] nl_MultLoop_acc_734_nl;
  wire[22:0] MultLoop_acc_1316_nl;
  wire[23:0] nl_MultLoop_acc_1316_nl;
  wire[17:0] MultLoop_acc_2334_nl;
  wire[18:0] nl_MultLoop_acc_2334_nl;
  wire[24:0] MultLoop_acc_718_nl;
  wire[25:0] nl_MultLoop_acc_718_nl;
  wire[17:0] MultLoop_acc_4151_nl;
  wire[18:0] nl_MultLoop_acc_4151_nl;
  wire[21:0] MultLoop_acc_2325_nl;
  wire[22:0] nl_MultLoop_acc_2325_nl;
  wire[17:0] MultLoop_acc_2324_nl;
  wire[18:0] nl_MultLoop_acc_2324_nl;
  wire[20:0] MultLoop_acc_1317_nl;
  wire[21:0] nl_MultLoop_acc_1317_nl;
  wire[17:0] MultLoop_acc_2327_nl;
  wire[18:0] nl_MultLoop_acc_2327_nl;
  wire[12:0] MultLoop_acc_4152_nl;
  wire[13:0] nl_MultLoop_acc_4152_nl;
  wire[17:0] MultLoop_acc_4154_nl;
  wire[18:0] nl_MultLoop_acc_4154_nl;
  wire[20:0] MultLoop_acc_2330_nl;
  wire[21:0] nl_MultLoop_acc_2330_nl;
  wire[17:0] MultLoop_acc_2329_nl;
  wire[18:0] nl_MultLoop_acc_2329_nl;
  wire[24:0] MultLoop_acc_722_nl;
  wire[25:0] nl_MultLoop_acc_722_nl;
  wire[23:0] MultLoop_acc_2332_nl;
  wire[25:0] nl_MultLoop_acc_2332_nl;
  wire[22:0] MultLoop_acc_715_nl;
  wire[23:0] nl_MultLoop_acc_715_nl;
  wire[20:0] MultLoop_acc_2338_nl;
  wire[21:0] nl_MultLoop_acc_2338_nl;
  wire[17:0] MultLoop_acc_4159_nl;
  wire[18:0] nl_MultLoop_acc_4159_nl;
  wire[18:0] MultLoop_acc_4670_nl;
  wire[19:0] nl_MultLoop_acc_4670_nl;
  wire[17:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl;
  wire[19:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl;
  wire[26:0] MultLoop_acc_407_nl;
  wire[28:0] nl_MultLoop_acc_407_nl;
  wire[23:0] MultLoop_acc_404_nl;
  wire[25:0] nl_MultLoop_acc_404_nl;
  wire[25:0] MultLoop_acc_402_nl;
  wire[26:0] nl_MultLoop_acc_402_nl;
  wire[21:0] MultLoop_acc_3088_nl;
  wire[22:0] nl_MultLoop_acc_3088_nl;
  wire[19:0] MultLoop_acc_3087_nl;
  wire[20:0] nl_MultLoop_acc_3087_nl;
  wire[21:0] MultLoop_acc_398_nl;
  wire[22:0] nl_MultLoop_acc_398_nl;
  wire[15:0] MultLoop_acc_4350_nl;
  wire[16:0] nl_MultLoop_acc_4350_nl;
  wire[26:0] MultLoop_acc_419_nl;
  wire[28:0] nl_MultLoop_acc_419_nl;
  wire[26:0] MultLoop_acc_414_nl;
  wire[28:0] nl_MultLoop_acc_414_nl;
  wire[20:0] MultLoop_acc_1219_nl;
  wire[21:0] nl_MultLoop_acc_1219_nl;
  wire[17:0] MultLoop_acc_3078_nl;
  wire[18:0] nl_MultLoop_acc_3078_nl;
  wire[25:0] MultLoop_acc_409_nl;
  wire[27:0] nl_MultLoop_acc_409_nl;
  wire[22:0] MultLoop_acc_1215_nl;
  wire[23:0] nl_MultLoop_acc_1215_nl;
  wire[17:0] MultLoop_acc_3091_nl;
  wire[18:0] nl_MultLoop_acc_3091_nl;
  wire[17:0] MultLoop_acc_389_nl;
  wire[18:0] nl_MultLoop_acc_389_nl;
  wire[17:0] MultLoop_acc_4353_nl;
  wire[18:0] nl_MultLoop_acc_4353_nl;
  wire[21:0] MultLoop_acc_3026_nl;
  wire[22:0] nl_MultLoop_acc_3026_nl;
  wire[17:0] MultLoop_acc_4355_nl;
  wire[18:0] nl_MultLoop_acc_4355_nl;
  wire[18:0] MultLoop_acc_4679_nl;
  wire[19:0] nl_MultLoop_acc_4679_nl;
  wire[23:0] MultLoop_acc_405_nl;
  wire[24:0] nl_MultLoop_acc_405_nl;
  wire[22:0] MultLoop_acc_397_nl;
  wire[23:0] nl_MultLoop_acc_397_nl;
  wire[20:0] MultLoop_acc_3031_nl;
  wire[21:0] nl_MultLoop_acc_3031_nl;
  wire[21:0] MultLoop_acc_1212_nl;
  wire[22:0] nl_MultLoop_acc_1212_nl;
  wire[17:0] MultLoop_acc_3033_nl;
  wire[18:0] nl_MultLoop_acc_3033_nl;
  wire[13:0] MultLoop_acc_4357_nl;
  wire[14:0] nl_MultLoop_acc_4357_nl;
  wire[18:0] MultLoop_acc_1226_nl;
  wire[19:0] nl_MultLoop_acc_1226_nl;
  wire[21:0] MultLoop_acc_1223_nl;
  wire[22:0] nl_MultLoop_acc_1223_nl;
  wire[17:0] MultLoop_acc_3034_nl;
  wire[18:0] nl_MultLoop_acc_3034_nl;
  wire[20:0] MultLoop_acc_1224_nl;
  wire[21:0] nl_MultLoop_acc_1224_nl;
  wire[17:0] MultLoop_acc_3035_nl;
  wire[18:0] nl_MultLoop_acc_3035_nl;
  wire[19:0] MultLoop_acc_1221_nl;
  wire[20:0] nl_MultLoop_acc_1221_nl;
  wire[17:0] MultLoop_acc_3036_nl;
  wire[18:0] nl_MultLoop_acc_3036_nl;
  wire[20:0] MultLoop_acc_403_nl;
  wire[21:0] nl_MultLoop_acc_403_nl;
  wire[18:0] MultLoop_acc_3038_nl;
  wire[19:0] nl_MultLoop_acc_3038_nl;
  wire[24:0] MultLoop_acc_393_nl;
  wire[25:0] nl_MultLoop_acc_393_nl;
  wire[23:0] MultLoop_acc_3040_nl;
  wire[24:0] nl_MultLoop_acc_3040_nl;
  wire[20:0] MultLoop_acc_1213_nl;
  wire[21:0] nl_MultLoop_acc_1213_nl;
  wire[17:0] MultLoop_acc_3042_nl;
  wire[18:0] nl_MultLoop_acc_3042_nl;
  wire[14:0] MultLoop_acc_4359_nl;
  wire[15:0] nl_MultLoop_acc_4359_nl;
  wire[21:0] MultLoop_acc_390_nl;
  wire[22:0] nl_MultLoop_acc_390_nl;
  wire[18:0] MultLoop_acc_3044_nl;
  wire[19:0] nl_MultLoop_acc_3044_nl;
  wire[23:0] MultLoop_acc_1228_nl;
  wire[24:0] nl_MultLoop_acc_1228_nl;
  wire[20:0] MultLoop_acc_3053_nl;
  wire[21:0] nl_MultLoop_acc_3053_nl;
  wire[17:0] MultLoop_acc_4362_nl;
  wire[18:0] nl_MultLoop_acc_4362_nl;
  wire[23:0] MultLoop_acc_3047_nl;
  wire[24:0] nl_MultLoop_acc_3047_nl;
  wire[19:0] MultLoop_acc_3046_nl;
  wire[20:0] nl_MultLoop_acc_3046_nl;
  wire[24:0] MultLoop_acc_382_nl;
  wire[25:0] nl_MultLoop_acc_382_nl;
  wire[21:0] MultLoop_acc_3050_nl;
  wire[22:0] nl_MultLoop_acc_3050_nl;
  wire[19:0] MultLoop_acc_3049_nl;
  wire[20:0] nl_MultLoop_acc_3049_nl;
  wire[17:0] MultLoop_acc_4366_nl;
  wire[18:0] nl_MultLoop_acc_4366_nl;
  wire[20:0] MultLoop_acc_3055_nl;
  wire[21:0] nl_MultLoop_acc_3055_nl;
  wire[22:0] MultLoop_acc_1220_nl;
  wire[23:0] nl_MultLoop_acc_1220_nl;
  wire[20:0] MultLoop_acc_3057_nl;
  wire[21:0] nl_MultLoop_acc_3057_nl;
  wire[18:0] MultLoop_acc_1218_nl;
  wire[19:0] nl_MultLoop_acc_1218_nl;
  wire[22:0] MultLoop_acc_401_nl;
  wire[23:0] nl_MultLoop_acc_401_nl;
  wire[20:0] MultLoop_acc_3060_nl;
  wire[21:0] nl_MultLoop_acc_3060_nl;
  wire[17:0] MultLoop_acc_3059_nl;
  wire[18:0] nl_MultLoop_acc_3059_nl;
  wire[18:0] MultLoop_acc_4680_nl;
  wire[19:0] nl_MultLoop_acc_4680_nl;
  wire[26:0] MultLoop_acc_423_nl;
  wire[28:0] nl_MultLoop_acc_423_nl;
  wire[17:0] MultLoop_acc_4369_nl;
  wire[18:0] nl_MultLoop_acc_4369_nl;
  wire[24:0] MultLoop_acc_3067_nl;
  wire[25:0] nl_MultLoop_acc_3067_nl;
  wire[20:0] MultLoop_acc_3066_nl;
  wire[21:0] nl_MultLoop_acc_3066_nl;
  wire[22:0] MultLoop_acc_1214_nl;
  wire[23:0] nl_MultLoop_acc_1214_nl;
  wire[18:0] MultLoop_acc_4635_nl;
  wire[19:0] nl_MultLoop_acc_4635_nl;
  wire[17:0] MultLoop_acc_385_nl;
  wire[18:0] nl_MultLoop_acc_385_nl;
  wire[17:0] MultLoop_acc_428_nl;
  wire[18:0] nl_MultLoop_acc_428_nl;
  wire[18:0] MultLoop_acc_1222_nl;
  wire[19:0] nl_MultLoop_acc_1222_nl;
  wire[17:0] MultLoop_acc_386_nl;
  wire[18:0] nl_MultLoop_acc_386_nl;
  wire[10:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl;
  wire[11:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl;
  wire[23:0] MultLoop_acc_1307_nl;
  wire[24:0] nl_MultLoop_acc_1307_nl;
  wire[17:0] MultLoop_acc_2411_nl;
  wire[18:0] nl_MultLoop_acc_2411_nl;
  wire[22:0] MultLoop_acc_1305_nl;
  wire[23:0] nl_MultLoop_acc_1305_nl;
  wire[20:0] MultLoop_acc_2413_nl;
  wire[21:0] nl_MultLoop_acc_2413_nl;
  wire[17:0] MultLoop_acc_4161_nl;
  wire[18:0] nl_MultLoop_acc_4161_nl;
  wire[21:0] MultLoop_acc_2408_nl;
  wire[23:0] nl_MultLoop_acc_2408_nl;
  wire[17:0] MultLoop_acc_2406_nl;
  wire[18:0] nl_MultLoop_acc_2406_nl;
  wire[23:0] MultLoop_acc_4671_nl;
  wire[24:0] nl_MultLoop_acc_4671_nl;
  wire[24:0] MultLoop_acc_682_nl;
  wire[25:0] nl_MultLoop_acc_682_nl;
  wire[23:0] MultLoop_acc_1306_nl;
  wire[24:0] nl_MultLoop_acc_1306_nl;
  wire[22:0] MultLoop_acc_2416_nl;
  wire[23:0] nl_MultLoop_acc_2416_nl;
  wire[19:0] MultLoop_acc_2415_nl;
  wire[21:0] nl_MultLoop_acc_2415_nl;
  wire[17:0] MultLoop_acc_4164_nl;
  wire[18:0] nl_MultLoop_acc_4164_nl;
  wire[21:0] MultLoop_acc_2418_nl;
  wire[22:0] nl_MultLoop_acc_2418_nl;
  wire[23:0] MultLoop_acc_1310_nl;
  wire[24:0] nl_MultLoop_acc_1310_nl;
  wire[19:0] MultLoop_acc_2425_nl;
  wire[20:0] nl_MultLoop_acc_2425_nl;
  wire[18:0] MultLoop_acc_4168_nl;
  wire[19:0] nl_MultLoop_acc_4168_nl;
  wire[24:0] MultLoop_acc_677_nl;
  wire[25:0] nl_MultLoop_acc_677_nl;
  wire[20:0] MultLoop_acc_2427_nl;
  wire[21:0] nl_MultLoop_acc_2427_nl;
  wire[21:0] MultLoop_acc_1303_nl;
  wire[22:0] nl_MultLoop_acc_1303_nl;
  wire[17:0] MultLoop_acc_4166_nl;
  wire[18:0] nl_MultLoop_acc_4166_nl;
  wire[22:0] MultLoop_acc_2422_nl;
  wire[23:0] nl_MultLoop_acc_2422_nl;
  wire[19:0] MultLoop_acc_2421_nl;
  wire[20:0] nl_MultLoop_acc_2421_nl;
  wire[26:0] MultLoop_acc_663_nl;
  wire[28:0] nl_MultLoop_acc_663_nl;
  wire[10:0] MultLoop_acc_4169_nl;
  wire[11:0] nl_MultLoop_acc_4169_nl;
  wire[17:0] MultLoop_acc_694_nl;
  wire[18:0] nl_MultLoop_acc_694_nl;
  wire[19:0] MultLoop_acc_665_nl;
  wire[20:0] nl_MultLoop_acc_665_nl;
  wire[18:0] MultLoop_acc_2353_nl;
  wire[19:0] nl_MultLoop_acc_2353_nl;
  wire[13:0] MultLoop_acc_4170_nl;
  wire[14:0] nl_MultLoop_acc_4170_nl;
  wire[17:0] MultLoop_acc_698_nl;
  wire[18:0] nl_MultLoop_acc_698_nl;
  wire[17:0] MultLoop_acc_4172_nl;
  wire[18:0] nl_MultLoop_acc_4172_nl;
  wire[20:0] MultLoop_acc_2355_nl;
  wire[21:0] nl_MultLoop_acc_2355_nl;
  wire[18:0] MultLoop_acc_1304_nl;
  wire[19:0] nl_MultLoop_acc_1304_nl;
  wire[22:0] MultLoop_acc_1314_nl;
  wire[23:0] nl_MultLoop_acc_1314_nl;
  wire[19:0] MultLoop_acc_2357_nl;
  wire[20:0] nl_MultLoop_acc_2357_nl;
  wire[17:0] MultLoop_acc_2356_nl;
  wire[18:0] nl_MultLoop_acc_2356_nl;
  wire[24:0] MultLoop_acc_703_nl;
  wire[25:0] nl_MultLoop_acc_703_nl;
  wire[21:0] MultLoop_acc_2360_nl;
  wire[22:0] nl_MultLoop_acc_2360_nl;
  wire[19:0] MultLoop_acc_2359_nl;
  wire[20:0] nl_MultLoop_acc_2359_nl;
  wire[19:0] MultLoop_acc_704_nl;
  wire[20:0] nl_MultLoop_acc_704_nl;
  wire[18:0] MultLoop_acc_2362_nl;
  wire[19:0] nl_MultLoop_acc_2362_nl;
  wire[24:0] MultLoop_acc_690_nl;
  wire[26:0] nl_MultLoop_acc_690_nl;
  wire[23:0] MultLoop_acc_680_nl;
  wire[24:0] nl_MultLoop_acc_680_nl;
  wire[21:0] MultLoop_acc_2366_nl;
  wire[22:0] nl_MultLoop_acc_2366_nl;
  wire[24:0] MultLoop_acc_681_nl;
  wire[25:0] nl_MultLoop_acc_681_nl;
  wire[21:0] MultLoop_acc_2369_nl;
  wire[22:0] nl_MultLoop_acc_2369_nl;
  wire[19:0] MultLoop_acc_2368_nl;
  wire[20:0] nl_MultLoop_acc_2368_nl;
  wire[12:0] MultLoop_acc_4176_nl;
  wire[13:0] nl_MultLoop_acc_4176_nl;
  wire[18:0] MultLoop_acc_4622_nl;
  wire[19:0] nl_MultLoop_acc_4622_nl;
  wire[17:0] MultLoop_acc_4178_nl;
  wire[18:0] nl_MultLoop_acc_4178_nl;
  wire[22:0] MultLoop_acc_2373_nl;
  wire[23:0] nl_MultLoop_acc_2373_nl;
  wire[19:0] MultLoop_acc_2372_nl;
  wire[20:0] nl_MultLoop_acc_2372_nl;
  wire[17:0] MultLoop_acc_675_nl;
  wire[18:0] nl_MultLoop_acc_675_nl;
  wire[17:0] MultLoop_acc_673_nl;
  wire[18:0] nl_MultLoop_acc_673_nl;
  wire[10:0] MultLoop_acc_4179_nl;
  wire[11:0] nl_MultLoop_acc_4179_nl;
  wire[20:0] MultLoop_acc_678_nl;
  wire[21:0] nl_MultLoop_acc_678_nl;
  wire[16:0] MultLoop_acc_4180_nl;
  wire[17:0] nl_MultLoop_acc_4180_nl;
  wire[21:0] MultLoop_acc_709_nl;
  wire[22:0] nl_MultLoop_acc_709_nl;
  wire[19:0] MultLoop_acc_2376_nl;
  wire[20:0] nl_MultLoop_acc_2376_nl;
  wire[17:0] MultLoop_acc_708_nl;
  wire[18:0] nl_MultLoop_acc_708_nl;
  wire[21:0] MultLoop_acc_706_nl;
  wire[22:0] nl_MultLoop_acc_706_nl;
  wire[19:0] MultLoop_acc_2379_nl;
  wire[20:0] nl_MultLoop_acc_2379_nl;
  wire[17:0] MultLoop_acc_2378_nl;
  wire[18:0] nl_MultLoop_acc_2378_nl;
  wire[10:0] MultLoop_acc_4182_nl;
  wire[11:0] nl_MultLoop_acc_4182_nl;
  wire[20:0] MultLoop_acc_1313_nl;
  wire[21:0] nl_MultLoop_acc_1313_nl;
  wire[17:0] MultLoop_acc_2380_nl;
  wire[18:0] nl_MultLoop_acc_2380_nl;
  wire[25:0] MultLoop_acc_702_nl;
  wire[27:0] nl_MultLoop_acc_702_nl;
  wire[18:0] MultLoop_acc_4623_nl;
  wire[19:0] nl_MultLoop_acc_4623_nl;
  wire[24:0] MultLoop_acc_700_nl;
  wire[25:0] nl_MultLoop_acc_700_nl;
  wire[23:0] MultLoop_acc_2386_nl;
  wire[24:0] nl_MultLoop_acc_2386_nl;
  wire[25:0] MultLoop_acc_696_nl;
  wire[26:0] nl_MultLoop_acc_696_nl;
  wire[24:0] MultLoop_acc_2389_nl;
  wire[26:0] nl_MultLoop_acc_2389_nl;
  wire[25:0] MultLoop_acc_695_nl;
  wire[26:0] nl_MultLoop_acc_695_nl;
  wire[22:0] MultLoop_acc_2391_nl;
  wire[23:0] nl_MultLoop_acc_2391_nl;
  wire[22:0] MultLoop_acc_692_nl;
  wire[23:0] nl_MultLoop_acc_692_nl;
  wire[21:0] MultLoop_acc_2394_nl;
  wire[23:0] nl_MultLoop_acc_2394_nl;
  wire[25:0] MultLoop_acc_691_nl;
  wire[26:0] nl_MultLoop_acc_691_nl;
  wire[17:0] MultLoop_acc_4187_nl;
  wire[18:0] nl_MultLoop_acc_4187_nl;
  wire[22:0] MultLoop_acc_2399_nl;
  wire[23:0] nl_MultLoop_acc_2399_nl;
  wire[19:0] MultLoop_acc_2398_nl;
  wire[20:0] nl_MultLoop_acc_2398_nl;
  wire[17:0] MultLoop_acc_2397_nl;
  wire[18:0] nl_MultLoop_acc_2397_nl;
  wire[22:0] MultLoop_acc_689_nl;
  wire[23:0] nl_MultLoop_acc_689_nl;
  wire[20:0] MultLoop_acc_2402_nl;
  wire[22:0] nl_MultLoop_acc_2402_nl;
  wire[22:0] MultLoop_acc_1309_nl;
  wire[23:0] nl_MultLoop_acc_1309_nl;
  wire[19:0] MultLoop_acc_2404_nl;
  wire[20:0] nl_MultLoop_acc_2404_nl;
  wire[26:0] MultLoop_acc_465_nl;
  wire[27:0] nl_MultLoop_acc_465_nl;
  wire[18:0] MultLoop_acc_4314_nl;
  wire[19:0] nl_MultLoop_acc_4314_nl;
  wire[20:0] MultLoop_acc_4634_nl;
  wire[21:0] nl_MultLoop_acc_4634_nl;
  wire[24:0] MultLoop_acc_1234_nl;
  wire[25:0] nl_MultLoop_acc_1234_nl;
  wire[21:0] MultLoop_acc_2969_nl;
  wire[22:0] nl_MultLoop_acc_2969_nl;
  wire[19:0] MultLoop_acc_2968_nl;
  wire[20:0] nl_MultLoop_acc_2968_nl;
  wire[22:0] MultLoop_acc_455_nl;
  wire[23:0] nl_MultLoop_acc_455_nl;
  wire[14:0] MultLoop_acc_4315_nl;
  wire[15:0] nl_MultLoop_acc_4315_nl;
  wire[16:0] MultLoop_434_MultLoop_acc_3_nl;
  wire[17:0] nl_MultLoop_434_MultLoop_acc_3_nl;
  wire[15:0] MultLoop_acc_2976_nl;
  wire[16:0] nl_MultLoop_acc_2976_nl;
  wire[22:0] MultLoop_acc_430_nl;
  wire[23:0] nl_MultLoop_acc_430_nl;
  wire[20:0] MultLoop_acc_2973_nl;
  wire[22:0] nl_MultLoop_acc_2973_nl;
  wire[11:0] MultLoop_acc_4316_nl;
  wire[12:0] nl_MultLoop_acc_4316_nl;
  wire[25:0] MultLoop_acc_429_nl;
  wire[27:0] nl_MultLoop_acc_429_nl;
  wire[11:0] MultLoop_acc_4317_nl;
  wire[12:0] nl_MultLoop_acc_4317_nl;
  wire[23:0] MultLoop_acc_1229_nl;
  wire[24:0] nl_MultLoop_acc_1229_nl;
  wire[19:0] MultLoop_acc_2979_nl;
  wire[20:0] nl_MultLoop_acc_2979_nl;
  wire[17:0] MultLoop_acc_4320_nl;
  wire[18:0] nl_MultLoop_acc_4320_nl;
  wire[17:0] MultLoop_acc_4322_nl;
  wire[18:0] nl_MultLoop_acc_4322_nl;
  wire[21:0] MultLoop_acc_2909_nl;
  wire[23:0] nl_MultLoop_acc_2909_nl;
  wire[12:0] MultLoop_acc_4321_nl;
  wire[13:0] nl_MultLoop_acc_4321_nl;
  wire[21:0] MultLoop_acc_462_nl;
  wire[22:0] nl_MultLoop_acc_462_nl;
  wire[20:0] MultLoop_acc_2912_nl;
  wire[22:0] nl_MultLoop_acc_2912_nl;
  wire[17:0] MultLoop_acc_474_nl;
  wire[18:0] nl_MultLoop_acc_474_nl;
  wire[20:0] MultLoop_acc_1231_nl;
  wire[21:0] nl_MultLoop_acc_1231_nl;
  wire[17:0] MultLoop_acc_2913_nl;
  wire[18:0] nl_MultLoop_acc_2913_nl;
  wire[20:0] MultLoop_acc_440_nl;
  wire[21:0] nl_MultLoop_acc_440_nl;
  wire[18:0] MultLoop_acc_2915_nl;
  wire[19:0] nl_MultLoop_acc_2915_nl;
  wire[12:0] MultLoop_acc_4324_nl;
  wire[13:0] nl_MultLoop_acc_4324_nl;
  wire[22:0] MultLoop_acc_472_nl;
  wire[23:0] nl_MultLoop_acc_472_nl;
  wire[19:0] MultLoop_acc_2917_nl;
  wire[20:0] nl_MultLoop_acc_2917_nl;
  wire[13:0] MultLoop_acc_4325_nl;
  wire[14:0] nl_MultLoop_acc_4325_nl;
  wire[21:0] MultLoop_acc_1238_nl;
  wire[22:0] nl_MultLoop_acc_1238_nl;
  wire[17:0] MultLoop_acc_2919_nl;
  wire[18:0] nl_MultLoop_acc_2919_nl;
  wire[12:0] MultLoop_acc_4326_nl;
  wire[13:0] nl_MultLoop_acc_4326_nl;
  wire[24:0] MultLoop_acc_467_nl;
  wire[25:0] nl_MultLoop_acc_467_nl;
  wire[21:0] MultLoop_acc_2921_nl;
  wire[22:0] nl_MultLoop_acc_2921_nl;
  wire[24:0] MultLoop_acc_460_nl;
  wire[25:0] nl_MultLoop_acc_460_nl;
  wire[24:0] MultLoop_acc_456_nl;
  wire[26:0] nl_MultLoop_acc_456_nl;
  wire[24:0] MultLoop_acc_450_nl;
  wire[25:0] nl_MultLoop_acc_450_nl;
  wire[23:0] MultLoop_acc_2926_nl;
  wire[24:0] nl_MultLoop_acc_2926_nl;
  wire[24:0] MultLoop_acc_446_nl;
  wire[25:0] nl_MultLoop_acc_446_nl;
  wire[20:0] MultLoop_acc_2927_nl;
  wire[21:0] nl_MultLoop_acc_2927_nl;
  wire[22:0] MultLoop_acc_1230_nl;
  wire[23:0] nl_MultLoop_acc_1230_nl;
  wire[17:0] MultLoop_acc_2929_nl;
  wire[18:0] nl_MultLoop_acc_2929_nl;
  wire[12:0] MultLoop_acc_4328_nl;
  wire[13:0] nl_MultLoop_acc_4328_nl;
  wire[22:0] MultLoop_acc_437_nl;
  wire[23:0] nl_MultLoop_acc_437_nl;
  wire[19:0] MultLoop_acc_2930_nl;
  wire[20:0] nl_MultLoop_acc_2930_nl;
  wire[24:0] MultLoop_acc_438_nl;
  wire[25:0] nl_MultLoop_acc_438_nl;
  wire[21:0] MultLoop_acc_2933_nl;
  wire[22:0] nl_MultLoop_acc_2933_nl;
  wire[19:0] MultLoop_acc_2932_nl;
  wire[20:0] nl_MultLoop_acc_2932_nl;
  wire[24:0] MultLoop_acc_436_nl;
  wire[25:0] nl_MultLoop_acc_436_nl;
  wire[22:0] MultLoop_acc_2934_nl;
  wire[23:0] nl_MultLoop_acc_2934_nl;
  wire[21:0] MultLoop_acc_1233_nl;
  wire[22:0] nl_MultLoop_acc_1233_nl;
  wire[20:0] MultLoop_acc_2945_nl;
  wire[21:0] nl_MultLoop_acc_2945_nl;
  wire[17:0] MultLoop_acc_2944_nl;
  wire[18:0] nl_MultLoop_acc_2944_nl;
  wire[17:0] MultLoop_acc_4333_nl;
  wire[18:0] nl_MultLoop_acc_4333_nl;
  wire[21:0] MultLoop_acc_2947_nl;
  wire[22:0] nl_MultLoop_acc_2947_nl;
  wire[25:0] MultLoop_acc_473_nl;
  wire[26:0] nl_MultLoop_acc_473_nl;
  wire[22:0] MultLoop_acc_2938_nl;
  wire[23:0] nl_MultLoop_acc_2938_nl;
  wire[20:0] MultLoop_acc_2937_nl;
  wire[21:0] nl_MultLoop_acc_2937_nl;
  wire[23:0] MultLoop_acc_1236_nl;
  wire[24:0] nl_MultLoop_acc_1236_nl;
  wire[21:0] MultLoop_acc_2940_nl;
  wire[22:0] nl_MultLoop_acc_2940_nl;
  wire[17:0] MultLoop_acc_2939_nl;
  wire[18:0] nl_MultLoop_acc_2939_nl;
  wire[22:0] MultLoop_acc_453_nl;
  wire[23:0] nl_MultLoop_acc_453_nl;
  wire[21:0] MultLoop_acc_2943_nl;
  wire[23:0] nl_MultLoop_acc_2943_nl;
  wire[17:0] MultLoop_acc_452_nl;
  wire[18:0] nl_MultLoop_acc_452_nl;
  wire[18:0] MultLoop_acc_4334_nl;
  wire[19:0] nl_MultLoop_acc_4334_nl;
  wire[21:0] MultLoop_acc_2948_nl;
  wire[22:0] nl_MultLoop_acc_2948_nl;
  wire[17:0] MultLoop_acc_448_nl;
  wire[18:0] nl_MultLoop_acc_448_nl;
  wire[25:0] MultLoop_acc_445_nl;
  wire[27:0] nl_MultLoop_acc_445_nl;
  wire[22:0] MultLoop_acc_1232_nl;
  wire[23:0] nl_MultLoop_acc_1232_nl;
  wire[19:0] MultLoop_acc_2952_nl;
  wire[21:0] nl_MultLoop_acc_2952_nl;
  wire[17:0] MultLoop_acc_4337_nl;
  wire[18:0] nl_MultLoop_acc_4337_nl;
  wire[24:0] MultLoop_acc_2955_nl;
  wire[25:0] nl_MultLoop_acc_2955_nl;
  wire[19:0] MultLoop_acc_2954_nl;
  wire[20:0] nl_MultLoop_acc_2954_nl;
  wire[22:0] MultLoop_acc_441_nl;
  wire[23:0] nl_MultLoop_acc_441_nl;
  wire[21:0] MultLoop_acc_2958_nl;
  wire[23:0] nl_MultLoop_acc_2958_nl;
  wire[22:0] MultLoop_acc_433_nl;
  wire[23:0] nl_MultLoop_acc_433_nl;
  wire[20:0] MultLoop_acc_2961_nl;
  wire[21:0] nl_MultLoop_acc_2961_nl;
  wire[17:0] MultLoop_acc_4341_nl;
  wire[18:0] nl_MultLoop_acc_4341_nl;
  wire[20:0] MultLoop_acc_2963_nl;
  wire[21:0] nl_MultLoop_acc_2963_nl;
  wire[19:0] MultLoop_acc_466_nl;
  wire[20:0] nl_MultLoop_acc_466_nl;
  wire[18:0] MultLoop_acc_2904_nl;
  wire[19:0] nl_MultLoop_acc_2904_nl;
  wire[13:0] MultLoop_acc_4342_nl;
  wire[14:0] nl_MultLoop_acc_4342_nl;
  wire[23:0] MultLoop_acc_1293_nl;
  wire[24:0] nl_MultLoop_acc_1293_nl;
  wire[19:0] MultLoop_acc_2551_nl;
  wire[21:0] nl_MultLoop_acc_2551_nl;
  wire[23:0] MultLoop_acc_1292_nl;
  wire[24:0] nl_MultLoop_acc_1292_nl;
  wire[20:0] MultLoop_acc_2554_nl;
  wire[22:0] nl_MultLoop_acc_2554_nl;
  wire[23:0] MultLoop_acc_1291_nl;
  wire[24:0] nl_MultLoop_acc_1291_nl;
  wire[19:0] MultLoop_acc_2557_nl;
  wire[21:0] nl_MultLoop_acc_2557_nl;
  wire[15:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl;
  wire[17:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl;
  wire[20:0] MultLoop_acc_659_nl;
  wire[21:0] nl_MultLoop_acc_659_nl;
  wire[18:0] MultLoop_acc_2480_nl;
  wire[19:0] nl_MultLoop_acc_2480_nl;
  wire[13:0] MultLoop_acc_4192_nl;
  wire[14:0] nl_MultLoop_acc_4192_nl;
  wire[23:0] MultLoop_acc_654_nl;
  wire[24:0] nl_MultLoop_acc_654_nl;
  wire[20:0] MultLoop_acc_2481_nl;
  wire[21:0] nl_MultLoop_acc_2481_nl;
  wire[21:0] MultLoop_acc_655_nl;
  wire[22:0] nl_MultLoop_acc_655_nl;
  wire[19:0] MultLoop_acc_2484_nl;
  wire[20:0] nl_MultLoop_acc_2484_nl;
  wire[17:0] MultLoop_acc_2483_nl;
  wire[18:0] nl_MultLoop_acc_2483_nl;
  wire[22:0] MultLoop_acc_644_nl;
  wire[23:0] nl_MultLoop_acc_644_nl;
  wire[14:0] MultLoop_acc_4194_nl;
  wire[15:0] nl_MultLoop_acc_4194_nl;
  wire[17:0] MultLoop_acc_645_nl;
  wire[18:0] nl_MultLoop_acc_645_nl;
  wire[22:0] MultLoop_acc_639_nl;
  wire[23:0] nl_MultLoop_acc_639_nl;
  wire[14:0] MultLoop_acc_4195_nl;
  wire[15:0] nl_MultLoop_acc_4195_nl;
  wire[18:0] MultLoop_acc_1301_nl;
  wire[19:0] nl_MultLoop_acc_1301_nl;
  wire[22:0] MultLoop_acc_4672_nl;
  wire[23:0] nl_MultLoop_acc_4672_nl;
  wire[22:0] MultLoop_acc_657_nl;
  wire[23:0] nl_MultLoop_acc_657_nl;
  wire[21:0] MultLoop_acc_2491_nl;
  wire[23:0] nl_MultLoop_acc_2491_nl;
  wire[11:0] MultLoop_acc_4197_nl;
  wire[12:0] nl_MultLoop_acc_4197_nl;
  wire[20:0] MultLoop_acc_4673_nl;
  wire[21:0] nl_MultLoop_acc_4673_nl;
  wire[24:0] MultLoop_acc_649_nl;
  wire[25:0] nl_MultLoop_acc_649_nl;
  wire[23:0] MultLoop_acc_2495_nl;
  wire[25:0] nl_MultLoop_acc_2495_nl;
  wire[24:0] MultLoop_acc_643_nl;
  wire[26:0] nl_MultLoop_acc_643_nl;
  wire[22:0] MultLoop_acc_1296_nl;
  wire[23:0] nl_MultLoop_acc_1296_nl;
  wire[21:0] MultLoop_acc_2499_nl;
  wire[22:0] nl_MultLoop_acc_2499_nl;
  wire[22:0] MultLoop_acc_1295_nl;
  wire[23:0] nl_MultLoop_acc_1295_nl;
  wire[20:0] MultLoop_acc_2501_nl;
  wire[21:0] nl_MultLoop_acc_2501_nl;
  wire[24:0] MultLoop_acc_637_nl;
  wire[25:0] nl_MultLoop_acc_637_nl;
  wire[22:0] MultLoop_acc_2503_nl;
  wire[24:0] nl_MultLoop_acc_2503_nl;
  wire[21:0] MultLoop_acc_632_nl;
  wire[22:0] nl_MultLoop_acc_632_nl;
  wire[18:0] MultLoop_acc_2505_nl;
  wire[19:0] nl_MultLoop_acc_2505_nl;
  wire[22:0] MultLoop_acc_622_nl;
  wire[23:0] nl_MultLoop_acc_622_nl;
  wire[20:0] MultLoop_acc_2508_nl;
  wire[21:0] nl_MultLoop_acc_2508_nl;
  wire[17:0] MultLoop_acc_2507_nl;
  wire[18:0] nl_MultLoop_acc_2507_nl;
  wire[20:0] MultLoop_acc_1289_nl;
  wire[21:0] nl_MultLoop_acc_1289_nl;
  wire[18:0] MultLoop_acc_2509_nl;
  wire[19:0] nl_MultLoop_acc_2509_nl;
  wire[17:0] MultLoop_acc_4202_nl;
  wire[18:0] nl_MultLoop_acc_4202_nl;
  wire[21:0] MultLoop_acc_2512_nl;
  wire[23:0] nl_MultLoop_acc_2512_nl;
  wire[12:0] MultLoop_acc_4201_nl;
  wire[13:0] nl_MultLoop_acc_4201_nl;
  wire[17:0] MultLoop_acc_4204_nl;
  wire[18:0] nl_MultLoop_acc_4204_nl;
  wire[23:0] MultLoop_acc_2515_nl;
  wire[24:0] nl_MultLoop_acc_2515_nl;
  wire[20:0] MultLoop_acc_2514_nl;
  wire[21:0] nl_MultLoop_acc_2514_nl;
  wire[14:0] MultLoop_625_MultLoop_acc_3_nl;
  wire[15:0] nl_MultLoop_625_MultLoop_acc_3_nl;
  wire[22:0] MultLoop_acc_616_nl;
  wire[23:0] nl_MultLoop_acc_616_nl;
  wire[20:0] MultLoop_acc_2518_nl;
  wire[21:0] nl_MultLoop_acc_2518_nl;
  wire[17:0] MultLoop_acc_4207_nl;
  wire[18:0] nl_MultLoop_acc_4207_nl;
  wire[18:0] MultLoop_acc_4674_nl;
  wire[19:0] nl_MultLoop_acc_4674_nl;
  wire[22:0] MultLoop_acc_1300_nl;
  wire[23:0] nl_MultLoop_acc_1300_nl;
  wire[20:0] MultLoop_acc_2523_nl;
  wire[21:0] nl_MultLoop_acc_2523_nl;
  wire[17:0] MultLoop_acc_4209_nl;
  wire[18:0] nl_MultLoop_acc_4209_nl;
  wire[21:0] MultLoop_acc_2527_nl;
  wire[22:0] nl_MultLoop_acc_2527_nl;
  wire[19:0] MultLoop_acc_2526_nl;
  wire[20:0] nl_MultLoop_acc_2526_nl;
  wire[21:0] MultLoop_acc_1297_nl;
  wire[22:0] nl_MultLoop_acc_1297_nl;
  wire[18:0] MultLoop_acc_2537_nl;
  wire[19:0] nl_MultLoop_acc_2537_nl;
  wire[17:0] MultLoop_acc_641_nl;
  wire[18:0] nl_MultLoop_acc_641_nl;
  wire[23:0] MultLoop_acc_651_nl;
  wire[25:0] nl_MultLoop_acc_651_nl;
  wire[23:0] MultLoop_acc_646_nl;
  wire[25:0] nl_MultLoop_acc_646_nl;
  wire[13:0] MultLoop_acc_4211_nl;
  wire[14:0] nl_MultLoop_acc_4211_nl;
  wire[22:0] MultLoop_acc_647_nl;
  wire[23:0] nl_MultLoop_acc_647_nl;
  wire[20:0] MultLoop_acc_2534_nl;
  wire[21:0] nl_MultLoop_acc_2534_nl;
  wire[17:0] MultLoop_acc_2533_nl;
  wire[18:0] nl_MultLoop_acc_2533_nl;
  wire[22:0] MultLoop_acc_1298_nl;
  wire[23:0] nl_MultLoop_acc_1298_nl;
  wire[21:0] MultLoop_acc_2536_nl;
  wire[22:0] nl_MultLoop_acc_2536_nl;
  wire[17:0] MultLoop_acc_4214_nl;
  wire[18:0] nl_MultLoop_acc_4214_nl;
  wire[23:0] MultLoop_acc_2540_nl;
  wire[25:0] nl_MultLoop_acc_2540_nl;
  wire[17:0] MultLoop_acc_629_nl;
  wire[18:0] nl_MultLoop_acc_629_nl;
  wire[22:0] MultLoop_acc_1290_nl;
  wire[23:0] nl_MultLoop_acc_1290_nl;
  wire[20:0] MultLoop_acc_2542_nl;
  wire[22:0] nl_MultLoop_acc_2542_nl;
  wire[22:0] MultLoop_acc_625_nl;
  wire[23:0] nl_MultLoop_acc_625_nl;
  wire[19:0] MultLoop_acc_2544_nl;
  wire[20:0] nl_MultLoop_acc_2544_nl;
  wire[23:0] MultLoop_acc_4624_nl;
  wire[24:0] nl_MultLoop_acc_4624_nl;
  wire[17:0] MultLoop_acc_631_nl;
  wire[18:0] nl_MultLoop_acc_631_nl;
  wire[19:0] MultLoop_acc_628_nl;
  wire[20:0] nl_MultLoop_acc_628_nl;
  wire[18:0] MultLoop_acc_2478_nl;
  wire[19:0] nl_MultLoop_acc_2478_nl;
  wire[14:0] MultLoop_acc_4216_nl;
  wire[15:0] nl_MultLoop_acc_4216_nl;
  wire[11:0] nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl;
  wire[13:0] nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl;
  wire[17:0] MultLoop_acc_627_nl;
  wire[18:0] nl_MultLoop_acc_627_nl;
  wire[0:0] nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl;
  wire[24:0] MultLoop_acc_1302_nl;
  wire[25:0] nl_MultLoop_acc_1302_nl;
  wire[17:0] MultLoop_acc_2547_nl;
  wire[18:0] nl_MultLoop_acc_2547_nl;
  wire[18:0] MultLoop_acc_4218_nl;
  wire[19:0] nl_MultLoop_acc_4218_nl;
  wire[21:0] MultLoop_acc_1251_nl;
  wire[22:0] nl_MultLoop_acc_1251_nl;
  wire[17:0] MultLoop_acc_2849_nl;
  wire[18:0] nl_MultLoop_acc_2849_nl;
  wire[20:0] MultLoop_acc_482_nl;
  wire[21:0] nl_MultLoop_acc_482_nl;
  wire[18:0] MultLoop_acc_2843_nl;
  wire[19:0] nl_MultLoop_acc_2843_nl;
  wire[15:0] MultLoop_482_MultLoop_acc_3_nl;
  wire[16:0] nl_MultLoop_482_MultLoop_acc_3_nl;
  wire[13:0] MultLoop_acc_2847_nl;
  wire[14:0] nl_MultLoop_acc_2847_nl;
  wire[18:0] MultLoop_acc_1239_nl;
  wire[19:0] nl_MultLoop_acc_1239_nl;
  wire[22:0] MultLoop_acc_477_nl;
  wire[23:0] nl_MultLoop_acc_477_nl;
  wire[21:0] MultLoop_acc_2846_nl;
  wire[23:0] nl_MultLoop_acc_2846_nl;
  wire[25:0] MultLoop_acc_505_nl;
  wire[26:0] nl_MultLoop_acc_505_nl;
  wire[22:0] MultLoop_acc_2852_nl;
  wire[23:0] nl_MultLoop_acc_2852_nl;
  wire[20:0] MultLoop_acc_2851_nl;
  wire[21:0] nl_MultLoop_acc_2851_nl;
  wire[23:0] MultLoop_acc_504_nl;
  wire[25:0] nl_MultLoop_acc_504_nl;
  wire[13:0] MultLoop_acc_4280_nl;
  wire[14:0] nl_MultLoop_acc_4280_nl;
  wire[20:0] MultLoop_acc_1245_nl;
  wire[21:0] nl_MultLoop_acc_1245_nl;
  wire[17:0] MultLoop_acc_2856_nl;
  wire[18:0] nl_MultLoop_acc_2856_nl;
  wire[10:0] MultLoop_acc_4281_nl;
  wire[11:0] nl_MultLoop_acc_4281_nl;
  wire[19:0] MultLoop_acc_483_nl;
  wire[20:0] nl_MultLoop_acc_483_nl;
  wire[18:0] MultLoop_acc_2858_nl;
  wire[19:0] nl_MultLoop_acc_2858_nl;
  wire[14:0] MultLoop_acc_4282_nl;
  wire[15:0] nl_MultLoop_acc_4282_nl;
  wire[21:0] MultLoop_acc_500_nl;
  wire[22:0] nl_MultLoop_acc_500_nl;
  wire[19:0] MultLoop_acc_2787_nl;
  wire[20:0] nl_MultLoop_acc_2787_nl;
  wire[17:0] MultLoop_acc_2786_nl;
  wire[18:0] nl_MultLoop_acc_2786_nl;
  wire[12:0] MultLoop_acc_4285_nl;
  wire[13:0] nl_MultLoop_acc_4285_nl;
  wire[17:0] MultLoop_acc_4287_nl;
  wire[18:0] nl_MultLoop_acc_4287_nl;
  wire[19:0] MultLoop_acc_2789_nl;
  wire[20:0] nl_MultLoop_acc_2789_nl;
  wire[20:0] MultLoop_acc_487_nl;
  wire[21:0] nl_MultLoop_acc_487_nl;
  wire[16:0] MultLoop_acc_4283_nl;
  wire[17:0] nl_MultLoop_acc_4283_nl;
  wire[11:0] MultLoop_acc_2860_nl;
  wire[13:0] nl_MultLoop_acc_2860_nl;
  wire[20:0] MultLoop_acc_495_nl;
  wire[21:0] nl_MultLoop_acc_495_nl;
  wire[16:0] MultLoop_acc_4284_nl;
  wire[17:0] nl_MultLoop_acc_4284_nl;
  wire[23:0] MultLoop_acc_518_nl;
  wire[25:0] nl_MultLoop_acc_518_nl;
  wire[21:0] MultLoop_acc_519_nl;
  wire[22:0] nl_MultLoop_acc_519_nl;
  wire[19:0] MultLoop_acc_2794_nl;
  wire[20:0] nl_MultLoop_acc_2794_nl;
  wire[17:0] MultLoop_acc_2793_nl;
  wire[18:0] nl_MultLoop_acc_2793_nl;
  wire[20:0] MultLoop_acc_1247_nl;
  wire[21:0] nl_MultLoop_acc_1247_nl;
  wire[18:0] MultLoop_acc_2795_nl;
  wire[19:0] nl_MultLoop_acc_2795_nl;
  wire[17:0] MultLoop_acc_4291_nl;
  wire[18:0] nl_MultLoop_acc_4291_nl;
  wire[20:0] MultLoop_acc_2797_nl;
  wire[21:0] nl_MultLoop_acc_2797_nl;
  wire[23:0] MultLoop_acc_501_nl;
  wire[24:0] nl_MultLoop_acc_501_nl;
  wire[21:0] MultLoop_acc_2799_nl;
  wire[22:0] nl_MultLoop_acc_2799_nl;
  wire[21:0] MultLoop_acc_1246_nl;
  wire[22:0] nl_MultLoop_acc_1246_nl;
  wire[17:0] MultLoop_acc_2801_nl;
  wire[18:0] nl_MultLoop_acc_2801_nl;
  wire[17:0] MultLoop_acc_497_nl;
  wire[18:0] nl_MultLoop_acc_497_nl;
  wire[18:0] MultLoop_acc_4631_nl;
  wire[19:0] nl_MultLoop_acc_4631_nl;
  wire[17:0] MultLoop_acc_4294_nl;
  wire[18:0] nl_MultLoop_acc_4294_nl;
  wire[21:0] MultLoop_acc_2805_nl;
  wire[23:0] nl_MultLoop_acc_2805_nl;
  wire[19:0] MultLoop_acc_1240_nl;
  wire[20:0] nl_MultLoop_acc_1240_nl;
  wire[17:0] MultLoop_acc_2806_nl;
  wire[18:0] nl_MultLoop_acc_2806_nl;
  wire[21:0] MultLoop_acc_521_nl;
  wire[22:0] nl_MultLoop_acc_521_nl;
  wire[19:0] MultLoop_acc_2810_nl;
  wire[20:0] nl_MultLoop_acc_2810_nl;
  wire[17:0] MultLoop_acc_2809_nl;
  wire[18:0] nl_MultLoop_acc_2809_nl;
  wire[17:0] MultLoop_acc_4298_nl;
  wire[18:0] nl_MultLoop_acc_4298_nl;
  wire[22:0] MultLoop_acc_2813_nl;
  wire[24:0] nl_MultLoop_acc_2813_nl;
  wire[18:0] MultLoop_acc_4632_nl;
  wire[19:0] nl_MultLoop_acc_4632_nl;
  wire[19:0] MultLoop_acc_4633_nl;
  wire[20:0] nl_MultLoop_acc_4633_nl;
  wire[19:0] MultLoop_acc_494_nl;
  wire[20:0] nl_MultLoop_acc_494_nl;
  wire[18:0] MultLoop_acc_2783_nl;
  wire[19:0] nl_MultLoop_acc_2783_nl;
  wire[14:0] MultLoop_acc_4295_nl;
  wire[15:0] nl_MultLoop_acc_4295_nl;
  wire[17:0] MultLoop_acc_4304_nl;
  wire[18:0] nl_MultLoop_acc_4304_nl;
  wire[18:0] MultLoop_acc_4677_nl;
  wire[19:0] nl_MultLoop_acc_4677_nl;
  wire[22:0] MultLoop_acc_516_nl;
  wire[23:0] nl_MultLoop_acc_516_nl;
  wire[20:0] MultLoop_acc_2816_nl;
  wire[22:0] nl_MultLoop_acc_2816_nl;
  wire[10:0] MultLoop_acc_4299_nl;
  wire[11:0] nl_MultLoop_acc_4299_nl;
  wire[20:0] MultLoop_acc_514_nl;
  wire[21:0] nl_MultLoop_acc_514_nl;
  wire[16:0] MultLoop_acc_4300_nl;
  wire[17:0] nl_MultLoop_acc_4300_nl;
  wire[22:0] MultLoop_acc_515_nl;
  wire[24:0] nl_MultLoop_acc_515_nl;
  wire[14:0] MultLoop_acc_4301_nl;
  wire[15:0] nl_MultLoop_acc_4301_nl;
  wire[23:0] MultLoop_acc_1250_nl;
  wire[24:0] nl_MultLoop_acc_1250_nl;
  wire[20:0] MultLoop_acc_2822_nl;
  wire[21:0] nl_MultLoop_acc_2822_nl;
  wire[17:0] MultLoop_acc_2821_nl;
  wire[18:0] nl_MultLoop_acc_2821_nl;
  wire[11:0] MultLoop_acc_4302_nl;
  wire[12:0] nl_MultLoop_acc_4302_nl;
  wire[17:0] MultLoop_acc_4306_nl;
  wire[18:0] nl_MultLoop_acc_4306_nl;
  wire[19:0] MultLoop_acc_4678_nl;
  wire[20:0] nl_MultLoop_acc_4678_nl;
  wire[18:0] MultLoop_acc_1248_nl;
  wire[19:0] nl_MultLoop_acc_1248_nl;
  wire[18:0] MultLoop_acc_4310_nl;
  wire[19:0] nl_MultLoop_acc_4310_nl;
  wire[24:0] MultLoop_acc_489_nl;
  wire[26:0] nl_MultLoop_acc_489_nl;
  wire[17:0] MultLoop_acc_4308_nl;
  wire[18:0] nl_MultLoop_acc_4308_nl;
  wire[22:0] MultLoop_acc_2833_nl;
  wire[23:0] nl_MultLoop_acc_2833_nl;
  wire[19:0] MultLoop_acc_2832_nl;
  wire[20:0] nl_MultLoop_acc_2832_nl;
  wire[17:0] MultLoop_acc_2831_nl;
  wire[18:0] nl_MultLoop_acc_2831_nl;
  wire[22:0] MultLoop_acc_502_nl;
  wire[23:0] nl_MultLoop_acc_502_nl;
  wire[14:0] MultLoop_acc_4309_nl;
  wire[15:0] nl_MultLoop_acc_4309_nl;
  wire[20:0] MultLoop_acc_1244_nl;
  wire[21:0] nl_MultLoop_acc_1244_nl;
  wire[18:0] MultLoop_acc_2835_nl;
  wire[19:0] nl_MultLoop_acc_2835_nl;
  wire[17:0] MultLoop_acc_491_nl;
  wire[18:0] nl_MultLoop_acc_491_nl;
  wire[23:0] MultLoop_acc_1242_nl;
  wire[24:0] nl_MultLoop_acc_1242_nl;
  wire[19:0] MultLoop_acc_2841_nl;
  wire[21:0] nl_MultLoop_acc_2841_nl;
  wire[23:0] MultLoop_acc_1287_nl;
  wire[24:0] nl_MultLoop_acc_1287_nl;
  wire[17:0] MultLoop_acc_4222_nl;
  wire[18:0] nl_MultLoop_acc_4222_nl;
  wire[22:0] MultLoop_acc_2602_nl;
  wire[24:0] nl_MultLoop_acc_2602_nl;
  wire[13:0] MultLoop_acc_1268_nl;
  wire[14:0] nl_MultLoop_acc_1268_nl;
  wire[22:0] MultLoop_acc_1271_nl;
  wire[23:0] nl_MultLoop_acc_1271_nl;
  wire[19:0] MultLoop_acc_2595_nl;
  wire[20:0] nl_MultLoop_acc_2595_nl;
  wire[17:0] MultLoop_acc_2594_nl;
  wire[18:0] nl_MultLoop_acc_2594_nl;
  wire[20:0] MultLoop_acc_1272_nl;
  wire[21:0] nl_MultLoop_acc_1272_nl;
  wire[17:0] MultLoop_acc_2596_nl;
  wire[18:0] nl_MultLoop_acc_2596_nl;
  wire[21:0] MultLoop_acc_1270_nl;
  wire[22:0] nl_MultLoop_acc_1270_nl;
  wire[17:0] MultLoop_acc_2598_nl;
  wire[18:0] nl_MultLoop_acc_2598_nl;
  wire[25:0] MultLoop_acc_575_nl;
  wire[26:0] nl_MultLoop_acc_575_nl;
  wire[25:0] MultLoop_acc_608_nl;
  wire[27:0] nl_MultLoop_acc_608_nl;
  wire[22:0] MultLoop_acc_1281_nl;
  wire[23:0] nl_MultLoop_acc_1281_nl;
  wire[20:0] MultLoop_acc_2609_nl;
  wire[21:0] nl_MultLoop_acc_2609_nl;
  wire[17:0] MultLoop_acc_2608_nl;
  wire[18:0] nl_MultLoop_acc_2608_nl;
  wire[18:0] MultLoop_acc_4226_nl;
  wire[19:0] nl_MultLoop_acc_4226_nl;
  wire[19:0] MultLoop_acc_2610_nl;
  wire[20:0] nl_MultLoop_acc_2610_nl;
  wire[25:0] MultLoop_acc_593_nl;
  wire[27:0] nl_MultLoop_acc_593_nl;
  wire[11:0] MultLoop_acc_4227_nl;
  wire[12:0] nl_MultLoop_acc_4227_nl;
  wire[22:0] MultLoop_acc_1278_nl;
  wire[23:0] nl_MultLoop_acc_1278_nl;
  wire[17:0] MultLoop_acc_2614_nl;
  wire[18:0] nl_MultLoop_acc_2614_nl;
  wire[21:0] MultLoop_acc_1277_nl;
  wire[22:0] nl_MultLoop_acc_1277_nl;
  wire[17:0] MultLoop_acc_2616_nl;
  wire[18:0] nl_MultLoop_acc_2616_nl;
  wire[22:0] MultLoop_acc_1269_nl;
  wire[23:0] nl_MultLoop_acc_1269_nl;
  wire[19:0] MultLoop_acc_2619_nl;
  wire[21:0] nl_MultLoop_acc_2619_nl;
  wire[19:0] MultLoop_acc_1286_nl;
  wire[20:0] nl_MultLoop_acc_1286_nl;
  wire[17:0] MultLoop_acc_2559_nl;
  wire[18:0] nl_MultLoop_acc_2559_nl;
  wire[19:0] MultLoop_acc_598_nl;
  wire[20:0] nl_MultLoop_acc_598_nl;
  wire[18:0] MultLoop_acc_2561_nl;
  wire[19:0] nl_MultLoop_acc_2561_nl;
  wire[17:0] MultLoop_acc_571_nl;
  wire[18:0] nl_MultLoop_acc_571_nl;
  wire[22:0] MultLoop_acc_615_nl;
  wire[23:0] nl_MultLoop_acc_615_nl;
  wire[14:0] MultLoop_acc_4232_nl;
  wire[15:0] nl_MultLoop_acc_4232_nl;
  wire[22:0] MultLoop_acc_1284_nl;
  wire[23:0] nl_MultLoop_acc_1284_nl;
  wire[17:0] MultLoop_acc_2563_nl;
  wire[18:0] nl_MultLoop_acc_2563_nl;
  wire[20:0] MultLoop_acc_610_nl;
  wire[21:0] nl_MultLoop_acc_610_nl;
  wire[18:0] MultLoop_acc_2565_nl;
  wire[19:0] nl_MultLoop_acc_2565_nl;
  wire[18:0] MultLoop_acc_4625_nl;
  wire[19:0] nl_MultLoop_acc_4625_nl;
  wire[22:0] MultLoop_acc_4626_nl;
  wire[23:0] nl_MultLoop_acc_4626_nl;
  wire[22:0] MultLoop_acc_1282_nl;
  wire[23:0] nl_MultLoop_acc_1282_nl;
  wire[21:0] MultLoop_acc_2569_nl;
  wire[22:0] nl_MultLoop_acc_2569_nl;
  wire[18:0] MultLoop_acc_4627_nl;
  wire[19:0] nl_MultLoop_acc_4627_nl;
  wire[20:0] MultLoop_acc_601_nl;
  wire[21:0] nl_MultLoop_acc_601_nl;
  wire[16:0] MultLoop_acc_4234_nl;
  wire[17:0] nl_MultLoop_acc_4234_nl;
  wire[17:0] MultLoop_acc_4236_nl;
  wire[18:0] nl_MultLoop_acc_4236_nl;
  wire[21:0] MultLoop_acc_2573_nl;
  wire[22:0] nl_MultLoop_acc_2573_nl;
  wire[21:0] MultLoop_acc_1276_nl;
  wire[22:0] nl_MultLoop_acc_1276_nl;
  wire[20:0] MultLoop_acc_2575_nl;
  wire[21:0] nl_MultLoop_acc_2575_nl;
  wire[23:0] MultLoop_acc_580_nl;
  wire[25:0] nl_MultLoop_acc_580_nl;
  wire[13:0] MultLoop_acc_4237_nl;
  wire[14:0] nl_MultLoop_acc_4237_nl;
  wire[21:0] MultLoop_acc_1273_nl;
  wire[22:0] nl_MultLoop_acc_1273_nl;
  wire[17:0] MultLoop_acc_2578_nl;
  wire[18:0] nl_MultLoop_acc_2578_nl;
  wire[20:0] MultLoop_acc_591_nl;
  wire[21:0] nl_MultLoop_acc_591_nl;
  wire[11:0] MultLoop_acc_2620_nl;
  wire[12:0] nl_MultLoop_acc_2620_nl;
  wire[21:0] MultLoop_acc_611_nl;
  wire[22:0] nl_MultLoop_acc_611_nl;
  wire[15:0] MultLoop_acc_4238_nl;
  wire[16:0] nl_MultLoop_acc_4238_nl;
  wire[19:0] MultLoop_acc_585_nl;
  wire[20:0] nl_MultLoop_acc_585_nl;
  wire[24:0] MultLoop_acc_605_nl;
  wire[25:0] nl_MultLoop_acc_605_nl;
  wire[20:0] MultLoop_acc_2579_nl;
  wire[21:0] nl_MultLoop_acc_2579_nl;
  wire[18:0] MultLoop_acc_4239_nl;
  wire[19:0] nl_MultLoop_acc_4239_nl;
  wire[22:0] MultLoop_acc_2581_nl;
  wire[24:0] nl_MultLoop_acc_2581_nl;
  wire[17:0] MultLoop_acc_596_nl;
  wire[18:0] nl_MultLoop_acc_596_nl;
  wire[18:0] MultLoop_acc_4629_nl;
  wire[19:0] nl_MultLoop_acc_4629_nl;
  wire[20:0] MultLoop_acc_4628_nl;
  wire[21:0] nl_MultLoop_acc_4628_nl;
  wire[17:0] MultLoop_acc_4675_nl;
  wire[18:0] nl_MultLoop_acc_4675_nl;
  wire[17:0] MultLoop_acc_4242_nl;
  wire[18:0] nl_MultLoop_acc_4242_nl;
  wire[19:0] MultLoop_acc_2587_nl;
  wire[20:0] nl_MultLoop_acc_2587_nl;
  wire[17:0] MultLoop_acc_2586_nl;
  wire[18:0] nl_MultLoop_acc_2586_nl;
  wire[17:0] MultLoop_acc_4244_nl;
  wire[18:0] nl_MultLoop_acc_4244_nl;
  wire[23:0] MultLoop_acc_2590_nl;
  wire[25:0] nl_MultLoop_acc_2590_nl;
  wire[25:0] MultLoop_acc_581_nl;
  wire[26:0] nl_MultLoop_acc_581_nl;
  wire[24:0] MultLoop_acc_2593_nl;
  wire[25:0] nl_MultLoop_acc_2593_nl;
  wire[20:0] MultLoop_acc_1266_nl;
  wire[21:0] nl_MultLoop_acc_1266_nl;
  wire[18:0] MultLoop_acc_2723_nl;
  wire[19:0] nl_MultLoop_acc_2723_nl;
  wire[20:0] MultLoop_acc_4247_nl;
  wire[21:0] nl_MultLoop_acc_4247_nl;
  wire[17:0] MultLoop_acc_4246_nl;
  wire[18:0] nl_MultLoop_acc_4246_nl;
  wire[19:0] MultLoop_acc_2725_nl;
  wire[20:0] nl_MultLoop_acc_2725_nl;
  wire[20:0] MultLoop_acc_4250_nl;
  wire[21:0] nl_MultLoop_acc_4250_nl;
  wire[17:0] MultLoop_acc_4249_nl;
  wire[18:0] nl_MultLoop_acc_4249_nl;
  wire[21:0] MultLoop_acc_2729_nl;
  wire[23:0] nl_MultLoop_acc_2729_nl;
  wire[10:0] MultLoop_acc_4248_nl;
  wire[11:0] nl_MultLoop_acc_4248_nl;
  wire[23:0] MultLoop_acc_523_nl;
  wire[25:0] nl_MultLoop_acc_523_nl;
  wire[13:0] MultLoop_acc_4251_nl;
  wire[14:0] nl_MultLoop_acc_4251_nl;
  wire[20:0] MultLoop_acc_1267_nl;
  wire[21:0] nl_MultLoop_acc_1267_nl;
  wire[17:0] MultLoop_acc_2667_nl;
  wire[18:0] nl_MultLoop_acc_2667_nl;
  wire[23:0] MultLoop_acc_567_nl;
  wire[24:0] nl_MultLoop_acc_567_nl;
  wire[22:0] MultLoop_acc_559_nl;
  wire[23:0] nl_MultLoop_acc_559_nl;
  wire[19:0] MultLoop_acc_4630_nl;
  wire[20:0] nl_MultLoop_acc_4630_nl;
  wire[17:0] MultLoop_acc_4254_nl;
  wire[18:0] nl_MultLoop_acc_4254_nl;
  wire[22:0] MultLoop_acc_2672_nl;
  wire[23:0] nl_MultLoop_acc_2672_nl;
  wire[19:0] MultLoop_acc_2671_nl;
  wire[20:0] nl_MultLoop_acc_2671_nl;
  wire[23:0] MultLoop_acc_546_nl;
  wire[24:0] nl_MultLoop_acc_546_nl;
  wire[20:0] MultLoop_acc_2673_nl;
  wire[21:0] nl_MultLoop_acc_2673_nl;
  wire[22:0] MultLoop_acc_540_nl;
  wire[23:0] nl_MultLoop_acc_540_nl;
  wire[21:0] MultLoop_acc_538_nl;
  wire[22:0] nl_MultLoop_acc_538_nl;
  wire[15:0] MultLoop_acc_4255_nl;
  wire[16:0] nl_MultLoop_acc_4255_nl;
  wire[17:0] MultLoop_acc_4257_nl;
  wire[18:0] nl_MultLoop_acc_4257_nl;
  wire[21:0] MultLoop_acc_2676_nl;
  wire[22:0] nl_MultLoop_acc_2676_nl;
  wire[18:0] MultLoop_acc_1255_nl;
  wire[19:0] nl_MultLoop_acc_1255_nl;
  wire[17:0] MultLoop_acc_535_nl;
  wire[18:0] nl_MultLoop_acc_535_nl;
  wire[17:0] MultLoop_acc_4259_nl;
  wire[18:0] nl_MultLoop_acc_4259_nl;
  wire[22:0] MultLoop_acc_2679_nl;
  wire[23:0] nl_MultLoop_acc_2679_nl;
  wire[19:0] MultLoop_acc_2678_nl;
  wire[20:0] nl_MultLoop_acc_2678_nl;
  wire[18:0] MultLoop_acc_1261_nl;
  wire[19:0] nl_MultLoop_acc_1261_nl;
  wire[17:0] MultLoop_acc_544_nl;
  wire[18:0] nl_MultLoop_acc_544_nl;
  wire[21:0] MultLoop_acc_1257_nl;
  wire[22:0] nl_MultLoop_acc_1257_nl;
  wire[19:0] MultLoop_acc_2681_nl;
  wire[20:0] nl_MultLoop_acc_2681_nl;
  wire[17:0] MultLoop_acc_4261_nl;
  wire[18:0] nl_MultLoop_acc_4261_nl;
  wire[20:0] MultLoop_acc_2683_nl;
  wire[21:0] nl_MultLoop_acc_2683_nl;
  wire[11:0] MultLoop_acc_4260_nl;
  wire[12:0] nl_MultLoop_acc_4260_nl;
  wire[21:0] MultLoop_acc_1254_nl;
  wire[22:0] nl_MultLoop_acc_1254_nl;
  wire[18:0] MultLoop_acc_2684_nl;
  wire[19:0] nl_MultLoop_acc_2684_nl;
  wire[14:0] MultLoop_acc_2743_nl;
  wire[17:0] nl_MultLoop_acc_2743_nl;
  wire[20:0] MultLoop_acc_1259_nl;
  wire[21:0] nl_MultLoop_acc_1259_nl;
  wire[17:0] MultLoop_acc_2666_nl;
  wire[18:0] nl_MultLoop_acc_2666_nl;
  wire[14:0] MultLoop_acc_4263_nl;
  wire[15:0] nl_MultLoop_acc_4263_nl;
  wire[9:0] MultLoop_acc_2733_nl;
  wire[10:0] nl_MultLoop_acc_2733_nl;
  wire[20:0] MultLoop_acc_1253_nl;
  wire[21:0] nl_MultLoop_acc_1253_nl;
  wire[21:0] MultLoop_acc_530_nl;
  wire[22:0] nl_MultLoop_acc_530_nl;
  wire[19:0] MultLoop_acc_2688_nl;
  wire[20:0] nl_MultLoop_acc_2688_nl;
  wire[17:0] MultLoop_acc_2687_nl;
  wire[18:0] nl_MultLoop_acc_2687_nl;
  wire[24:0] MultLoop_acc_568_nl;
  wire[25:0] nl_MultLoop_acc_568_nl;
  wire[19:0] MultLoop_acc_2689_nl;
  wire[20:0] nl_MultLoop_acc_2689_nl;
  wire[20:0] MultLoop_acc_564_nl;
  wire[21:0] nl_MultLoop_acc_564_nl;
  wire[18:0] MultLoop_acc_2691_nl;
  wire[19:0] nl_MultLoop_acc_2691_nl;
  wire[10:0] MultLoop_acc_4264_nl;
  wire[11:0] nl_MultLoop_acc_4264_nl;
  wire[23:0] MultLoop_acc_562_nl;
  wire[24:0] nl_MultLoop_acc_562_nl;
  wire[20:0] MultLoop_acc_2692_nl;
  wire[21:0] nl_MultLoop_acc_2692_nl;
  wire[23:0] MultLoop_acc_1265_nl;
  wire[24:0] nl_MultLoop_acc_1265_nl;
  wire[19:0] MultLoop_acc_2694_nl;
  wire[20:0] nl_MultLoop_acc_2694_nl;
  wire[22:0] MultLoop_acc_1262_nl;
  wire[23:0] nl_MultLoop_acc_1262_nl;
  wire[17:0] MultLoop_acc_2703_nl;
  wire[18:0] nl_MultLoop_acc_2703_nl;
  wire[25:0] MultLoop_acc_553_nl;
  wire[26:0] nl_MultLoop_acc_553_nl;
  wire[21:0] MultLoop_acc_2705_nl;
  wire[22:0] nl_MultLoop_acc_2705_nl;
  wire[19:0] MultLoop_acc_2704_nl;
  wire[20:0] nl_MultLoop_acc_2704_nl;
  wire[23:0] MultLoop_acc_1264_nl;
  wire[24:0] nl_MultLoop_acc_1264_nl;
  wire[21:0] MultLoop_acc_2696_nl;
  wire[22:0] nl_MultLoop_acc_2696_nl;
  wire[21:0] MultLoop_acc_1263_nl;
  wire[22:0] nl_MultLoop_acc_1263_nl;
  wire[17:0] MultLoop_acc_2697_nl;
  wire[18:0] nl_MultLoop_acc_2697_nl;
  wire[18:0] MultLoop_acc_4265_nl;
  wire[19:0] nl_MultLoop_acc_4265_nl;
  wire[21:0] MultLoop_acc_2698_nl;
  wire[22:0] nl_MultLoop_acc_2698_nl;
  wire[22:0] MultLoop_acc_554_nl;
  wire[23:0] nl_MultLoop_acc_554_nl;
  wire[19:0] MultLoop_acc_2701_nl;
  wire[20:0] nl_MultLoop_acc_2701_nl;
  wire[17:0] MultLoop_acc_2700_nl;
  wire[18:0] nl_MultLoop_acc_2700_nl;
  wire[10:0] MultLoop_acc_4266_nl;
  wire[11:0] nl_MultLoop_acc_4266_nl;
  wire[21:0] MultLoop_acc_1260_nl;
  wire[22:0] nl_MultLoop_acc_1260_nl;
  wire[19:0] MultLoop_acc_2707_nl;
  wire[21:0] nl_MultLoop_acc_2707_nl;
  wire[17:0] MultLoop_acc_4269_nl;
  wire[18:0] nl_MultLoop_acc_4269_nl;
  wire[22:0] MultLoop_acc_2709_nl;
  wire[23:0] nl_MultLoop_acc_2709_nl;
  wire[18:0] MultLoop_acc_4275_nl;
  wire[19:0] nl_MultLoop_acc_4275_nl;
  wire[19:0] MultLoop_acc_2722_nl;
  wire[20:0] nl_MultLoop_acc_2722_nl;
  wire[17:0] MultLoop_acc_526_nl;
  wire[18:0] nl_MultLoop_acc_526_nl;
  wire[17:0] MultLoop_acc_4274_nl;
  wire[18:0] nl_MultLoop_acc_4274_nl;
  wire[18:0] MultLoop_acc_4676_nl;
  wire[19:0] nl_MultLoop_acc_4676_nl;
  wire[23:0] MultLoop_acc_1256_nl;
  wire[24:0] nl_MultLoop_acc_1256_nl;
  wire[21:0] MultLoop_acc_2711_nl;
  wire[23:0] nl_MultLoop_acc_2711_nl;
  wire[17:0] MultLoop_acc_4271_nl;
  wire[18:0] nl_MultLoop_acc_4271_nl;
  wire[19:0] MultLoop_acc_2714_nl;
  wire[20:0] nl_MultLoop_acc_2714_nl;
  wire[17:0] MultLoop_acc_2713_nl;
  wire[18:0] nl_MultLoop_acc_2713_nl;
  wire[22:0] MultLoop_acc_531_nl;
  wire[23:0] nl_MultLoop_acc_531_nl;
  wire[19:0] MultLoop_acc_2717_nl;
  wire[20:0] nl_MultLoop_acc_2717_nl;
  wire[17:0] MultLoop_acc_2716_nl;
  wire[18:0] nl_MultLoop_acc_2716_nl;
  wire[19:0] MultLoop_acc_1252_nl;
  wire[20:0] nl_MultLoop_acc_1252_nl;
  wire[17:0] MultLoop_acc_2718_nl;
  wire[18:0] nl_MultLoop_acc_2718_nl;
  wire[18:0] MultLoop_acc_3683_nl;
  wire[19:0] nl_MultLoop_acc_3683_nl;
  wire[20:0] MultLoop_acc_3532_nl;
  wire[21:0] nl_MultLoop_acc_3532_nl;
  wire[20:0] MultLoop_acc_3281_nl;
  wire[21:0] nl_MultLoop_acc_3281_nl;
  wire[18:0] MultLoop_acc_1943_nl;
  wire[19:0] nl_MultLoop_acc_1943_nl;
  wire[20:0] MultLoop_acc_1811_nl;
  wire[21:0] nl_MultLoop_acc_1811_nl;
  wire[17:0] MultLoop_acc_1810_nl;
  wire[18:0] nl_MultLoop_acc_1810_nl;
  wire[18:0] MultLoop_acc_4587_nl;
  wire[19:0] nl_MultLoop_acc_4587_nl;
  wire[11:0] MultLoop_acc_4103_nl;
  wire[12:0] nl_MultLoop_acc_4103_nl;
  wire[19:0] MultLoop_acc_3190_nl;
  wire[20:0] nl_MultLoop_acc_3190_nl;
  wire[17:0] MultLoop_acc_3189_nl;
  wire[18:0] nl_MultLoop_acc_3189_nl;
  wire[20:0] MultLoop_acc_3338_nl;
  wire[21:0] nl_MultLoop_acc_3338_nl;
  wire[19:0] MultLoop_acc_1753_nl;
  wire[20:0] nl_MultLoop_acc_1753_nl;
  wire[17:0] MultLoop_acc_25_nl;
  wire[18:0] nl_MultLoop_acc_25_nl;
  wire[19:0] MultLoop_acc_3761_nl;
  wire[20:0] nl_MultLoop_acc_3761_nl;
  wire[17:0] MultLoop_acc_67_nl;
  wire[18:0] nl_MultLoop_acc_67_nl;
  wire[18:0] MultLoop_acc_4588_nl;
  wire[19:0] nl_MultLoop_acc_4588_nl;
  wire[20:0] MultLoop_acc_2317_nl;
  wire[21:0] nl_MultLoop_acc_2317_nl;
  wire[18:0] MultLoop_acc_1097_nl;
  wire[19:0] nl_MultLoop_acc_1097_nl;
  wire[19:0] MultLoop_acc_87_nl;
  wire[20:0] nl_MultLoop_acc_87_nl;
  wire[18:0] MultLoop_acc_1478_nl;
  wire[19:0] nl_MultLoop_acc_1478_nl;
  wire[17:0] MultLoop_acc_3181_nl;
  wire[18:0] nl_MultLoop_acc_3181_nl;
  wire[18:0] MultLoop_acc_1095_nl;
  wire[19:0] nl_MultLoop_acc_1095_nl;
  wire[17:0] MultLoop_acc_3918_nl;
  wire[18:0] nl_MultLoop_acc_3918_nl;
  wire[21:0] MultLoop_acc_1484_nl;
  wire[22:0] nl_MultLoop_acc_1484_nl;
  wire[10:0] MultLoop_acc_3917_nl;
  wire[11:0] nl_MultLoop_acc_3917_nl;
  wire[20:0] MultLoop_acc_447_nl;
  wire[21:0] nl_MultLoop_acc_447_nl;
  wire[23:0] MultLoop_acc_119_nl;
  wire[24:0] nl_MultLoop_acc_119_nl;
  wire[21:0] MultLoop_acc_1482_nl;
  wire[22:0] nl_MultLoop_acc_1482_nl;
  wire[19:0] MultLoop_acc_1481_nl;
  wire[20:0] nl_MultLoop_acc_1481_nl;
  wire[17:0] MultLoop_acc_123_nl;
  wire[18:0] nl_MultLoop_acc_123_nl;
  wire[19:0] MultLoop_acc_4589_nl;
  wire[20:0] nl_MultLoop_acc_4589_nl;
  wire[19:0] MultLoop_acc_3556_nl;
  wire[21:0] nl_MultLoop_acc_3556_nl;
  wire[22:0] MultLoop_acc_1145_nl;
  wire[23:0] nl_MultLoop_acc_1145_nl;
  wire[20:0] MultLoop_acc_1547_nl;
  wire[21:0] nl_MultLoop_acc_1547_nl;
  wire[17:0] MultLoop_acc_1546_nl;
  wire[18:0] nl_MultLoop_acc_1546_nl;
  wire[20:0] MultLoop_acc_2409_nl;
  wire[21:0] nl_MultLoop_acc_2409_nl;
  wire[21:0] MultLoop_acc_1128_nl;
  wire[22:0] nl_MultLoop_acc_1128_nl;
  wire[20:0] MultLoop_acc_1490_nl;
  wire[21:0] nl_MultLoop_acc_1490_nl;
  wire[17:0] MultLoop_acc_1489_nl;
  wire[18:0] nl_MultLoop_acc_1489_nl;
  wire[12:0] MultLoop_acc_4181_nl;
  wire[13:0] nl_MultLoop_acc_4181_nl;
  wire[22:0] MultLoop_acc_181_nl;
  wire[23:0] nl_MultLoop_acc_181_nl;
  wire[20:0] MultLoop_acc_1492_nl;
  wire[21:0] nl_MultLoop_acc_1492_nl;
  wire[13:0] MultLoop_acc_3921_nl;
  wire[14:0] nl_MultLoop_acc_3921_nl;
  wire[17:0] MultLoop_acc_3920_nl;
  wire[18:0] nl_MultLoop_acc_3920_nl;
  wire[20:0] MultLoop_acc_1488_nl;
  wire[21:0] nl_MultLoop_acc_1488_nl;
  wire[12:0] MultLoop_acc_3919_nl;
  wire[13:0] nl_MultLoop_acc_3919_nl;
  wire[21:0] MultLoop_acc_2026_nl;
  wire[23:0] nl_MultLoop_acc_2026_nl;
  wire[23:0] MultLoop_acc_149_nl;
  wire[24:0] nl_MultLoop_acc_149_nl;
  wire[22:0] MultLoop_acc_1486_nl;
  wire[23:0] nl_MultLoop_acc_1486_nl;
  wire[21:0] MultLoop_acc_3213_nl;
  wire[22:0] nl_MultLoop_acc_3213_nl;
  wire[20:0] MultLoop_acc_2252_nl;
  wire[21:0] nl_MultLoop_acc_2252_nl;
  wire[21:0] MultLoop_acc_1154_nl;
  wire[22:0] nl_MultLoop_acc_1154_nl;
  wire[19:0] MultLoop_acc_1494_nl;
  wire[21:0] nl_MultLoop_acc_1494_nl;
  wire[18:0] MultLoop_acc_2040_nl;
  wire[19:0] nl_MultLoop_acc_2040_nl;
  wire[22:0] MultLoop_acc_434_nl;
  wire[23:0] nl_MultLoop_acc_434_nl;
  wire[21:0] MultLoop_acc_2935_nl;
  wire[22:0] nl_MultLoop_acc_2935_nl;
  wire[18:0] MultLoop_acc_2807_nl;
  wire[19:0] nl_MultLoop_acc_2807_nl;
  wire[21:0] MultLoop_acc_1543_nl;
  wire[22:0] nl_MultLoop_acc_1543_nl;
  wire[18:0] MultLoop_acc_1152_nl;
  wire[19:0] nl_MultLoop_acc_1152_nl;
  wire[21:0] MultLoop_acc_1848_nl;
  wire[23:0] nl_MultLoop_acc_1848_nl;
  wire[18:0] MultLoop_acc_1541_nl;
  wire[19:0] nl_MultLoop_acc_1541_nl;
  wire[19:0] MultLoop_acc_3062_nl;
  wire[20:0] nl_MultLoop_acc_3062_nl;
  wire[20:0] MultLoop_acc_1715_nl;
  wire[21:0] nl_MultLoop_acc_1715_nl;
  wire[18:0] MultLoop_acc_1476_nl;
  wire[19:0] nl_MultLoop_acc_1476_nl;
  wire[21:0] MultLoop_acc_307_nl;
  wire[22:0] nl_MultLoop_acc_307_nl;
  wire[15:0] MultLoop_acc_3922_nl;
  wire[16:0] nl_MultLoop_acc_3922_nl;
  wire[20:0] MultLoop_acc_334_nl;
  wire[21:0] nl_MultLoop_acc_334_nl;
  wire[18:0] MultLoop_acc_1499_nl;
  wire[19:0] nl_MultLoop_acc_1499_nl;
  wire[13:0] MultLoop_acc_3924_nl;
  wire[14:0] nl_MultLoop_acc_3924_nl;
  wire[20:0] MultLoop_acc_2145_nl;
  wire[21:0] nl_MultLoop_acc_2145_nl;
  wire[21:0] MultLoop_acc_335_nl;
  wire[22:0] nl_MultLoop_acc_335_nl;
  wire[15:0] MultLoop_acc_4391_nl;
  wire[16:0] nl_MultLoop_acc_4391_nl;
  wire[18:0] MultLoop_acc_4594_nl;
  wire[19:0] nl_MultLoop_acc_4594_nl;
  wire[19:0] MultLoop_acc_2836_nl;
  wire[20:0] nl_MultLoop_acc_2836_nl;
  wire[19:0] MultLoop_acc_343_nl;
  wire[20:0] nl_MultLoop_acc_343_nl;
  wire[17:0] MultLoop_acc_340_nl;
  wire[18:0] nl_MultLoop_acc_340_nl;
  wire[20:0] MultLoop_acc_2289_nl;
  wire[21:0] nl_MultLoop_acc_2289_nl;
  wire[20:0] MultLoop_acc_355_nl;
  wire[21:0] nl_MultLoop_acc_355_nl;
  wire[19:0] MultLoop_acc_1204_nl;
  wire[20:0] nl_MultLoop_acc_1204_nl;
  wire[17:0] MultLoop_acc_1501_nl;
  wire[18:0] nl_MultLoop_acc_1501_nl;
  wire[19:0] MultLoop_acc_1200_nl;
  wire[20:0] nl_MultLoop_acc_1200_nl;
  wire[17:0] MultLoop_acc_1500_nl;
  wire[18:0] nl_MultLoop_acc_1500_nl;
  wire[19:0] MultLoop_acc_2802_nl;
  wire[20:0] nl_MultLoop_acc_2802_nl;
  wire[20:0] MultLoop_acc_410_nl;
  wire[21:0] nl_MultLoop_acc_410_nl;
  wire[23:0] MultLoop_acc_408_nl;
  wire[24:0] nl_MultLoop_acc_408_nl;
  wire[22:0] MultLoop_acc_1507_nl;
  wire[23:0] nl_MultLoop_acc_1507_nl;
  wire[19:0] MultLoop_acc_2906_nl;
  wire[20:0] nl_MultLoop_acc_2906_nl;
  wire[22:0] MultLoop_acc_400_nl;
  wire[24:0] nl_MultLoop_acc_400_nl;
  wire[14:0] MultLoop_acc_3926_nl;
  wire[15:0] nl_MultLoop_acc_3926_nl;
  wire[21:0] MultLoop_acc_1227_nl;
  wire[22:0] nl_MultLoop_acc_1227_nl;
  wire[17:0] MultLoop_acc_1509_nl;
  wire[18:0] nl_MultLoop_acc_1509_nl;
  wire[13:0] MultLoop_acc_3927_nl;
  wire[14:0] nl_MultLoop_acc_3927_nl;
  wire[10:0] Result_acc_202_nl;
  wire[11:0] nl_Result_acc_202_nl;
  wire[20:0] MultLoop_acc_4590_nl;
  wire[21:0] nl_MultLoop_acc_4590_nl;
  wire[21:0] MultLoop_acc_471_nl;
  wire[22:0] nl_MultLoop_acc_471_nl;
  wire[20:0] MultLoop_acc_1237_nl;
  wire[21:0] nl_MultLoop_acc_1237_nl;
  wire[17:0] MultLoop_acc_1511_nl;
  wire[18:0] nl_MultLoop_acc_1511_nl;
  wire[11:0] MultLoop_acc_3928_nl;
  wire[12:0] nl_MultLoop_acc_3928_nl;
  wire[10:0] MultLoop_acc_4157_nl;
  wire[11:0] nl_MultLoop_acc_4157_nl;
  wire[20:0] MultLoop_acc_2669_nl;
  wire[21:0] nl_MultLoop_acc_2669_nl;
  wire[20:0] MultLoop_acc_1866_nl;
  wire[21:0] nl_MultLoop_acc_1866_nl;
  wire[11:0] MultLoop_acc_3986_nl;
  wire[12:0] nl_MultLoop_acc_3986_nl;
  wire[17:0] MultLoop_acc_3930_nl;
  wire[18:0] nl_MultLoop_acc_3930_nl;
  wire[24:0] MultLoop_acc_1516_nl;
  wire[25:0] nl_MultLoop_acc_1516_nl;
  wire[21:0] MultLoop_acc_1515_nl;
  wire[22:0] nl_MultLoop_acc_1515_nl;
  wire[17:0] MultLoop_acc_506_nl;
  wire[18:0] nl_MultLoop_acc_506_nl;
  wire[19:0] MultLoop_acc_2340_nl;
  wire[20:0] nl_MultLoop_acc_2340_nl;
  wire[24:0] MultLoop_acc_528_nl;
  wire[26:0] nl_MultLoop_acc_528_nl;
  wire[23:0] MultLoop_acc_541_nl;
  wire[24:0] nl_MultLoop_acc_541_nl;
  wire[22:0] MultLoop_acc_1521_nl;
  wire[23:0] nl_MultLoop_acc_1521_nl;
  wire[20:0] MultLoop_acc_1275_nl;
  wire[21:0] nl_MultLoop_acc_1275_nl;
  wire[17:0] MultLoop_acc_1528_nl;
  wire[18:0] nl_MultLoop_acc_1528_nl;
  wire[14:0] MultLoop_acc_3934_nl;
  wire[15:0] nl_MultLoop_acc_3934_nl;
  wire[19:0] MultLoop_acc_579_nl;
  wire[20:0] nl_MultLoop_acc_579_nl;
  wire[18:0] MultLoop_acc_1526_nl;
  wire[19:0] nl_MultLoop_acc_1526_nl;
  wire[13:0] MultLoop_acc_3933_nl;
  wire[14:0] nl_MultLoop_acc_3933_nl;
  wire[21:0] MultLoop_acc_570_nl;
  wire[22:0] nl_MultLoop_acc_570_nl;
  wire[19:0] MultLoop_acc_1524_nl;
  wire[20:0] nl_MultLoop_acc_1524_nl;
  wire[17:0] MultLoop_acc_1523_nl;
  wire[18:0] nl_MultLoop_acc_1523_nl;
  wire[10:0] MultLoop_acc_3932_nl;
  wire[11:0] nl_MultLoop_acc_3932_nl;
  wire[11:0] MultLoop_acc_3935_nl;
  wire[12:0] nl_MultLoop_acc_3935_nl;
  wire[22:0] MultLoop_acc_1730_nl;
  wire[23:0] nl_MultLoop_acc_1730_nl;
  wire[20:0] MultLoop_acc_1816_nl;
  wire[21:0] nl_MultLoop_acc_1816_nl;
  wire[23:0] MultLoop_acc_713_nl;
  wire[24:0] nl_MultLoop_acc_713_nl;
  wire[20:0] MultLoop_acc_1532_nl;
  wire[21:0] nl_MultLoop_acc_1532_nl;
  wire[17:0] MultLoop_acc_785_nl;
  wire[18:0] nl_MultLoop_acc_785_nl;
  wire[19:0] MultLoop_acc_4663_nl;
  wire[20:0] nl_MultLoop_acc_4663_nl;
  wire[25:0] MultLoop_acc_826_nl;
  wire[27:0] nl_MultLoop_acc_826_nl;
  wire[11:0] MultLoop_acc_3937_nl;
  wire[12:0] nl_MultLoop_acc_3937_nl;
  wire[18:0] MultLoop_acc_1479_nl;
  wire[19:0] nl_MultLoop_acc_1479_nl;
  wire[18:0] MultLoop_acc_4592_nl;
  wire[19:0] nl_MultLoop_acc_4592_nl;
  wire[18:0] MultLoop_acc_4593_nl;
  wire[19:0] nl_MultLoop_acc_4593_nl;
  wire[22:0] MultLoop_acc_1350_nl;
  wire[23:0] nl_MultLoop_acc_1350_nl;
  wire[17:0] MultLoop_acc_1540_nl;
  wire[18:0] nl_MultLoop_acc_1540_nl;
  wire[21:0] MultLoop_acc_807_nl;
  wire[22:0] nl_MultLoop_acc_807_nl;
  wire[19:0] MultLoop_acc_1537_nl;
  wire[21:0] nl_MultLoop_acc_1537_nl;
  wire[20:0] MultLoop_acc_1512_nl;
  wire[21:0] nl_MultLoop_acc_1512_nl;
  wire[20:0] Result_acc_102_nl;
  wire[21:0] nl_Result_acc_102_nl;
  wire[18:0] MultLoop_acc_1993_nl;
  wire[19:0] nl_MultLoop_acc_1993_nl;
  wire[22:0] MultLoop_acc_856_nl;
  wire[23:0] nl_MultLoop_acc_856_nl;
  wire[14:0] MultLoop_acc_3938_nl;
  wire[15:0] nl_MultLoop_acc_3938_nl;
  wire[19:0] Result_acc_154_nl;
  wire[20:0] nl_Result_acc_154_nl;
  wire[18:0] MultLoop_acc_4591_nl;
  wire[19:0] nl_MultLoop_acc_4591_nl;
  wire[17:0] MultLoop_acc_150_nl;
  wire[18:0] nl_MultLoop_acc_150_nl;
  wire[21:0] MultLoop_acc_1191_nl;
  wire[22:0] nl_MultLoop_acc_1191_nl;
  wire[17:0] MultLoop_acc_1497_nl;
  wire[18:0] nl_MultLoop_acc_1497_nl;
  wire[23:0] MultLoop_acc_1211_nl;
  wire[24:0] nl_MultLoop_acc_1211_nl;
  wire[20:0] MultLoop_acc_1504_nl;
  wire[21:0] nl_MultLoop_acc_1504_nl;
  wire[19:0] MultLoop_acc_1243_nl;
  wire[20:0] nl_MultLoop_acc_1243_nl;
  wire[17:0] MultLoop_acc_1513_nl;
  wire[18:0] nl_MultLoop_acc_1513_nl;
  wire[19:0] MultLoop_acc_1315_nl;
  wire[20:0] nl_MultLoop_acc_1315_nl;
  wire[17:0] MultLoop_acc_1529_nl;
  wire[18:0] nl_MultLoop_acc_1529_nl;
  wire[22:0] MultLoop_acc_1324_nl;
  wire[23:0] nl_MultLoop_acc_1324_nl;
  wire[20:0] MultLoop_acc_1535_nl;
  wire[21:0] nl_MultLoop_acc_1535_nl;
  wire[17:0] MultLoop_acc_1534_nl;
  wire[18:0] nl_MultLoop_acc_1534_nl;
  wire[12:0] MultLoop_acc_3936_nl;
  wire[13:0] nl_MultLoop_acc_3936_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [431:0] nl_res_rsci_d;
  assign nl_res_rsci_d = {res_rsci_d_431_414 , res_rsci_d_413_396 , res_rsci_d_395_378
      , res_rsci_d_377_360 , res_rsci_d_359_342 , res_rsci_d_341_324 , res_rsci_d_323_306
      , res_rsci_d_305_288 , res_rsci_d_287_270 , res_rsci_d_269_252 , res_rsci_d_251_234
      , res_rsci_d_233_216 , res_rsci_d_215_198 , res_rsci_d_197_180 , res_rsci_d_179_162
      , res_rsci_d_161_144 , res_rsci_d_143_126 , res_rsci_d_125_108 , res_rsci_d_107_90
      , res_rsci_d_89_72 , res_rsci_d_71_54 , res_rsci_d_53_36 , res_rsci_d_35_18
      , res_rsci_d_17_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd864)) data_rsci (
      .dat(data_rsc_dat),
      .idat(data_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd2),
  .width(32'sd432)) res_rsci (
      .d(nl_res_rsci_d[431:0]),
      .z(res_rsc_z)
    );
  assign nl_MultLoop_acc_3683_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_16_19(data_rsci_idat[17:2]);
  assign MultLoop_acc_3683_nl = nl_MultLoop_acc_3683_nl[18:0];
  assign MultLoop_acc_3683_itm_18_3_1 = readslicef_19_16_3((MultLoop_acc_3683_nl));
  assign nl_MultLoop_acc_3532_nl = ({(data_rsci_idat[647:630]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_2568_cse_1);
  assign MultLoop_acc_3532_nl = nl_MultLoop_acc_3532_nl[20:0];
  assign MultLoop_acc_3532_itm_20_5_1 = readslicef_21_16_5((MultLoop_acc_3532_nl));
  assign nl_MultLoop_acc_3283_cse = conv_s2s_18_19(data_rsci_idat[503:486]) + conv_s2s_16_19(data_rsci_idat[503:488]);
  assign MultLoop_acc_3283_cse = nl_MultLoop_acc_3283_cse[18:0];
  assign nl_MultLoop_acc_3105_cse = conv_s2s_18_19(data_rsci_idat[485:468]) + conv_s2s_16_19(data_rsci_idat[485:470]);
  assign MultLoop_acc_3105_cse = nl_MultLoop_acc_3105_cse[18:0];
  assign nl_MultLoop_acc_2133_cse_1 = (~ (data_rsci_idat[521:504])) + conv_s2s_16_18(data_rsci_idat[521:506]);
  assign MultLoop_acc_2133_cse_1 = nl_MultLoop_acc_2133_cse_1[17:0];
  assign nl_MultLoop_acc_2535_cse_1 = (~ (data_rsci_idat[485:468])) + conv_s2s_16_18(data_rsci_idat[485:470]);
  assign MultLoop_acc_2535_cse_1 = nl_MultLoop_acc_2535_cse_1[17:0];
  assign nl_MultLoop_acc_4229_cse_1 = conv_s2u_10_11(data_rsci_idat[377:368]) + 11'b00000000001;
  assign MultLoop_acc_4229_cse_1 = nl_MultLoop_acc_4229_cse_1[10:0];
  assign nl_MultLoop_acc_2591_cse_1 = conv_s2s_18_19(data_rsci_idat[251:234]) + conv_s2s_16_19(data_rsci_idat[251:236]);
  assign MultLoop_acc_2591_cse_1 = nl_MultLoop_acc_2591_cse_1[18:0];
  assign nl_MultLoop_acc_3099_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[215:198]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[215:198]));
  assign MultLoop_acc_3099_cse_1 = nl_MultLoop_acc_3099_cse_1[21:0];
  assign nl_MultLoop_acc_1946_cse_1 = (~ (data_rsci_idat[791:774])) + conv_s2s_15_18(data_rsci_idat[791:777]);
  assign MultLoop_acc_1946_cse_1 = nl_MultLoop_acc_1946_cse_1[17:0];
  assign nl_MultLoop_acc_3961_cse_1 = conv_s2u_12_13(data_rsci_idat[863:852]) + 13'b0000000000001;
  assign MultLoop_acc_3961_cse_1 = nl_MultLoop_acc_3961_cse_1[12:0];
  assign nl_Result_acc_192_cse_1 = conv_s2u_12_13(data_rsci_idat[773:762]) + 13'b0000000000001;
  assign Result_acc_192_cse_1 = nl_Result_acc_192_cse_1[12:0];
  assign nl_MultLoop_acc_3281_nl = ({(data_rsci_idat[647:630]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[647:630]));
  assign MultLoop_acc_3281_nl = nl_MultLoop_acc_3281_nl[20:0];
  assign MultLoop_acc_3281_itm_20_6 = readslicef_21_15_6((MultLoop_acc_3281_nl));
  assign nl_MultLoop_acc_1943_nl = conv_s2s_18_19(data_rsci_idat[629:612]) + conv_s2s_14_19(data_rsci_idat[629:616]);
  assign MultLoop_acc_1943_nl = nl_MultLoop_acc_1943_nl[18:0];
  assign MultLoop_acc_1943_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1943_nl));
  assign nl_MultLoop_acc_3661_cse_1 = conv_s2s_18_19(data_rsci_idat[323:306]) + conv_s2s_15_19(data_rsci_idat[323:309]);
  assign MultLoop_acc_3661_cse_1 = nl_MultLoop_acc_3661_cse_1[18:0];
  assign nl_MultLoop_acc_2387_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[593:576]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[593:576]));
  assign MultLoop_acc_2387_cse_1 = nl_MultLoop_acc_2387_cse_1[20:0];
  assign nl_MultLoop_acc_1810_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_16_18(data_rsci_idat[557:542]);
  assign MultLoop_acc_1810_nl = nl_MultLoop_acc_1810_nl[17:0];
  assign nl_MultLoop_acc_1811_nl = conv_s2s_20_21({(~ (data_rsci_idat[557:540]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1810_nl);
  assign MultLoop_acc_1811_nl = nl_MultLoop_acc_1811_nl[20:0];
  assign MultLoop_acc_1811_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1811_nl));
  assign nl_MultLoop_acc_4587_nl = conv_s2u_17_19(MultLoop_acc_1476_itm_18_2) + conv_s2u_18_19(data_rsci_idat[431:414]);
  assign MultLoop_acc_4587_nl = nl_MultLoop_acc_4587_nl[18:0];
  assign MultLoop_acc_4587_itm_18_3 = readslicef_19_16_3((MultLoop_acc_4587_nl));
  assign nl_MultLoop_acc_4103_nl = conv_s2s_11_12(data_rsci_idat[719:709]) + 12'b000000000001;
  assign MultLoop_acc_4103_nl = nl_MultLoop_acc_4103_nl[11:0];
  assign nl_MultLoop_acc_2220_cse_1 = conv_s2s_18_19(data_rsci_idat[719:702]) + conv_s2s_17_19({(MultLoop_acc_4103_nl)
      , (data_rsci_idat[708:704])});
  assign MultLoop_acc_2220_cse_1 = nl_MultLoop_acc_2220_cse_1[18:0];
  assign nl_MultLoop_acc_3189_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_16_18(data_rsci_idat[395:380]);
  assign MultLoop_acc_3189_nl = nl_MultLoop_acc_3189_nl[17:0];
  assign nl_MultLoop_acc_3190_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3189_nl);
  assign MultLoop_acc_3190_nl = nl_MultLoop_acc_3190_nl[19:0];
  assign MultLoop_acc_3190_itm_19_4 = readslicef_20_16_4((MultLoop_acc_3190_nl));
  assign nl_MultLoop_acc_3338_nl = conv_s2s_20_21({(~ (data_rsci_idat[35:18])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_3338_nl = nl_MultLoop_acc_3338_nl[20:0];
  assign MultLoop_acc_3338_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_3338_nl));
  assign nl_MultLoop_acc_1753_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[53:36]));
  assign MultLoop_acc_1753_nl = nl_MultLoop_acc_1753_nl[19:0];
  assign MultLoop_acc_1753_itm_19_4 = readslicef_20_16_4((MultLoop_acc_1753_nl));
  assign nl_MultLoop_acc_1722_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[17:0]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[17:0]));
  assign MultLoop_acc_1722_cse_1 = nl_MultLoop_acc_1722_cse_1[20:0];
  assign nl_MultLoop_acc_25_nl = conv_s2u_14_18(data_rsci_idat[413:400]) - (data_rsci_idat[413:396]);
  assign MultLoop_acc_25_nl = nl_MultLoop_acc_25_nl[17:0];
  assign MultLoop_acc_25_itm_17_5 = readslicef_18_13_5((MultLoop_acc_25_nl));
  assign nl_MultLoop_acc_3761_nl = ({(data_rsci_idat[107:90]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[107:90]));
  assign MultLoop_acc_3761_nl = nl_MultLoop_acc_3761_nl[19:0];
  assign MultLoop_acc_3761_itm_19_6 = readslicef_20_14_6((MultLoop_acc_3761_nl));
  assign nl_MultLoop_acc_67_nl = conv_s2u_13_18(data_rsci_idat[341:329]) - (data_rsci_idat[341:324]);
  assign MultLoop_acc_67_nl = nl_MultLoop_acc_67_nl[17:0];
  assign MultLoop_acc_67_itm_17_3 = readslicef_18_15_3((MultLoop_acc_67_nl));
  assign nl_MultLoop_acc_4588_nl = conv_s2u_16_19(MultLoop_acc_1479_itm_18_3) + conv_s2u_18_19(data_rsci_idat[809:792]);
  assign MultLoop_acc_4588_nl = nl_MultLoop_acc_4588_nl[18:0];
  assign MultLoop_acc_4588_itm_18_2 = readslicef_19_17_2((MultLoop_acc_4588_nl));
  assign nl_MultLoop_acc_4212_cse_1 = conv_s2u_10_11(data_rsci_idat[575:566]) + 11'b00000000001;
  assign MultLoop_acc_4212_cse_1 = nl_MultLoop_acc_4212_cse_1[10:0];
  assign nl_MultLoop_acc_1611_cse_1 = conv_s2s_18_19(data_rsci_idat[269:252]) + conv_s2s_16_19(data_rsci_idat[269:254]);
  assign MultLoop_acc_1611_cse_1 = nl_MultLoop_acc_1611_cse_1[18:0];
  assign nl_MultLoop_acc_4167_cse_1 = conv_s2u_10_11(data_rsci_idat[539:530]) + 11'b00000000001;
  assign MultLoop_acc_4167_cse_1 = nl_MultLoop_acc_4167_cse_1[10:0];
  assign nl_MultLoop_acc_2317_nl = ({(data_rsci_idat[503:486]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[503:486]));
  assign MultLoop_acc_2317_nl = nl_MultLoop_acc_2317_nl[20:0];
  assign MultLoop_acc_2317_itm_20_5 = readslicef_21_16_5((MultLoop_acc_2317_nl));
  assign nl_MultLoop_acc_2584_cse_1 = conv_s2s_18_19(data_rsci_idat[431:414]) + conv_s2s_17_19({MultLoop_MultLoop_conc_794_16_5
      , (data_rsci_idat[420:416])});
  assign MultLoop_acc_2584_cse_1 = nl_MultLoop_acc_2584_cse_1[18:0];
  assign nl_MultLoop_acc_3636_cse_1 = ({(data_rsci_idat[863:846]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[863:846]));
  assign MultLoop_acc_3636_cse_1 = nl_MultLoop_acc_3636_cse_1[19:0];
  assign nl_MultLoop_acc_1097_nl = conv_s2u_14_19(data_rsci_idat[593:580]) + conv_s2u_18_19(data_rsci_idat[593:576]);
  assign MultLoop_acc_1097_nl = nl_MultLoop_acc_1097_nl[18:0];
  assign MultLoop_acc_1097_itm_18_4 = readslicef_19_15_4((MultLoop_acc_1097_nl));
  assign nl_MultLoop_acc_2057_cse_1 = conv_s2s_18_19(data_rsci_idat[287:270]) + conv_s2s_16_19(data_rsci_idat[287:272]);
  assign MultLoop_acc_2057_cse_1 = nl_MultLoop_acc_2057_cse_1[18:0];
  assign nl_MultLoop_acc_1478_nl = conv_s2s_18_19(data_rsci_idat[719:702]) + conv_s2s_15_19({MultLoop_acc_3916_cse_1
      , (data_rsci_idat[707:706])});
  assign MultLoop_acc_1478_nl = nl_MultLoop_acc_1478_nl[18:0];
  assign nl_MultLoop_acc_87_nl = conv_s2u_19_20(MultLoop_acc_1478_nl) + ({(~ (data_rsci_idat[719:702]))
      , 2'b00});
  assign MultLoop_acc_87_nl = nl_MultLoop_acc_87_nl[19:0];
  assign MultLoop_acc_87_itm_19_4 = readslicef_20_16_4((MultLoop_acc_87_nl));
  assign nl_MultLoop_acc_3181_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_16_18(data_rsci_idat[611:596]);
  assign MultLoop_acc_3181_nl = nl_MultLoop_acc_3181_nl[17:0];
  assign nl_MultLoop_acc_3182_cse_1 = ({(data_rsci_idat[611:594]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3181_nl);
  assign MultLoop_acc_3182_cse_1 = nl_MultLoop_acc_3182_cse_1[19:0];
  assign nl_MultLoop_acc_2307_cse_1 = (~ (data_rsci_idat[773:756])) + conv_s2s_16_18(data_rsci_idat[773:758]);
  assign MultLoop_acc_2307_cse_1 = nl_MultLoop_acc_2307_cse_1[17:0];
  assign nl_MultLoop_acc_2685_cse_1 = (~ (data_rsci_idat[125:108])) + conv_s2s_16_18(data_rsci_idat[125:110]);
  assign MultLoop_acc_2685_cse_1 = nl_MultLoop_acc_2685_cse_1[17:0];
  assign nl_MultLoop_acc_1095_nl = conv_s2u_13_19(data_rsci_idat[521:509]) + conv_s2u_18_19(data_rsci_idat[521:504]);
  assign MultLoop_acc_1095_nl = nl_MultLoop_acc_1095_nl[18:0];
  assign MultLoop_acc_1095_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1095_nl));
  assign nl_MultLoop_acc_3917_nl =  -conv_s2s_10_11(data_rsci_idat[467:458]);
  assign MultLoop_acc_3917_nl = nl_MultLoop_acc_3917_nl[10:0];
  assign nl_MultLoop_acc_1484_nl = ({(data_rsci_idat[467:450]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_3917_nl)
      , (~ (data_rsci_idat[457:450]))});
  assign MultLoop_acc_1484_nl = nl_MultLoop_acc_1484_nl[21:0];
  assign nl_MultLoop_acc_3918_nl = conv_s2u_14_18(readslicef_22_14_8((MultLoop_acc_1484_nl)))
      + (~ (data_rsci_idat[467:450]));
  assign MultLoop_acc_3918_nl = nl_MultLoop_acc_3918_nl[17:0];
  assign MultLoop_acc_3918_itm_17_2 = readslicef_18_16_2((MultLoop_acc_3918_nl));
  assign nl_MultLoop_acc_447_nl = conv_s2s_18_21(~ (data_rsci_idat[341:324])) + ({(data_rsci_idat[341:324])
      , 3'b001});
  assign MultLoop_acc_447_nl = nl_MultLoop_acc_447_nl[20:0];
  assign MultLoop_acc_447_itm_20_7 = readslicef_21_14_7((MultLoop_acc_447_nl));
  assign nl_MultLoop_acc_1949_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[737:720]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_820_18_8 , (~ (data_rsci_idat[727:720]))});
  assign MultLoop_acc_1949_cse_1 = nl_MultLoop_acc_1949_cse_1[20:0];
  assign nl_Result_acc_214_cse_1 = conv_s2u_10_11(data_rsci_idat[755:746]) + 11'b00000000001;
  assign Result_acc_214_cse_1 = nl_Result_acc_214_cse_1[10:0];
  assign nl_MultLoop_acc_1481_nl = ({(data_rsci_idat[431:414]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[431:414]));
  assign MultLoop_acc_1481_nl = nl_MultLoop_acc_1481_nl[19:0];
  assign nl_MultLoop_acc_1482_nl = ({(~ (data_rsci_idat[431:414])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_1481_nl);
  assign MultLoop_acc_1482_nl = nl_MultLoop_acc_1482_nl[21:0];
  assign nl_MultLoop_acc_119_nl = conv_s2s_22_24(MultLoop_acc_1482_nl) + ({(data_rsci_idat[431:414])
      , 6'b010000});
  assign MultLoop_acc_119_nl = nl_MultLoop_acc_119_nl[23:0];
  assign MultLoop_acc_119_itm_23_9 = readslicef_24_15_9((MultLoop_acc_119_nl));
  assign nl_MultLoop_acc_4083_cse_1 = conv_s2u_11_12(data_rsci_idat[791:781]) + 12'b000000000001;
  assign MultLoop_acc_4083_cse_1 = nl_MultLoop_acc_4083_cse_1[11:0];
  assign nl_MultLoop_acc_123_nl = conv_s2u_16_18(data_rsci_idat[503:488]) - (data_rsci_idat[503:486]);
  assign MultLoop_acc_123_nl = nl_MultLoop_acc_123_nl[17:0];
  assign MultLoop_acc_123_itm_17_3 = readslicef_18_15_3((MultLoop_acc_123_nl));
  assign nl_MultLoop_acc_3946_cse_1 = conv_s2u_12_13(data_rsci_idat[413:402]) + 13'b0000000000001;
  assign MultLoop_acc_3946_cse_1 = nl_MultLoop_acc_3946_cse_1[12:0];
  assign nl_MultLoop_acc_4589_nl = conv_s2u_19_20(MultLoop_acc_1480_cse_1[20:2])
      + ({(data_rsci_idat[305:288]) , 2'b01});
  assign MultLoop_acc_4589_nl = nl_MultLoop_acc_4589_nl[19:0];
  assign MultLoop_acc_4589_itm_19_4 = readslicef_20_16_4((MultLoop_acc_4589_nl));
  assign nl_MultLoop_acc_3556_nl = ({(~ (data_rsci_idat[35:18])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[35:18])
      + conv_s2s_16_20(data_rsci_idat[35:20]);
  assign MultLoop_acc_3556_nl = nl_MultLoop_acc_3556_nl[19:0];
  assign MultLoop_acc_3556_itm_19_2_1 = readslicef_20_18_2((MultLoop_acc_3556_nl));
  assign nl_Result_acc_178_cse_1 = conv_s2u_10_11(data_rsci_idat[827:818]) + 11'b00000000001;
  assign Result_acc_178_cse_1 = nl_Result_acc_178_cse_1[10:0];
  assign nl_MultLoop_acc_4233_cse_1 = conv_s2u_11_12(data_rsci_idat[773:763]) + 12'b000000000001;
  assign MultLoop_acc_4233_cse_1 = nl_MultLoop_acc_4233_cse_1[11:0];
  assign nl_MultLoop_acc_1546_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18({MultLoop_MultLoop_conc_798_16_4
      , (data_rsci_idat[167:164])});
  assign MultLoop_acc_1546_nl = nl_MultLoop_acc_1546_nl[17:0];
  assign nl_MultLoop_acc_1547_nl = conv_s2s_20_21({(~ (data_rsci_idat[179:162]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1546_nl);
  assign MultLoop_acc_1547_nl = nl_MultLoop_acc_1547_nl[20:0];
  assign nl_MultLoop_acc_1145_nl = conv_s2u_21_23(MultLoop_acc_1547_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[179:162])) , 4'b0100});
  assign MultLoop_acc_1145_nl = nl_MultLoop_acc_1145_nl[22:0];
  assign MultLoop_acc_1145_itm_22_7 = readslicef_23_16_7((MultLoop_acc_1145_nl));
  assign nl_MultLoop_acc_1618_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[107:90]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_822_18_7 , (~ (data_rsci_idat[96:90]))});
  assign MultLoop_acc_1618_cse_1 = nl_MultLoop_acc_1618_cse_1[20:0];
  assign nl_MultLoop_acc_2424_cse_1 = conv_s2s_18_19(data_rsci_idat[539:522]) + conv_s2s_16_19({MultLoop_acc_4167_cse_1
      , (data_rsci_idat[529:525])});
  assign MultLoop_acc_2424_cse_1 = nl_MultLoop_acc_2424_cse_1[18:0];
  assign nl_MultLoop_acc_2079_cse_1 = (~ (data_rsci_idat[125:108])) + conv_s2s_14_18(data_rsci_idat[125:112]);
  assign MultLoop_acc_2079_cse_1 = nl_MultLoop_acc_2079_cse_1[17:0];
  assign nl_MultLoop_acc_2568_cse_1 = (~ (data_rsci_idat[647:630])) + conv_s2s_16_18(data_rsci_idat[647:632]);
  assign MultLoop_acc_2568_cse_1 = nl_MultLoop_acc_2568_cse_1[17:0];
  assign nl_MultLoop_acc_2520_cse_1 = ({(data_rsci_idat[773:756]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_846_18_8
      , (~ (data_rsci_idat[763:756]))});
  assign MultLoop_acc_2520_cse_1 = nl_MultLoop_acc_2520_cse_1[19:0];
  assign nl_MultLoop_acc_1720_cse_1 = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[143:126]));
  assign MultLoop_acc_1720_cse_1 = nl_MultLoop_acc_1720_cse_1[20:0];
  assign nl_MultLoop_acc_2409_nl = conv_s2s_20_21({(~ (data_rsci_idat[377:360]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_2409_nl = nl_MultLoop_acc_2409_nl[20:0];
  assign MultLoop_acc_2409_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_2409_nl));
  assign nl_MultLoop_acc_1489_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_16_18(data_rsci_idat[359:344]);
  assign MultLoop_acc_1489_nl = nl_MultLoop_acc_1489_nl[17:0];
  assign nl_MultLoop_acc_1490_nl = conv_s2s_20_21({(~ (data_rsci_idat[359:342]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1489_nl);
  assign MultLoop_acc_1490_nl = nl_MultLoop_acc_1490_nl[20:0];
  assign nl_MultLoop_acc_1128_nl = conv_s2u_21_22(MultLoop_acc_1490_nl) + ({(data_rsci_idat[359:342])
      , 4'b0100});
  assign MultLoop_acc_1128_nl = nl_MultLoop_acc_1128_nl[21:0];
  assign MultLoop_acc_1128_itm_21_7 = readslicef_22_15_7((MultLoop_acc_1128_nl));
  assign nl_MultLoop_acc_4181_nl = conv_s2s_12_13(data_rsci_idat[845:834]) + 13'b0000000000001;
  assign MultLoop_acc_4181_nl = nl_MultLoop_acc_4181_nl[12:0];
  assign nl_MultLoop_acc_2375_cse_1 = (~ (data_rsci_idat[845:828])) + conv_s2s_17_18({(MultLoop_acc_4181_nl)
      , (data_rsci_idat[833:830])});
  assign MultLoop_acc_2375_cse_1 = nl_MultLoop_acc_2375_cse_1[17:0];
  assign nl_MultLoop_acc_3921_nl =  -conv_s2s_13_14(data_rsci_idat[665:653]);
  assign MultLoop_acc_3921_nl = nl_MultLoop_acc_3921_nl[13:0];
  assign nl_MultLoop_acc_1492_nl = ({(data_rsci_idat[665:648]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_3921_nl)
      , (~ (data_rsci_idat[652:648]))});
  assign MultLoop_acc_1492_nl = nl_MultLoop_acc_1492_nl[20:0];
  assign nl_MultLoop_acc_181_nl = conv_s2s_21_23(MultLoop_acc_1492_nl) + ({(~ (data_rsci_idat[665:648]))
      , 5'b00000});
  assign MultLoop_acc_181_nl = nl_MultLoop_acc_181_nl[22:0];
  assign MultLoop_acc_181_itm_22_8 = readslicef_23_15_8((MultLoop_acc_181_nl));
  assign nl_MultLoop_acc_3919_nl =  -conv_s2s_12_13(data_rsci_idat[215:204]);
  assign MultLoop_acc_3919_nl = nl_MultLoop_acc_3919_nl[12:0];
  assign nl_MultLoop_acc_1488_nl = ({(data_rsci_idat[215:198]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_3919_nl)
      , (~ (data_rsci_idat[203:198]))});
  assign MultLoop_acc_1488_nl = nl_MultLoop_acc_1488_nl[20:0];
  assign nl_MultLoop_acc_3920_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_1488_nl)))
      + (~ (data_rsci_idat[215:198]));
  assign MultLoop_acc_3920_nl = nl_MultLoop_acc_3920_nl[17:0];
  assign MultLoop_acc_3920_itm_17_2 = readslicef_18_16_2((MultLoop_acc_3920_nl));
  assign nl_MultLoop_acc_3063_cse_1 = (~ (data_rsci_idat[269:252])) + conv_s2s_15_18(data_rsci_idat[269:255]);
  assign MultLoop_acc_3063_cse_1 = nl_MultLoop_acc_3063_cse_1[17:0];
  assign nl_MultLoop_acc_2026_nl = ({(data_rsci_idat[233:216]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[233:216])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_2026_nl = nl_MultLoop_acc_2026_nl[21:0];
  assign MultLoop_acc_2026_itm_21_6 = readslicef_22_16_6((MultLoop_acc_2026_nl));
  assign nl_MultLoop_acc_1486_nl = conv_s2s_22_23({(~ (data_rsci_idat[89:72])) ,
      4'b0100}) + conv_s2s_21_23(MultLoop_acc_1485_cse_1);
  assign MultLoop_acc_1486_nl = nl_MultLoop_acc_1486_nl[22:0];
  assign nl_MultLoop_acc_149_nl = conv_s2s_23_24(MultLoop_acc_1486_nl) + ({(data_rsci_idat[89:72])
      , 6'b010000});
  assign MultLoop_acc_149_nl = nl_MultLoop_acc_149_nl[23:0];
  assign MultLoop_acc_149_itm_23_8 = readslicef_24_16_8((MultLoop_acc_149_nl));
  assign nl_MultLoop_acc_3187_cse_1 = conv_s2s_18_19(data_rsci_idat[467:450]) + conv_s2s_16_19(data_rsci_idat[467:452]);
  assign MultLoop_acc_3187_cse_1 = nl_MultLoop_acc_3187_cse_1[18:0];
  assign nl_MultLoop_acc_3974_cse_1 = conv_s2u_10_11(data_rsci_idat[233:224]) + 11'b00000000001;
  assign MultLoop_acc_3974_cse_1 = nl_MultLoop_acc_3974_cse_1[10:0];
  assign nl_MultLoop_acc_3213_nl = conv_s2s_21_22({(~ (data_rsci_idat[251:234]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[251:234]));
  assign MultLoop_acc_3213_nl = nl_MultLoop_acc_3213_nl[21:0];
  assign MultLoop_acc_3213_itm_21_3_1 = readslicef_22_19_3((MultLoop_acc_3213_nl));
  assign nl_MultLoop_acc_2390_cse_1 = ({(data_rsci_idat[575:558]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[575:558]));
  assign MultLoop_acc_2390_cse_1 = nl_MultLoop_acc_2390_cse_1[20:0];
  assign nl_MultLoop_acc_2252_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[125:108]));
  assign MultLoop_acc_2252_nl = nl_MultLoop_acc_2252_nl[20:0];
  assign MultLoop_acc_2252_itm_20_5 = readslicef_21_16_5((MultLoop_acc_2252_nl));
  assign nl_MultLoop_acc_1494_nl = ({(~ (data_rsci_idat[611:594])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[611:594])
      + conv_s2s_15_20(data_rsci_idat[611:597]);
  assign MultLoop_acc_1494_nl = nl_MultLoop_acc_1494_nl[19:0];
  assign nl_MultLoop_acc_1154_nl = conv_s2u_20_22(MultLoop_acc_1494_nl) + ({(data_rsci_idat[611:594])
      , 4'b0100});
  assign MultLoop_acc_1154_nl = nl_MultLoop_acc_1154_nl[21:0];
  assign MultLoop_acc_1154_itm_21_6 = readslicef_22_16_6((MultLoop_acc_1154_nl));
  assign nl_Result_acc_190_cse_1 = conv_s2u_12_13(data_rsci_idat[503:492]) + 13'b0000000000001;
  assign Result_acc_190_cse_1 = nl_Result_acc_190_cse_1[12:0];
  assign nl_MultLoop_acc_2040_nl = conv_s2s_18_19(data_rsci_idat[755:738]) + conv_s2s_15_19(data_rsci_idat[755:741]);
  assign MultLoop_acc_2040_nl = nl_MultLoop_acc_2040_nl[18:0];
  assign MultLoop_acc_2040_itm_18_3 = readslicef_19_16_3((MultLoop_acc_2040_nl));
  assign nl_MultLoop_acc_1822_cse_1 = conv_s2s_18_19(data_rsci_idat[863:846]) + conv_s2s_17_19({MultLoop_acc_3961_cse_1
      , (data_rsci_idat[851:848])});
  assign MultLoop_acc_1822_cse_1 = nl_MultLoop_acc_1822_cse_1[18:0];
  assign nl_MultLoop_acc_4122_cse_1 = conv_s2u_10_11(data_rsci_idat[341:332]) + 11'b00000000001;
  assign MultLoop_acc_4122_cse_1 = nl_MultLoop_acc_4122_cse_1[10:0];
  assign nl_MultLoop_acc_2935_nl = conv_s2s_21_22({(~ (data_rsci_idat[107:90])) ,
      3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_2935_nl = nl_MultLoop_acc_2935_nl[21:0];
  assign nl_MultLoop_acc_434_nl = conv_s2s_22_23(MultLoop_acc_2935_nl) + ({(data_rsci_idat[107:90])
      , 5'b01000});
  assign MultLoop_acc_434_nl = nl_MultLoop_acc_434_nl[22:0];
  assign MultLoop_acc_434_itm_22_7 = readslicef_23_16_7((MultLoop_acc_434_nl));
  assign nl_MultLoop_acc_2807_nl = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_14_19(data_rsci_idat[71:58]);
  assign MultLoop_acc_2807_nl = nl_MultLoop_acc_2807_nl[18:0];
  assign MultLoop_acc_2807_itm_18_2 = readslicef_19_17_2((MultLoop_acc_2807_nl));
  assign nl_MultLoop_acc_1543_nl = ({(data_rsci_idat[719:702]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[719:702]));
  assign MultLoop_acc_1543_nl = nl_MultLoop_acc_1543_nl[21:0];
  assign MultLoop_acc_1543_itm_21_6 = readslicef_22_16_6((MultLoop_acc_1543_nl));
  assign nl_MultLoop_acc_1152_nl = conv_s2u_15_19(data_rsci_idat[557:543]) + conv_s2u_18_19(data_rsci_idat[557:540]);
  assign MultLoop_acc_1152_nl = nl_MultLoop_acc_1152_nl[18:0];
  assign MultLoop_acc_1152_itm_18_3 = readslicef_19_16_3((MultLoop_acc_1152_nl));
  assign nl_MultLoop_acc_3941_cse_1 = conv_s2u_11_12(data_rsci_idat[251:241]) + 12'b000000000001;
  assign MultLoop_acc_3941_cse_1 = nl_MultLoop_acc_3941_cse_1[11:0];
  assign nl_MultLoop_acc_4011_cse_1 = conv_s2u_10_11(data_rsci_idat[863:854]) + 11'b00000000001;
  assign MultLoop_acc_4011_cse_1 = nl_MultLoop_acc_4011_cse_1[10:0];
  assign nl_MultLoop_acc_2385_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[683:666]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[683:666]));
  assign MultLoop_acc_2385_cse_1 = nl_MultLoop_acc_2385_cse_1[20:0];
  assign nl_Result_acc_143_cse_1 = (~ (data_rsci_idat[845:828])) + conv_s2s_16_18(data_rsci_idat[845:830]);
  assign Result_acc_143_cse_1 = nl_Result_acc_143_cse_1[17:0];
  assign nl_MultLoop_acc_2566_cse_1 = conv_s2s_18_19(data_rsci_idat[719:702]) + conv_s2s_16_19(data_rsci_idat[719:704]);
  assign MultLoop_acc_2566_cse_1 = nl_MultLoop_acc_2566_cse_1[18:0];
  assign nl_MultLoop_acc_1743_cse_1 = ({(data_rsci_idat[665:648]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[665:648]));
  assign MultLoop_acc_1743_cse_1 = nl_MultLoop_acc_1743_cse_1[20:0];
  assign nl_MultLoop_acc_1848_nl = ({(data_rsci_idat[125:108]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_1848_nl = nl_MultLoop_acc_1848_nl[21:0];
  assign MultLoop_acc_1848_itm_21_6 = readslicef_22_16_6((MultLoop_acc_1848_nl));
  assign nl_Result_acc_111_cse_1 = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_16_19(data_rsci_idat[107:92]);
  assign Result_acc_111_cse_1 = nl_Result_acc_111_cse_1[18:0];
  assign nl_MultLoop_acc_2574_cse_1 = (~ (data_rsci_idat[341:324])) + conv_s2s_16_18(data_rsci_idat[341:326]);
  assign MultLoop_acc_2574_cse_1 = nl_MultLoop_acc_2574_cse_1[17:0];
  assign nl_MultLoop_acc_1541_nl = conv_s2s_18_19(data_rsci_idat[701:684]) + conv_s2s_16_19(data_rsci_idat[701:686]);
  assign MultLoop_acc_1541_nl = nl_MultLoop_acc_1541_nl[18:0];
  assign MultLoop_acc_1541_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1541_nl));
  assign nl_MultLoop_acc_1480_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[305:288]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_1480_cse_1 = nl_MultLoop_acc_1480_cse_1[20:0];
  assign nl_MultLoop_acc_3062_nl = ({(data_rsci_idat[341:324]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2574_cse_1);
  assign MultLoop_acc_3062_nl = nl_MultLoop_acc_3062_nl[19:0];
  assign MultLoop_acc_3062_itm_19_4 = readslicef_20_16_4((MultLoop_acc_3062_nl));
  assign nl_Result_acc_152_cse_1 = (~ (data_rsci_idat[593:576])) + conv_s2s_15_18(data_rsci_idat[593:579]);
  assign Result_acc_152_cse_1 = nl_Result_acc_152_cse_1[17:0];
  assign nl_MultLoop_acc_2073_cse_1 = conv_s2s_18_19(data_rsci_idat[665:648]) + conv_s2s_16_19(data_rsci_idat[665:650]);
  assign MultLoop_acc_2073_cse_1 = nl_MultLoop_acc_2073_cse_1[18:0];
  assign nl_MultLoop_acc_1715_nl = conv_s2s_20_21({(~ (data_rsci_idat[485:468]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[485:468]));
  assign MultLoop_acc_1715_nl = nl_MultLoop_acc_1715_nl[20:0];
  assign MultLoop_acc_1715_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1715_nl));
  assign nl_MultLoop_acc_1476_nl = conv_s2s_18_19(data_rsci_idat[431:414]) + conv_s2s_15_19(data_rsci_idat[431:417]);
  assign MultLoop_acc_1476_nl = nl_MultLoop_acc_1476_nl[18:0];
  assign MultLoop_acc_1476_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1476_nl));
  assign nl_MultLoop_acc_3922_nl =  -conv_s2s_15_16(data_rsci_idat[359:345]);
  assign MultLoop_acc_3922_nl = nl_MultLoop_acc_3922_nl[15:0];
  assign nl_MultLoop_acc_307_nl = conv_s2s_19_22({(MultLoop_acc_3922_nl) , (~ (data_rsci_idat[344:342]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[359:342])) , 3'b001});
  assign MultLoop_acc_307_nl = nl_MultLoop_acc_307_nl[21:0];
  assign MultLoop_acc_307_itm_21_7 = readslicef_22_15_7((MultLoop_acc_307_nl));
  assign nl_MultLoop_acc_2522_cse_1 = conv_s2s_18_19(data_rsci_idat[737:720]) + conv_s2s_16_19(data_rsci_idat[737:722]);
  assign MultLoop_acc_2522_cse_1 = nl_MultLoop_acc_2522_cse_1[18:0];
  assign nl_MultLoop_acc_2967_cse_1 = conv_s2s_18_19(data_rsci_idat[521:504]) + conv_s2s_16_19(data_rsci_idat[521:506]);
  assign MultLoop_acc_2967_cse_1 = nl_MultLoop_acc_2967_cse_1[18:0];
  assign nl_MultLoop_acc_2412_cse_1 = conv_s2s_18_19(data_rsci_idat[125:108]) + conv_s2s_16_19(data_rsci_idat[125:110]);
  assign MultLoop_acc_2412_cse_1 = nl_MultLoop_acc_2412_cse_1[18:0];
  assign nl_MultLoop_acc_1485_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[89:72]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_1485_cse_1 = nl_MultLoop_acc_1485_cse_1[20:0];
  assign nl_MultLoop_acc_3924_nl = conv_s2s_13_14(data_rsci_idat[863:851]) + 14'b00000000000001;
  assign MultLoop_acc_3924_nl = nl_MultLoop_acc_3924_nl[13:0];
  assign nl_MultLoop_acc_1499_nl = conv_s2s_18_19(data_rsci_idat[863:846]) + conv_s2s_17_19({(MultLoop_acc_3924_nl)
      , (data_rsci_idat[850:848])});
  assign MultLoop_acc_1499_nl = nl_MultLoop_acc_1499_nl[18:0];
  assign nl_MultLoop_acc_334_nl = conv_s2u_19_21(MultLoop_acc_1499_nl) + ({(~ (data_rsci_idat[863:846]))
      , 3'b000});
  assign MultLoop_acc_334_nl = nl_MultLoop_acc_334_nl[20:0];
  assign MultLoop_acc_334_itm_20_5 = readslicef_21_16_5((MultLoop_acc_334_nl));
  assign nl_MultLoop_acc_788_cse_1 = conv_s2s_18_20(~ (data_rsci_idat[557:540]))
      + ({(data_rsci_idat[557:540]) , 2'b01});
  assign MultLoop_acc_788_cse_1 = nl_MultLoop_acc_788_cse_1[19:0];
  assign nl_MultLoop_acc_2923_cse_1 = ({(data_rsci_idat[503:486]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[503:486]));
  assign MultLoop_acc_2923_cse_1 = nl_MultLoop_acc_2923_cse_1[19:0];
  assign nl_MultLoop_acc_2145_nl = ({(data_rsci_idat[233:216]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[233:216]));
  assign MultLoop_acc_2145_nl = nl_MultLoop_acc_2145_nl[20:0];
  assign MultLoop_acc_2145_itm_20_5 = readslicef_21_16_5((MultLoop_acc_2145_nl));
  assign nl_MultLoop_acc_4162_cse_1 = conv_s2u_11_12(data_rsci_idat[161:151]) + 12'b000000000001;
  assign MultLoop_acc_4162_cse_1 = nl_MultLoop_acc_4162_cse_1[11:0];
  assign nl_MultLoop_acc_4391_nl =  -conv_s2s_15_16(data_rsci_idat[17:3]);
  assign MultLoop_acc_4391_nl = nl_MultLoop_acc_4391_nl[15:0];
  assign nl_MultLoop_acc_335_nl = conv_s2s_19_22({(MultLoop_acc_4391_nl) , (~ (data_rsci_idat[2:0]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[17:0])) , 3'b001});
  assign MultLoop_acc_335_nl = nl_MultLoop_acc_335_nl[21:0];
  assign MultLoop_acc_335_itm_21_9 = readslicef_22_13_9((MultLoop_acc_335_nl));
  assign nl_MultLoop_acc_4594_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_16_19(MultLoop_acc_1753_itm_19_4);
  assign MultLoop_acc_4594_nl = nl_MultLoop_acc_4594_nl[18:0];
  assign MultLoop_acc_4594_itm_18_2 = readslicef_19_17_2((MultLoop_acc_4594_nl));
  assign nl_MultLoop_acc_1636_cse_1 = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({MultLoop_acc_3955_cse_1
      , (data_rsci_idat[60:56])});
  assign MultLoop_acc_1636_cse_1 = nl_MultLoop_acc_1636_cse_1[17:0];
  assign nl_MultLoop_acc_2836_nl = ({(data_rsci_idat[287:270]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[287:270]));
  assign MultLoop_acc_2836_nl = nl_MultLoop_acc_2836_nl[19:0];
  assign MultLoop_acc_2836_itm_19_6 = readslicef_20_14_6((MultLoop_acc_2836_nl));
  assign nl_MultLoop_acc_4146_cse_1 = conv_s2u_10_11(data_rsci_idat[557:548]) + 11'b00000000001;
  assign MultLoop_acc_4146_cse_1 = nl_MultLoop_acc_4146_cse_1[10:0];
  assign nl_MultLoop_acc_1962_cse_1 = conv_s2s_18_19(data_rsci_idat[539:522]) + conv_s2s_15_19(data_rsci_idat[539:525]);
  assign MultLoop_acc_1962_cse_1 = nl_MultLoop_acc_1962_cse_1[18:0];
  assign nl_Result_acc_206_cse_1 = conv_s2u_10_11(data_rsci_idat[719:710]) + 11'b00000000001;
  assign Result_acc_206_cse_1 = nl_Result_acc_206_cse_1[10:0];
  assign nl_MultLoop_acc_343_nl = conv_s2s_18_20(~ (data_rsci_idat[143:126])) + ({(data_rsci_idat[143:126])
      , 2'b01});
  assign MultLoop_acc_343_nl = nl_MultLoop_acc_343_nl[19:0];
  assign MultLoop_acc_343_itm_19_5 = readslicef_20_15_5((MultLoop_acc_343_nl));
  assign nl_MultLoop_acc_340_nl = conv_s2u_16_18(data_rsci_idat[89:74]) - (data_rsci_idat[89:72]);
  assign MultLoop_acc_340_nl = nl_MultLoop_acc_340_nl[17:0];
  assign MultLoop_acc_340_itm_17_3 = readslicef_18_15_3((MultLoop_acc_340_nl));
  assign nl_MultLoop_acc_2289_nl = ({(data_rsci_idat[809:792]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[809:792]));
  assign MultLoop_acc_2289_nl = nl_MultLoop_acc_2289_nl[20:0];
  assign MultLoop_acc_2289_itm_20_5 = readslicef_21_16_5((MultLoop_acc_2289_nl));
  assign nl_MultLoop_acc_355_nl = conv_s2s_18_21(~ (data_rsci_idat[359:342])) + ({(data_rsci_idat[359:342])
      , 3'b001});
  assign MultLoop_acc_355_nl = nl_MultLoop_acc_355_nl[20:0];
  assign MultLoop_acc_355_itm_20_6 = readslicef_21_15_6((MultLoop_acc_355_nl));
  assign nl_MultLoop_acc_1708_cse_1 = conv_s2s_18_19(data_rsci_idat[629:612]) + conv_s2s_16_19(data_rsci_idat[629:614]);
  assign MultLoop_acc_1708_cse_1 = nl_MultLoop_acc_1708_cse_1[18:0];
  assign nl_MultLoop_acc_1501_nl = (~ (data_rsci_idat[593:576])) + conv_s2s_14_18(data_rsci_idat[593:580]);
  assign MultLoop_acc_1501_nl = nl_MultLoop_acc_1501_nl[17:0];
  assign nl_MultLoop_acc_1204_nl = conv_s2u_18_20(MultLoop_acc_1501_nl) + ({(data_rsci_idat[593:576])
      , 2'b01});
  assign MultLoop_acc_1204_nl = nl_MultLoop_acc_1204_nl[19:0];
  assign MultLoop_acc_1204_itm_19_5 = readslicef_20_15_5((MultLoop_acc_1204_nl));
  assign nl_MultLoop_acc_1500_nl = (~ (data_rsci_idat[467:450])) + conv_s2s_16_18(data_rsci_idat[467:452]);
  assign MultLoop_acc_1500_nl = nl_MultLoop_acc_1500_nl[17:0];
  assign nl_MultLoop_acc_1200_nl = conv_s2u_18_20(MultLoop_acc_1500_nl) + ({(data_rsci_idat[467:450])
      , 2'b01});
  assign MultLoop_acc_1200_nl = nl_MultLoop_acc_1200_nl[19:0];
  assign MultLoop_acc_1200_itm_19_4 = readslicef_20_16_4((MultLoop_acc_1200_nl));
  assign nl_MultLoop_acc_2802_nl = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[251:234]));
  assign MultLoop_acc_2802_nl = nl_MultLoop_acc_2802_nl[19:0];
  assign MultLoop_acc_2802_itm_19_4 = readslicef_20_16_4((MultLoop_acc_2802_nl));
  assign nl_MultLoop_acc_410_nl = conv_s2s_18_21(~ (data_rsci_idat[539:522])) + ({(data_rsci_idat[539:522])
      , 3'b001});
  assign MultLoop_acc_410_nl = nl_MultLoop_acc_410_nl[20:0];
  assign MultLoop_acc_410_itm_20_7 = readslicef_21_14_7((MultLoop_acc_410_nl));
  assign nl_MultLoop_acc_2604_cse_1 = (~ (data_rsci_idat[845:828])) + conv_s2s_17_18({Result_acc_216_cse_1
      , (data_rsci_idat[834:830])});
  assign MultLoop_acc_2604_cse_1 = nl_MultLoop_acc_2604_cse_1[17:0];
  assign nl_MultLoop_acc_4032_cse_1 = conv_s2u_13_14(data_rsci_idat[413:401]) + 14'b00000000000001;
  assign MultLoop_acc_4032_cse_1 = nl_MultLoop_acc_4032_cse_1[13:0];
  assign nl_MultLoop_acc_2592_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[233:216]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_2592_cse_1 = nl_MultLoop_acc_2592_cse_1[21:0];
  assign nl_MultLoop_acc_1507_nl = conv_s2s_22_23({(~ (data_rsci_idat[503:486]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[503:486]));
  assign MultLoop_acc_1507_nl = nl_MultLoop_acc_1507_nl[22:0];
  assign nl_MultLoop_acc_408_nl = conv_s2s_23_24(MultLoop_acc_1507_nl) + ({(data_rsci_idat[503:486])
      , 6'b010000});
  assign MultLoop_acc_408_nl = nl_MultLoop_acc_408_nl[23:0];
  assign MultLoop_acc_408_itm_23_9 = readslicef_24_15_9((MultLoop_acc_408_nl));
  assign nl_MultLoop_acc_2906_nl = ({(data_rsci_idat[755:738]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_842_18_6
      , (~ (data_rsci_idat[743:738]))});
  assign MultLoop_acc_2906_nl = nl_MultLoop_acc_2906_nl[19:0];
  assign MultLoop_acc_2906_itm_19_4 = readslicef_20_16_4((MultLoop_acc_2906_nl));
  assign nl_MultLoop_acc_3926_nl =  -conv_s2s_14_15(data_rsci_idat[359:346]);
  assign MultLoop_acc_3926_nl = nl_MultLoop_acc_3926_nl[14:0];
  assign nl_MultLoop_acc_400_nl = conv_s2s_22_23({(~ (data_rsci_idat[359:342])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[359:342])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_3926_nl)
      , (~ (data_rsci_idat[345:342]))});
  assign MultLoop_acc_400_nl = nl_MultLoop_acc_400_nl[22:0];
  assign MultLoop_acc_400_itm_22_7 = readslicef_23_16_7((MultLoop_acc_400_nl));
  assign nl_MultLoop_acc_3927_nl = conv_s2s_13_14(data_rsci_idat[809:797]) + 14'b00000000000001;
  assign MultLoop_acc_3927_nl = nl_MultLoop_acc_3927_nl[13:0];
  assign nl_MultLoop_acc_1509_nl = (~ (data_rsci_idat[809:792])) + conv_s2s_17_18({(MultLoop_acc_3927_nl)
      , (data_rsci_idat[796:794])});
  assign MultLoop_acc_1509_nl = nl_MultLoop_acc_1509_nl[17:0];
  assign nl_MultLoop_acc_1227_nl = conv_s2u_18_22(MultLoop_acc_1509_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[809:792])) , 3'b001});
  assign MultLoop_acc_1227_nl = nl_MultLoop_acc_1227_nl[21:0];
  assign MultLoop_acc_1227_itm_21_5 = readslicef_22_17_5((MultLoop_acc_1227_nl));
  assign nl_MultLoop_acc_3976_cse_1 = conv_s2u_10_11(data_rsci_idat[287:278]) + 11'b00000000001;
  assign MultLoop_acc_3976_cse_1 = nl_MultLoop_acc_3976_cse_1[10:0];
  assign nl_Result_acc_202_nl =  -conv_s2s_10_11(data_rsci_idat[611:602]);
  assign Result_acc_202_nl = nl_Result_acc_202_nl[10:0];
  assign nl_Result_acc_129_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[611:594]))
      , 2'b01}) + conv_s2s_19_21({(Result_acc_202_nl) , (~ (data_rsci_idat[601:594]))});
  assign Result_acc_129_cse_1 = nl_Result_acc_129_cse_1[20:0];
  assign nl_MultLoop_acc_4094_cse_1 = conv_s2u_13_14(data_rsci_idat[575:563]) + 14'b00000000000001;
  assign MultLoop_acc_4094_cse_1 = nl_MultLoop_acc_4094_cse_1[13:0];
  assign nl_MultLoop_acc_1503_cse_1 = conv_s2s_18_19(data_rsci_idat[89:72]) + conv_s2s_17_19({MultLoop_acc_3925_cse_1
      , (data_rsci_idat[78:74])});
  assign MultLoop_acc_1503_cse_1 = nl_MultLoop_acc_1503_cse_1[18:0];
  assign nl_MultLoop_acc_4590_nl = conv_s2u_19_21(MultLoop_acc_1512_itm_20_2_1) +
      ({(data_rsci_idat[845:828]) , 3'b001});
  assign MultLoop_acc_4590_nl = nl_MultLoop_acc_4590_nl[20:0];
  assign MultLoop_acc_4590_itm_20_5 = readslicef_21_16_5((MultLoop_acc_4590_nl));
  assign nl_MultLoop_acc_471_nl = conv_s2s_18_22(~ (data_rsci_idat[773:756])) + ({(data_rsci_idat[773:756])
      , 4'b0001});
  assign MultLoop_acc_471_nl = nl_MultLoop_acc_471_nl[21:0];
  assign MultLoop_acc_471_itm_21_7 = readslicef_22_15_7((MultLoop_acc_471_nl));
  assign nl_MultLoop_acc_3928_nl = conv_s2s_11_12(data_rsci_idat[647:637]) + 12'b000000000001;
  assign MultLoop_acc_3928_nl = nl_MultLoop_acc_3928_nl[11:0];
  assign nl_MultLoop_acc_1511_nl = (~ (data_rsci_idat[647:630])) + conv_s2s_14_18({(MultLoop_acc_3928_nl)
      , (data_rsci_idat[636:635])});
  assign MultLoop_acc_1511_nl = nl_MultLoop_acc_1511_nl[17:0];
  assign nl_MultLoop_acc_1237_nl = conv_s2u_18_21(MultLoop_acc_1511_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[647:630])) , 2'b01});
  assign MultLoop_acc_1237_nl = nl_MultLoop_acc_1237_nl[20:0];
  assign MultLoop_acc_1237_itm_20_4 = readslicef_21_17_4((MultLoop_acc_1237_nl));
  assign nl_MultLoop_acc_4186_cse_1 = conv_s2u_10_11(data_rsci_idat[449:440]) + 11'b00000000001;
  assign MultLoop_acc_4186_cse_1 = nl_MultLoop_acc_4186_cse_1[10:0];
  assign nl_MultLoop_acc_2781_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[395:378]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[395:378]));
  assign MultLoop_acc_2781_cse_1 = nl_MultLoop_acc_2781_cse_1[21:0];
  assign nl_MultLoop_acc_1940_cse_1 = ({(data_rsci_idat[701:684]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[701:684]));
  assign MultLoop_acc_1940_cse_1 = nl_MultLoop_acc_1940_cse_1[19:0];
  assign nl_MultLoop_acc_4157_nl = conv_s2s_10_11(data_rsci_idat[53:44]) + 11'b00000000001;
  assign MultLoop_acc_4157_nl = nl_MultLoop_acc_4157_nl[10:0];
  assign nl_MultLoop_acc_2337_cse_1 = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_16_19({(MultLoop_acc_4157_nl)
      , (data_rsci_idat[43:39])});
  assign MultLoop_acc_2337_cse_1 = nl_MultLoop_acc_2337_cse_1[18:0];
  assign nl_MultLoop_acc_2669_nl = conv_s2s_20_21({(~ (data_rsci_idat[557:540]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[557:540]));
  assign MultLoop_acc_2669_nl = nl_MultLoop_acc_2669_nl[20:0];
  assign MultLoop_acc_2669_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_2669_nl));
  assign nl_MultLoop_acc_2525_cse_1 = conv_s2s_18_19(data_rsci_idat[629:612]) + conv_s2s_17_19({MultLoop_acc_4084_cse_1
      , (data_rsci_idat[619:614])});
  assign MultLoop_acc_2525_cse_1 = nl_MultLoop_acc_2525_cse_1[18:0];
  assign nl_MultLoop_acc_3986_nl =  -conv_s2s_11_12(data_rsci_idat[593:583]);
  assign MultLoop_acc_3986_nl = nl_MultLoop_acc_3986_nl[11:0];
  assign nl_MultLoop_acc_1866_nl = conv_s2s_20_21({(~ (data_rsci_idat[593:576]))
      , 2'b01}) + conv_s2s_19_21({(MultLoop_acc_3986_nl) , (~ (data_rsci_idat[582:576]))});
  assign MultLoop_acc_1866_nl = nl_MultLoop_acc_1866_nl[20:0];
  assign MultLoop_acc_1866_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1866_nl));
  assign nl_MultLoop_acc_1515_nl = ({(data_rsci_idat[809:792]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_682_18_8
      , (~ (data_rsci_idat[799:792]))});
  assign MultLoop_acc_1515_nl = nl_MultLoop_acc_1515_nl[21:0];
  assign nl_MultLoop_acc_1516_nl = conv_s2s_24_25({(data_rsci_idat[809:792]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_1515_nl);
  assign MultLoop_acc_1516_nl = nl_MultLoop_acc_1516_nl[24:0];
  assign nl_MultLoop_acc_3930_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_1516_nl)))
      + (~ (data_rsci_idat[809:792]));
  assign MultLoop_acc_3930_nl = nl_MultLoop_acc_3930_nl[17:0];
  assign MultLoop_acc_3930_itm_17_2 = readslicef_18_16_2((MultLoop_acc_3930_nl));
  assign nl_Result_acc_216_cse_1 = conv_s2u_11_12(data_rsci_idat[845:835]) + 12'b000000000001;
  assign Result_acc_216_cse_1 = nl_Result_acc_216_cse_1[11:0];
  assign nl_MultLoop_acc_506_nl = conv_s2u_16_18(data_rsci_idat[539:524]) - (data_rsci_idat[539:522]);
  assign MultLoop_acc_506_nl = nl_MultLoop_acc_506_nl[17:0];
  assign MultLoop_acc_506_itm_17_5 = readslicef_18_13_5((MultLoop_acc_506_nl));
  assign nl_MultLoop_acc_4015_cse_1 = conv_s2u_10_11(data_rsci_idat[17:8]) + 11'b00000000001;
  assign MultLoop_acc_4015_cse_1 = nl_MultLoop_acc_4015_cse_1[10:0];
  assign nl_MultLoop_acc_4076_cse_1 = conv_s2u_12_13(data_rsci_idat[755:744]) + 13'b0000000000001;
  assign MultLoop_acc_4076_cse_1 = nl_MultLoop_acc_4076_cse_1[12:0];
  assign nl_MultLoop_acc_4191_cse_1 = conv_s2u_10_11(data_rsci_idat[197:188]) + 11'b00000000001;
  assign MultLoop_acc_4191_cse_1 = nl_MultLoop_acc_4191_cse_1[10:0];
  assign nl_MultLoop_acc_4153_cse_1 = conv_s2u_10_11(data_rsci_idat[161:152]) + 11'b00000000001;
  assign MultLoop_acc_4153_cse_1 = nl_MultLoop_acc_4153_cse_1[10:0];
  assign nl_MultLoop_acc_2340_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_780_18_8
      , (~ (data_rsci_idat[25:18]))});
  assign MultLoop_acc_2340_nl = nl_MultLoop_acc_2340_nl[19:0];
  assign MultLoop_acc_2340_itm_19_4 = readslicef_20_16_4((MultLoop_acc_2340_nl));
  assign nl_MultLoop_acc_4021_cse_1 = conv_s2u_12_13(data_rsci_idat[143:132]) + 13'b0000000000001;
  assign MultLoop_acc_4021_cse_1 = nl_MultLoop_acc_4021_cse_1[12:0];
  assign nl_MultLoop_acc_528_nl = conv_s2s_24_25({(~ (data_rsci_idat[107:90])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[107:90])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[107:90])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_792_18_6
      , (~ (data_rsci_idat[95:90]))});
  assign MultLoop_acc_528_nl = nl_MultLoop_acc_528_nl[24:0];
  assign MultLoop_acc_528_itm_24_10 = readslicef_25_15_10((MultLoop_acc_528_nl));
  assign nl_MultLoop_acc_2500_cse_1 = conv_s2s_18_19(data_rsci_idat[377:360]) + conv_s2s_16_19(data_rsci_idat[377:362]);
  assign MultLoop_acc_2500_cse_1 = nl_MultLoop_acc_2500_cse_1[18:0];
  assign nl_MultLoop_acc_1521_nl = conv_s2s_22_23({(~ (data_rsci_idat[359:342]))
      , 4'b0100}) + conv_s2s_21_23(MultLoop_acc_1520_cse_1);
  assign MultLoop_acc_1521_nl = nl_MultLoop_acc_1521_nl[22:0];
  assign nl_MultLoop_acc_541_nl = conv_s2s_23_24(MultLoop_acc_1521_nl) + ({(data_rsci_idat[359:342])
      , 6'b010000});
  assign MultLoop_acc_541_nl = nl_MultLoop_acc_541_nl[23:0];
  assign MultLoop_acc_541_itm_23_8 = readslicef_24_16_8((MultLoop_acc_541_nl));
  assign nl_MultLoop_acc_1603_cse_1 = conv_s2s_21_22({(~ (data_rsci_idat[521:504]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[521:504]));
  assign MultLoop_acc_1603_cse_1 = nl_MultLoop_acc_1603_cse_1[21:0];
  assign nl_MultLoop_acc_3934_nl = conv_s2s_14_15(data_rsci_idat[269:256]) + 15'b000000000000001;
  assign MultLoop_acc_3934_nl = nl_MultLoop_acc_3934_nl[14:0];
  assign nl_MultLoop_acc_1528_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_17_18({(MultLoop_acc_3934_nl)
      , (data_rsci_idat[255:254])});
  assign MultLoop_acc_1528_nl = nl_MultLoop_acc_1528_nl[17:0];
  assign nl_MultLoop_acc_1275_nl = conv_s2u_18_21(MultLoop_acc_1528_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[269:252])) , 2'b01});
  assign MultLoop_acc_1275_nl = nl_MultLoop_acc_1275_nl[20:0];
  assign MultLoop_acc_1275_itm_20_5 = readslicef_21_16_5((MultLoop_acc_1275_nl));
  assign nl_MultLoop_acc_3933_nl = conv_s2s_13_14(data_rsci_idat[197:185]) + 14'b00000000000001;
  assign MultLoop_acc_3933_nl = nl_MultLoop_acc_3933_nl[13:0];
  assign nl_MultLoop_acc_1526_nl = conv_s2s_18_19(data_rsci_idat[197:180]) + conv_s2s_16_19({(MultLoop_acc_3933_nl)
      , (data_rsci_idat[184:183])});
  assign MultLoop_acc_1526_nl = nl_MultLoop_acc_1526_nl[18:0];
  assign nl_MultLoop_acc_579_nl = conv_s2u_19_20(MultLoop_acc_1526_nl) + ({(~ (data_rsci_idat[197:180]))
      , 2'b00});
  assign MultLoop_acc_579_nl = nl_MultLoop_acc_579_nl[19:0];
  assign MultLoop_acc_579_itm_19_4 = readslicef_20_16_4((MultLoop_acc_579_nl));
  assign nl_Result_acc_127_cse_1 = conv_s2s_18_19(data_rsci_idat[575:558]) + conv_s2s_16_19(data_rsci_idat[575:560]);
  assign Result_acc_127_cse_1 = nl_Result_acc_127_cse_1[18:0];
  assign nl_MultLoop_acc_3955_cse_1 = conv_s2u_11_12(data_rsci_idat[71:61]) + 12'b000000000001;
  assign MultLoop_acc_3955_cse_1 = nl_MultLoop_acc_3955_cse_1[11:0];
  assign nl_MultLoop_acc_4084_cse_1 = conv_s2u_10_11(data_rsci_idat[629:620]) + 11'b00000000001;
  assign MultLoop_acc_4084_cse_1 = nl_MultLoop_acc_4084_cse_1[10:0];
  assign nl_MultLoop_acc_3932_nl = conv_s2s_10_11(data_rsci_idat[35:26]) + 11'b00000000001;
  assign MultLoop_acc_3932_nl = nl_MultLoop_acc_3932_nl[10:0];
  assign nl_MultLoop_acc_1523_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_15_18({(MultLoop_acc_3932_nl)
      , (data_rsci_idat[25:22])});
  assign MultLoop_acc_1523_nl = nl_MultLoop_acc_1523_nl[17:0];
  assign nl_MultLoop_acc_1524_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1523_nl);
  assign MultLoop_acc_1524_nl = nl_MultLoop_acc_1524_nl[19:0];
  assign nl_MultLoop_acc_570_nl = conv_s2u_20_22(MultLoop_acc_1524_nl) + ({(~ (data_rsci_idat[35:18]))
      , 4'b0000});
  assign MultLoop_acc_570_nl = nl_MultLoop_acc_570_nl[21:0];
  assign MultLoop_acc_570_itm_21_6 = readslicef_22_16_6((MultLoop_acc_570_nl));
  assign nl_MultLoop_acc_1741_cse_1 = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_15_19(data_rsci_idat[35:21]);
  assign MultLoop_acc_1741_cse_1 = nl_MultLoop_acc_1741_cse_1[18:0];
  assign nl_MultLoop_acc_3935_nl = conv_s2s_11_12(data_rsci_idat[17:7]) + 12'b000000000001;
  assign MultLoop_acc_3935_nl = nl_MultLoop_acc_3935_nl[11:0];
  assign nl_MultLoop_acc_1531_cse_1 = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_17_19({(MultLoop_acc_3935_nl)
      , (data_rsci_idat[6:2])});
  assign MultLoop_acc_1531_cse_1 = nl_MultLoop_acc_1531_cse_1[18:0];
  assign nl_Result_acc_187_cse_1 = conv_s2u_11_12(data_rsci_idat[125:115]) + 12'b000000000001;
  assign Result_acc_187_cse_1 = nl_Result_acc_187_cse_1[11:0];
  assign nl_MultLoop_acc_2403_cse_1 = (~ (data_rsci_idat[413:396])) + conv_s2s_16_18(data_rsci_idat[413:398]);
  assign MultLoop_acc_2403_cse_1 = nl_MultLoop_acc_2403_cse_1[17:0];
  assign nl_MultLoop_acc_2030_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[809:792]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_690_18_6 , (~ (data_rsci_idat[797:792]))});
  assign MultLoop_acc_2030_cse_1 = nl_MultLoop_acc_2030_cse_1[20:0];
  assign nl_MultLoop_acc_3916_cse_1 = conv_s2u_12_13(data_rsci_idat[719:708]) + 13'b0000000000001;
  assign MultLoop_acc_3916_cse_1 = nl_MultLoop_acc_3916_cse_1[12:0];
  assign nl_MultLoop_acc_4150_cse_1 = conv_s2u_10_11(data_rsci_idat[269:260]) + 11'b00000000001;
  assign MultLoop_acc_4150_cse_1 = nl_MultLoop_acc_4150_cse_1[10:0];
  assign nl_MultLoop_acc_4030_cse_1 = conv_s2u_10_11(data_rsci_idat[467:458]) + 11'b00000000001;
  assign MultLoop_acc_4030_cse_1 = nl_MultLoop_acc_4030_cse_1[10:0];
  assign nl_MultLoop_acc_3987_cse_1 = conv_s2u_10_11(data_rsci_idat[521:512]) + 11'b00000000001;
  assign MultLoop_acc_3987_cse_1 = nl_MultLoop_acc_3987_cse_1[10:0];
  assign nl_MultLoop_acc_2259_cse_1 = (~ (data_rsci_idat[53:36])) + conv_s2s_15_18(data_rsci_idat[53:39]);
  assign MultLoop_acc_2259_cse_1 = nl_MultLoop_acc_2259_cse_1[17:0];
  assign nl_MultLoop_acc_1730_nl = ({(data_rsci_idat[395:378]) , 5'b00001}) + conv_s2s_18_23(~
      (data_rsci_idat[395:378]));
  assign MultLoop_acc_1730_nl = nl_MultLoop_acc_1730_nl[22:0];
  assign MultLoop_acc_1730_itm_22_7 = readslicef_23_16_7((MultLoop_acc_1730_nl));
  assign nl_MultLoop_acc_3925_cse_1 = conv_s2u_11_12(data_rsci_idat[89:79]) + 12'b000000000001;
  assign MultLoop_acc_3925_cse_1 = nl_MultLoop_acc_3925_cse_1[11:0];
  assign nl_Result_acc_163_cse_1 = conv_s2s_18_19(data_rsci_idat[755:738]) + conv_s2s_16_19({Result_acc_214_cse_1
      , (data_rsci_idat[745:741])});
  assign Result_acc_163_cse_1 = nl_Result_acc_163_cse_1[18:0];
  assign nl_MultLoop_acc_1816_nl = conv_s2s_20_21({(~ (data_rsci_idat[197:180]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_862_18_6 , (~ (data_rsci_idat[185:180]))});
  assign MultLoop_acc_1816_nl = nl_MultLoop_acc_1816_nl[20:0];
  assign MultLoop_acc_1816_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1816_nl));
  assign nl_MultLoop_acc_2035_cse_1 = (~ (data_rsci_idat[791:774])) + conv_s2s_16_18(data_rsci_idat[791:776]);
  assign MultLoop_acc_2035_cse_1 = nl_MultLoop_acc_2035_cse_1[17:0];
  assign nl_MultLoop_acc_1532_nl = ({(~ (data_rsci_idat[17:0])) , 3'b000}) + conv_s2s_19_21(MultLoop_acc_1531_cse_1);
  assign MultLoop_acc_1532_nl = nl_MultLoop_acc_1532_nl[20:0];
  assign nl_MultLoop_acc_713_nl = conv_s2u_21_24(MultLoop_acc_1532_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[17:0])) , 5'b01000});
  assign MultLoop_acc_713_nl = nl_MultLoop_acc_713_nl[23:0];
  assign MultLoop_acc_713_itm_23_8 = readslicef_24_16_8((MultLoop_acc_713_nl));
  assign nl_MultLoop_acc_785_nl = conv_s2u_13_18(data_rsci_idat[503:491]) - (data_rsci_idat[503:486]);
  assign MultLoop_acc_785_nl = nl_MultLoop_acc_785_nl[17:0];
  assign MultLoop_acc_785_itm_17_4 = readslicef_18_14_4((MultLoop_acc_785_nl));
  assign nl_MultLoop_acc_4663_nl = conv_s2u_19_20(MultLoop_acc_1715_itm_20_2_1) +
      ({(data_rsci_idat[485:468]) , 2'b01});
  assign MultLoop_acc_4663_nl = nl_MultLoop_acc_4663_nl[19:0];
  assign MultLoop_acc_4663_itm_19_4 = readslicef_20_16_4((MultLoop_acc_4663_nl));
  assign nl_Result_acc_183_cse_1 = conv_s2u_11_12(data_rsci_idat[701:691]) + 12'b000000000001;
  assign Result_acc_183_cse_1 = nl_Result_acc_183_cse_1[11:0];
  assign nl_MultLoop_acc_4075_cse_1 = conv_s2u_12_13(data_rsci_idat[287:276]) + 13'b0000000000001;
  assign MultLoop_acc_4075_cse_1 = nl_MultLoop_acc_4075_cse_1[12:0];
  assign nl_MultLoop_acc_1043_cse_1 = conv_s2s_18_20(~ (data_rsci_idat[17:0])) +
      ({(data_rsci_idat[17:0]) , 2'b01});
  assign MultLoop_acc_1043_cse_1 = nl_MultLoop_acc_1043_cse_1[19:0];
  assign nl_MultLoop_acc_3937_nl =  -conv_s2s_11_12(data_rsci_idat[359:349]);
  assign MultLoop_acc_3937_nl = nl_MultLoop_acc_3937_nl[11:0];
  assign nl_MultLoop_acc_826_nl = conv_s2s_25_26({(~ (data_rsci_idat[359:342])) ,
      7'b0001000}) + conv_s2s_21_26({(~ (data_rsci_idat[359:342])) , 3'b001}) + conv_s2s_19_26({(MultLoop_acc_3937_nl)
      , (~ (data_rsci_idat[348:342]))});
  assign MultLoop_acc_826_nl = nl_MultLoop_acc_826_nl[25:0];
  assign MultLoop_acc_826_itm_25_10 = readslicef_26_16_10((MultLoop_acc_826_nl));
  assign nl_MultLoop_acc_3989_cse_1 = conv_s2u_10_11(data_rsci_idat[305:296]) + 11'b00000000001;
  assign MultLoop_acc_3989_cse_1 = nl_MultLoop_acc_3989_cse_1[10:0];
  assign nl_MultLoop_acc_1735_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[251:234]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[251:234]));
  assign MultLoop_acc_1735_cse_1 = nl_MultLoop_acc_1735_cse_1[20:0];
  assign nl_MultLoop_acc_1479_nl = conv_s2s_18_19(data_rsci_idat[809:792]) + conv_s2s_16_19(data_rsci_idat[809:794]);
  assign MultLoop_acc_1479_nl = nl_MultLoop_acc_1479_nl[18:0];
  assign MultLoop_acc_1479_itm_18_3 = readslicef_19_16_3((MultLoop_acc_1479_nl));
  assign nl_MultLoop_acc_4592_nl = conv_s2u_17_19(MultLoop_acc_4591_itm_18_2) + conv_s2u_18_19(data_rsci_idat[701:684]);
  assign MultLoop_acc_4592_nl = nl_MultLoop_acc_4592_nl[18:0];
  assign MultLoop_acc_4592_itm_18_3 = readslicef_19_16_3((MultLoop_acc_4592_nl));
  assign nl_MultLoop_acc_4593_nl = conv_s2u_16_19(MultLoop_acc_1543_itm_21_6) + conv_s2u_18_19(data_rsci_idat[719:702]);
  assign MultLoop_acc_4593_nl = nl_MultLoop_acc_4593_nl[18:0];
  assign MultLoop_acc_4593_itm_18_3 = readslicef_19_16_3((MultLoop_acc_4593_nl));
  assign nl_MultLoop_acc_1540_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_16_18(data_rsci_idat[377:362]);
  assign MultLoop_acc_1540_nl = nl_MultLoop_acc_1540_nl[17:0];
  assign nl_MultLoop_acc_1350_nl = conv_s2u_18_23(MultLoop_acc_1540_nl) + ({(data_rsci_idat[377:360])
      , 5'b00001});
  assign MultLoop_acc_1350_nl = nl_MultLoop_acc_1350_nl[22:0];
  assign MultLoop_acc_1350_itm_22_7 = readslicef_23_16_7((MultLoop_acc_1350_nl));
  assign nl_MultLoop_acc_1537_nl = ({(~ (data_rsci_idat[17:0])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[17:0])
      + conv_s2s_15_20(data_rsci_idat[17:3]);
  assign MultLoop_acc_1537_nl = nl_MultLoop_acc_1537_nl[19:0];
  assign nl_MultLoop_acc_807_nl = conv_s2u_20_22(MultLoop_acc_1537_nl) + ({(data_rsci_idat[17:0])
      , 4'b0100});
  assign MultLoop_acc_807_nl = nl_MultLoop_acc_807_nl[21:0];
  assign MultLoop_acc_807_itm_21_6 = readslicef_22_16_6((MultLoop_acc_807_nl));
  assign nl_MultLoop_acc_1957_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[647:630]))
      , 2'b01}) + conv_s2s_19_21({MultLoop_MultLoop_conc_754_18_6 , (~ (data_rsci_idat[635:630]))});
  assign MultLoop_acc_1957_cse_1 = nl_MultLoop_acc_1957_cse_1[20:0];
  assign nl_MultLoop_acc_1723_cse_1 = ({(data_rsci_idat[773:756]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[773:756]));
  assign MultLoop_acc_1723_cse_1 = nl_MultLoop_acc_1723_cse_1[19:0];
  assign nl_MultLoop_acc_1727_cse_1 = conv_s2s_18_19(data_rsci_idat[575:558]) + conv_s2s_15_19(data_rsci_idat[575:561]);
  assign MultLoop_acc_1727_cse_1 = nl_MultLoop_acc_1727_cse_1[18:0];
  assign nl_MultLoop_acc_1512_nl = conv_s2s_20_21({(~ (data_rsci_idat[845:828]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[845:828]));
  assign MultLoop_acc_1512_nl = nl_MultLoop_acc_1512_nl[20:0];
  assign MultLoop_acc_1512_itm_20_2_1 = readslicef_21_19_2((MultLoop_acc_1512_nl));
  assign nl_Result_acc_102_nl = conv_s2s_20_21({(~ (data_rsci_idat[521:504])) , 2'b01})
      + conv_s2s_18_21(~ (data_rsci_idat[521:504]));
  assign Result_acc_102_nl = nl_Result_acc_102_nl[20:0];
  assign Result_acc_102_itm_20_2_1 = readslicef_21_19_2((Result_acc_102_nl));
  assign nl_MultLoop_acc_1993_nl = conv_s2s_18_19(data_rsci_idat[683:666]) + conv_s2s_13_19(data_rsci_idat[683:671]);
  assign MultLoop_acc_1993_nl = nl_MultLoop_acc_1993_nl[18:0];
  assign MultLoop_acc_1993_itm_18_2 = readslicef_19_17_2((MultLoop_acc_1993_nl));
  assign nl_MultLoop_acc_4036_cse_1 = conv_s2u_11_12(data_rsci_idat[197:187]) + 12'b000000000001;
  assign MultLoop_acc_4036_cse_1 = nl_MultLoop_acc_4036_cse_1[11:0];
  assign nl_MultLoop_acc_3938_nl =  -conv_s2s_14_15(data_rsci_idat[35:22]);
  assign MultLoop_acc_3938_nl = nl_MultLoop_acc_3938_nl[14:0];
  assign nl_MultLoop_acc_856_nl = conv_s2s_19_23({(MultLoop_acc_3938_nl) , (~ (data_rsci_idat[21:18]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[35:18])) , 4'b0001});
  assign MultLoop_acc_856_nl = nl_MultLoop_acc_856_nl[22:0];
  assign MultLoop_acc_856_itm_22_7 = readslicef_23_16_7((MultLoop_acc_856_nl));
  assign nl_MultLoop_acc_1626_cse_1 = (~ (data_rsci_idat[287:270])) + conv_s2s_16_18(data_rsci_idat[287:272]);
  assign MultLoop_acc_1626_cse_1 = nl_MultLoop_acc_1626_cse_1[17:0];
  assign nl_MultLoop_acc_1844_cse_1 = (~ (data_rsci_idat[161:144])) + conv_s2s_16_18(data_rsci_idat[161:146]);
  assign MultLoop_acc_1844_cse_1 = nl_MultLoop_acc_1844_cse_1[17:0];
  assign nl_MultLoop_acc_1702_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[431:414]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_1702_cse_1 = nl_MultLoop_acc_1702_cse_1[20:0];
  assign nl_Result_acc_154_nl = ({(data_rsci_idat[683:666]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[683:666]));
  assign Result_acc_154_nl = nl_Result_acc_154_nl[19:0];
  assign Result_acc_154_itm_19_4 = readslicef_20_16_4((Result_acc_154_nl));
  assign nl_MultLoop_acc_4591_nl = conv_s2u_18_19(data_rsci_idat[701:684]) + conv_s2u_17_19(MultLoop_acc_1541_itm_18_2);
  assign MultLoop_acc_4591_nl = nl_MultLoop_acc_4591_nl[18:0];
  assign MultLoop_acc_4591_itm_18_2 = readslicef_19_17_2((MultLoop_acc_4591_nl));
  assign nl_MultLoop_acc_1520_cse_1 = conv_s2s_20_21({(~ (data_rsci_idat[359:342]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[359:342]));
  assign MultLoop_acc_1520_cse_1 = nl_MultLoop_acc_1520_cse_1[20:0];
  assign nl_MultLoop_MultLoop_conc_674_18_5 =  -conv_s2s_13_14(data_rsci_idat[305:293]);
  assign MultLoop_MultLoop_conc_674_18_5 = nl_MultLoop_MultLoop_conc_674_18_5[13:0];
  assign nl_MultLoop_MultLoop_conc_676_18_6 =  -conv_s2s_12_13(data_rsci_idat[791:780]);
  assign MultLoop_MultLoop_conc_676_18_6 = nl_MultLoop_MultLoop_conc_676_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_678_18_7 =  -conv_s2s_11_12(data_rsci_idat[467:457]);
  assign MultLoop_MultLoop_conc_678_18_7 = nl_MultLoop_MultLoop_conc_678_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_680_16_6 = conv_s2s_10_11(data_rsci_idat[431:422])
      + 11'b00000000001;
  assign MultLoop_MultLoop_conc_680_16_6 = nl_MultLoop_MultLoop_conc_680_16_6[10:0];
  assign nl_MultLoop_MultLoop_conc_682_18_8 =  -conv_s2s_10_11(data_rsci_idat[809:800]);
  assign MultLoop_MultLoop_conc_682_18_8 = nl_MultLoop_MultLoop_conc_682_18_8[10:0];
  assign nl_MultLoop_acc_4133_itm =  -conv_s2s_11_12(data_rsci_idat[827:817]);
  assign MultLoop_acc_4133_itm = nl_MultLoop_acc_4133_itm[11:0];
  assign nl_MultLoop_MultLoop_conc_686_18_6 =  -conv_s2s_12_13(data_rsci_idat[575:564]);
  assign MultLoop_MultLoop_conc_686_18_6 = nl_MultLoop_MultLoop_conc_686_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_688_18_7 =  -conv_s2s_11_12(data_rsci_idat[773:763]);
  assign MultLoop_MultLoop_conc_688_18_7 = nl_MultLoop_MultLoop_conc_688_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_690_18_6 =  -conv_s2s_12_13(data_rsci_idat[809:798]);
  assign MultLoop_MultLoop_conc_690_18_6 = nl_MultLoop_MultLoop_conc_690_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_692_18_7 =  -conv_s2s_11_12(data_rsci_idat[485:475]);
  assign MultLoop_MultLoop_conc_692_18_7 = nl_MultLoop_MultLoop_conc_692_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_694_15_3 = conv_s2s_12_13(data_rsci_idat[107:96])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_694_15_3 = nl_MultLoop_MultLoop_conc_694_15_3[12:0];
  assign nl_MultLoop_MultLoop_conc_696_18_7 =  -conv_s2s_11_12(data_rsci_idat[845:835]);
  assign MultLoop_MultLoop_conc_696_18_7 = nl_MultLoop_MultLoop_conc_696_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_698_18_7 =  -conv_s2s_11_12(data_rsci_idat[197:187]);
  assign MultLoop_MultLoop_conc_698_18_7 = nl_MultLoop_MultLoop_conc_698_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_700_18_7 =  -conv_s2s_11_12(data_rsci_idat[557:547]);
  assign MultLoop_MultLoop_conc_700_18_7 = nl_MultLoop_MultLoop_conc_700_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_702_18_6 =  -conv_s2s_12_13(data_rsci_idat[233:222]);
  assign MultLoop_MultLoop_conc_702_18_6 = nl_MultLoop_MultLoop_conc_702_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_704_18_6 =  -conv_s2s_12_13(data_rsci_idat[593:582]);
  assign MultLoop_MultLoop_conc_704_18_6 = nl_MultLoop_MultLoop_conc_704_18_6[12:0];
  assign nl_MultLoop_acc_4688 = conv_s2s_20_21({(~ (data_rsci_idat[629:612])) , 2'b01})
      + conv_s2s_18_21(~ (data_rsci_idat[629:612]));
  assign MultLoop_acc_4688 = nl_MultLoop_acc_4688[20:0];
  assign nl_MultLoop_MultLoop_conc_706_16_4 = conv_s2s_12_13(data_rsci_idat[305:294])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_706_16_4 = nl_MultLoop_MultLoop_conc_706_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_708_18_6 =  -conv_s2s_12_13(data_rsci_idat[17:6]);
  assign MultLoop_MultLoop_conc_708_18_6 = nl_MultLoop_MultLoop_conc_708_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_714_15_2 = conv_s2s_13_14(data_rsci_idat[737:725])
      + 14'b00000000000001;
  assign MultLoop_MultLoop_conc_714_15_2 = nl_MultLoop_MultLoop_conc_714_15_2[13:0];
  assign nl_MultLoop_MultLoop_conc_716_18_7 =  -conv_s2s_11_12(data_rsci_idat[503:493]);
  assign MultLoop_MultLoop_conc_716_18_7 = nl_MultLoop_MultLoop_conc_716_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_718_18_8 =  -conv_s2s_10_11(data_rsci_idat[179:170]);
  assign MultLoop_MultLoop_conc_718_18_8 = nl_MultLoop_MultLoop_conc_718_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_720_18_7 =  -conv_s2s_11_12(data_rsci_idat[863:853]);
  assign MultLoop_MultLoop_conc_720_18_7 = nl_MultLoop_MultLoop_conc_720_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_722_18_8 =  -conv_s2s_10_11(data_rsci_idat[413:404]);
  assign MultLoop_MultLoop_conc_722_18_8 = nl_MultLoop_MultLoop_conc_722_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_724_18_6 =  -conv_s2s_12_13(data_rsci_idat[485:474]);
  assign MultLoop_MultLoop_conc_724_18_6 = nl_MultLoop_MultLoop_conc_724_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_726_18_7 =  -conv_s2s_11_12(data_rsci_idat[521:511]);
  assign MultLoop_MultLoop_conc_726_18_7 = nl_MultLoop_MultLoop_conc_726_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_728_18_8 =  -conv_s2s_10_11(data_rsci_idat[863:854]);
  assign MultLoop_MultLoop_conc_728_18_8 = nl_MultLoop_MultLoop_conc_728_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_730_18_7 =  -conv_s2s_11_12(data_rsci_idat[233:223]);
  assign MultLoop_MultLoop_conc_730_18_7 = nl_MultLoop_MultLoop_conc_730_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_732_14_2 = conv_s2s_12_13(data_rsci_idat[539:528])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_732_14_2 = nl_MultLoop_MultLoop_conc_732_14_2[12:0];
  assign nl_MultLoop_MultLoop_conc_734_18_7 =  -conv_s2s_11_12(data_rsci_idat[305:295]);
  assign MultLoop_MultLoop_conc_734_18_7 = nl_MultLoop_MultLoop_conc_734_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_736_16_5 = conv_s2s_11_12(data_rsci_idat[377:367])
      + 12'b000000000001;
  assign MultLoop_MultLoop_conc_736_16_5 = nl_MultLoop_MultLoop_conc_736_16_5[11:0];
  assign nl_MultLoop_MultLoop_conc_738_18_4 =  -conv_s2s_14_15(data_rsci_idat[791:778]);
  assign MultLoop_MultLoop_conc_738_18_4 = nl_MultLoop_MultLoop_conc_738_18_4[14:0];
  assign nl_MultLoop_MultLoop_conc_740_16_4 = conv_s2s_12_13(data_rsci_idat[791:780])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_740_16_4 = nl_MultLoop_MultLoop_conc_740_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_742_18_6 =  -conv_s2s_12_13(data_rsci_idat[503:492]);
  assign MultLoop_MultLoop_conc_742_18_6 = nl_MultLoop_MultLoop_conc_742_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_746_18_8 =  -conv_s2s_10_11(data_rsci_idat[215:206]);
  assign MultLoop_MultLoop_conc_746_18_8 = nl_MultLoop_MultLoop_conc_746_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_750_18_7 =  -conv_s2s_11_12(data_rsci_idat[611:601]);
  assign MultLoop_MultLoop_conc_750_18_7 = nl_MultLoop_MultLoop_conc_750_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_752_18_6 =  -conv_s2s_12_13(data_rsci_idat[287:276]);
  assign MultLoop_MultLoop_conc_752_18_6 = nl_MultLoop_MultLoop_conc_752_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_754_18_6 =  -conv_s2s_12_13(data_rsci_idat[647:636]);
  assign MultLoop_MultLoop_conc_754_18_6 = nl_MultLoop_MultLoop_conc_754_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_756_18_8 =  -conv_s2s_10_11(data_rsci_idat[665:656]);
  assign MultLoop_MultLoop_conc_756_18_8 = nl_MultLoop_MultLoop_conc_756_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_758_18_6 =  -conv_s2s_12_13(data_rsci_idat[71:60]);
  assign MultLoop_MultLoop_conc_758_18_6 = nl_MultLoop_MultLoop_conc_758_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_760_18_5 =  -conv_s2s_13_14(data_rsci_idat[773:761]);
  assign MultLoop_MultLoop_conc_760_18_5 = nl_MultLoop_MultLoop_conc_760_18_5[13:0];
  assign nl_MultLoop_MultLoop_conc_766_18_7 =  -conv_s2s_11_12(data_rsci_idat[629:619]);
  assign MultLoop_MultLoop_conc_766_18_7 = nl_MultLoop_MultLoop_conc_766_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_768_15_2 = conv_s2s_13_14(data_rsci_idat[449:437])
      + 14'b00000000000001;
  assign MultLoop_MultLoop_conc_768_15_2 = nl_MultLoop_MultLoop_conc_768_15_2[13:0];
  assign nl_MultLoop_MultLoop_conc_770_18_8 =  -conv_s2s_10_11(data_rsci_idat[251:242]);
  assign MultLoop_MultLoop_conc_770_18_8 = nl_MultLoop_MultLoop_conc_770_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_772_16_2 = conv_s2s_14_15(data_rsci_idat[593:580])
      + 15'b000000000000001;
  assign MultLoop_MultLoop_conc_772_16_2 = nl_MultLoop_MultLoop_conc_772_16_2[14:0];
  assign nl_MultLoop_MultLoop_conc_774_16_4 = conv_s2s_12_13(data_rsci_idat[611:600])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_774_16_4 = nl_MultLoop_MultLoop_conc_774_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_776_15_4 = conv_s2s_11_12(data_rsci_idat[611:601])
      + 12'b000000000001;
  assign MultLoop_MultLoop_conc_776_15_4 = nl_MultLoop_MultLoop_conc_776_15_4[11:0];
  assign nl_MultLoop_MultLoop_conc_778_16_6 = conv_s2s_10_11(data_rsci_idat[323:314])
      + 11'b00000000001;
  assign MultLoop_MultLoop_conc_778_16_6 = nl_MultLoop_MultLoop_conc_778_16_6[10:0];
  assign nl_MultLoop_MultLoop_conc_780_18_8 =  -conv_s2s_10_11(data_rsci_idat[35:26]);
  assign MultLoop_MultLoop_conc_780_18_8 = nl_MultLoop_MultLoop_conc_780_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_782_18_8 =  -conv_s2s_10_11(data_rsci_idat[701:692]);
  assign MultLoop_MultLoop_conc_782_18_8 = nl_MultLoop_MultLoop_conc_782_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_784_16_6 = conv_s2s_10_11(data_rsci_idat[683:674])
      + 11'b00000000001;
  assign MultLoop_MultLoop_conc_784_16_6 = nl_MultLoop_MultLoop_conc_784_16_6[10:0];
  assign nl_MultLoop_MultLoop_conc_786_18_7 =  -conv_s2s_11_12(data_rsci_idat[71:61]);
  assign MultLoop_MultLoop_conc_786_18_7 = nl_MultLoop_MultLoop_conc_786_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_788_18_5 =  -conv_s2s_13_14(data_rsci_idat[431:419]);
  assign MultLoop_MultLoop_conc_788_18_5 = nl_MultLoop_MultLoop_conc_788_18_5[13:0];
  assign nl_MultLoop_MultLoop_conc_790_16_4 = conv_s2s_12_13(data_rsci_idat[395:384])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_790_16_4 = nl_MultLoop_MultLoop_conc_790_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_792_18_6 =  -conv_s2s_12_13(data_rsci_idat[107:96]);
  assign MultLoop_MultLoop_conc_792_18_6 = nl_MultLoop_MultLoop_conc_792_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_794_16_5 = conv_s2s_11_12(data_rsci_idat[431:421])
      + 12'b000000000001;
  assign MultLoop_MultLoop_conc_794_16_5 = nl_MultLoop_MultLoop_conc_794_16_5[11:0];
  assign nl_MultLoop_MultLoop_conc_796_18_8 =  -conv_s2s_10_11(data_rsci_idat[485:476]);
  assign MultLoop_MultLoop_conc_796_18_8 = nl_MultLoop_MultLoop_conc_796_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_798_16_4 = conv_s2s_12_13(data_rsci_idat[179:168])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_798_16_4 = nl_MultLoop_MultLoop_conc_798_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_800_18_7 =  -conv_s2s_11_12(data_rsci_idat[377:367]);
  assign MultLoop_MultLoop_conc_800_18_7 = nl_MultLoop_MultLoop_conc_800_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_802_18_8 =  -conv_s2s_10_11(data_rsci_idat[53:44]);
  assign MultLoop_MultLoop_conc_802_18_8 = nl_MultLoop_MultLoop_conc_802_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_804_18_7 =  -conv_s2s_11_12(data_rsci_idat[89:79]);
  assign MultLoop_MultLoop_conc_804_18_7 = nl_MultLoop_MultLoop_conc_804_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_806_18_5 =  -conv_s2s_13_14(data_rsci_idat[449:437]);
  assign MultLoop_MultLoop_conc_806_18_5 = nl_MultLoop_MultLoop_conc_806_18_5[13:0];
  assign nl_MultLoop_acc_4690 = conv_s2s_22_23({(~ (data_rsci_idat[161:144])) , 4'b0001})
      + conv_s2s_18_23(~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_4690 = nl_MultLoop_acc_4690[22:0];
  assign nl_MultLoop_MultLoop_conc_810_15_2 = conv_s2s_13_14(data_rsci_idat[485:473])
      + 14'b00000000000001;
  assign MultLoop_MultLoop_conc_810_15_2 = nl_MultLoop_MultLoop_conc_810_15_2[13:0];
  assign nl_MultLoop_MultLoop_conc_814_18_8 =  -conv_s2s_10_11(data_rsci_idat[287:278]);
  assign MultLoop_MultLoop_conc_814_18_8 = nl_MultLoop_MultLoop_conc_814_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_816_18_7 =  -conv_s2s_11_12(data_rsci_idat[683:673]);
  assign MultLoop_MultLoop_conc_816_18_7 = nl_MultLoop_MultLoop_conc_816_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_818_18_7 =  -conv_s2s_11_12(data_rsci_idat[395:385]);
  assign MultLoop_MultLoop_conc_818_18_7 = nl_MultLoop_MultLoop_conc_818_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_820_18_8 =  -conv_s2s_10_11(data_rsci_idat[737:728]);
  assign MultLoop_MultLoop_conc_820_18_8 = nl_MultLoop_MultLoop_conc_820_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_822_18_7 =  -conv_s2s_11_12(data_rsci_idat[107:97]);
  assign MultLoop_MultLoop_conc_822_18_7 = nl_MultLoop_MultLoop_conc_822_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_824_18_6 =  -conv_s2s_12_13(data_rsci_idat[143:132]);
  assign MultLoop_MultLoop_conc_824_18_6 = nl_MultLoop_MultLoop_conc_824_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_826_18_5 =  -conv_s2s_13_14(data_rsci_idat[179:167]);
  assign MultLoop_MultLoop_conc_826_18_5 = nl_MultLoop_MultLoop_conc_826_18_5[13:0];
  assign nl_MultLoop_MultLoop_conc_828_18_7 =  -conv_s2s_11_12(data_rsci_idat[701:691]);
  assign MultLoop_MultLoop_conc_828_18_7 = nl_MultLoop_MultLoop_conc_828_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_830_18_6 =  -conv_s2s_12_13(data_rsci_idat[737:726]);
  assign MultLoop_MultLoop_conc_830_18_6 = nl_MultLoop_MultLoop_conc_830_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_832_18_7 =  -conv_s2s_11_12(data_rsci_idat[125:115]);
  assign MultLoop_MultLoop_conc_832_18_7 = nl_MultLoop_MultLoop_conc_832_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_834_18_5 =  -conv_s2s_13_14(data_rsci_idat[647:635]);
  assign MultLoop_MultLoop_conc_834_18_5 = nl_MultLoop_MultLoop_conc_834_18_5[13:0];
  assign nl_MultLoop_MultLoop_conc_836_18_8 =  -conv_s2s_10_11(data_rsci_idat[323:314]);
  assign MultLoop_MultLoop_conc_836_18_8 = nl_MultLoop_MultLoop_conc_836_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_838_18_4 =  -conv_s2s_14_15(data_rsci_idat[683:670]);
  assign MultLoop_MultLoop_conc_838_18_4 = nl_MultLoop_MultLoop_conc_838_18_4[14:0];
  assign nl_MultLoop_MultLoop_conc_840_18_7 =  -conv_s2s_11_12(data_rsci_idat[719:709]);
  assign MultLoop_MultLoop_conc_840_18_7 = nl_MultLoop_MultLoop_conc_840_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_842_18_6 =  -conv_s2s_12_13(data_rsci_idat[755:744]);
  assign MultLoop_MultLoop_conc_842_18_6 = nl_MultLoop_MultLoop_conc_842_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_844_18_7 =  -conv_s2s_11_12(data_rsci_idat[431:421]);
  assign MultLoop_MultLoop_conc_844_18_7 = nl_MultLoop_MultLoop_conc_844_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_846_18_8 =  -conv_s2s_10_11(data_rsci_idat[773:764]);
  assign MultLoop_MultLoop_conc_846_18_8 = nl_MultLoop_MultLoop_conc_846_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_848_18_7 =  -conv_s2s_11_12(data_rsci_idat[143:133]);
  assign MultLoop_MultLoop_conc_848_18_7 = nl_MultLoop_MultLoop_conc_848_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_850_18_6 =  -conv_s2s_12_13(data_rsci_idat[179:168]);
  assign MultLoop_MultLoop_conc_850_18_6 = nl_MultLoop_MultLoop_conc_850_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_852_18_6 =  -conv_s2s_12_13(data_rsci_idat[539:528]);
  assign MultLoop_MultLoop_conc_852_18_6 = nl_MultLoop_MultLoop_conc_852_18_6[12:0];
  assign nl_MultLoop_MultLoop_conc_854_18_8 =  -conv_s2s_10_11(data_rsci_idat[341:332]);
  assign MultLoop_MultLoop_conc_854_18_8 = nl_MultLoop_MultLoop_conc_854_18_8[10:0];
  assign nl_MultLoop_MultLoop_conc_856_18_7 =  -conv_s2s_11_12(data_rsci_idat[737:727]);
  assign MultLoop_MultLoop_conc_856_18_7 = nl_MultLoop_MultLoop_conc_856_18_7[11:0];
  assign nl_MultLoop_acc_4692 = ({(data_rsci_idat[449:432]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[449:432]));
  assign MultLoop_acc_4692 = nl_MultLoop_acc_4692[19:0];
  assign nl_MultLoop_MultLoop_conc_858_18_7 =  -conv_s2s_11_12(data_rsci_idat[809:799]);
  assign MultLoop_MultLoop_conc_858_18_7 = nl_MultLoop_MultLoop_conc_858_18_7[11:0];
  assign nl_MultLoop_MultLoop_conc_860_16_4 = conv_s2s_12_13(data_rsci_idat[485:474])
      + 13'b0000000000001;
  assign MultLoop_MultLoop_conc_860_16_4 = nl_MultLoop_MultLoop_conc_860_16_4[12:0];
  assign nl_MultLoop_MultLoop_conc_862_18_6 =  -conv_s2s_12_13(data_rsci_idat[197:186]);
  assign MultLoop_MultLoop_conc_862_18_6 = nl_MultLoop_MultLoop_conc_862_18_6[12:0];
  assign nl_MultLoop_acc_150_nl = conv_s2u_13_18(data_rsci_idat[107:95]) - (data_rsci_idat[107:90]);
  assign MultLoop_acc_150_nl = nl_MultLoop_acc_150_nl[17:0];
  assign MultLoop_acc_150_itm_17_4 = readslicef_18_14_4((MultLoop_acc_150_nl));
  assign nl_MultLoop_acc_1497_nl = (~ (data_rsci_idat[719:702])) + conv_s2s_16_18({MultLoop_acc_3916_cse_1
      , (data_rsci_idat[707:705])});
  assign MultLoop_acc_1497_nl = nl_MultLoop_acc_1497_nl[17:0];
  assign nl_MultLoop_acc_1191_nl = conv_s2u_18_22(MultLoop_acc_1497_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[719:702])) , 3'b001});
  assign MultLoop_acc_1191_nl = nl_MultLoop_acc_1191_nl[21:0];
  assign MultLoop_acc_1191_itm_21_7 = readslicef_22_15_7((MultLoop_acc_1191_nl));
  assign nl_MultLoop_acc_1504_nl = ({(~ (data_rsci_idat[89:72])) , 3'b000}) + conv_s2s_19_21(MultLoop_acc_1503_cse_1);
  assign MultLoop_acc_1504_nl = nl_MultLoop_acc_1504_nl[20:0];
  assign nl_MultLoop_acc_1211_nl = conv_s2u_21_24(MultLoop_acc_1504_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[89:72])) , 5'b01000});
  assign MultLoop_acc_1211_nl = nl_MultLoop_acc_1211_nl[23:0];
  assign MultLoop_acc_1211_itm_23_8 = readslicef_24_16_8((MultLoop_acc_1211_nl));
  assign nl_MultLoop_acc_1513_nl = (~ (data_rsci_idat[215:198])) + conv_s2s_16_18(data_rsci_idat[215:200]);
  assign MultLoop_acc_1513_nl = nl_MultLoop_acc_1513_nl[17:0];
  assign nl_MultLoop_acc_1243_nl = conv_s2u_18_20(MultLoop_acc_1513_nl) + ({(data_rsci_idat[215:198])
      , 2'b01});
  assign MultLoop_acc_1243_nl = nl_MultLoop_acc_1243_nl[19:0];
  assign MultLoop_acc_1243_itm_19_6 = readslicef_20_14_6((MultLoop_acc_1243_nl));
  assign nl_MultLoop_asn_1479 = (~ (data_rsci_idat[683:666])) + conv_s2s_16_18(Result_acc_154_itm_19_4);
  assign MultLoop_asn_1479 = nl_MultLoop_asn_1479[17:0];
  assign nl_MultLoop_acc_1529_nl = (~ (data_rsci_idat[863:846])) + conv_s2s_16_18(data_rsci_idat[863:848]);
  assign MultLoop_acc_1529_nl = nl_MultLoop_acc_1529_nl[17:0];
  assign nl_MultLoop_acc_1315_nl = conv_s2u_18_20(MultLoop_acc_1529_nl) + ({(data_rsci_idat[863:846])
      , 2'b01});
  assign MultLoop_acc_1315_nl = nl_MultLoop_acc_1315_nl[19:0];
  assign MultLoop_acc_1315_itm_19_4 = readslicef_20_16_4((MultLoop_acc_1315_nl));
  assign nl_MultLoop_acc_3936_nl = conv_s2s_12_13(data_rsci_idat[647:636]) + 13'b0000000000001;
  assign MultLoop_acc_3936_nl = nl_MultLoop_acc_3936_nl[12:0];
  assign nl_MultLoop_acc_1534_nl = (~ (data_rsci_idat[647:630])) + conv_s2s_17_18({(MultLoop_acc_3936_nl)
      , (data_rsci_idat[635:632])});
  assign MultLoop_acc_1534_nl = nl_MultLoop_acc_1534_nl[17:0];
  assign nl_MultLoop_acc_1535_nl = conv_s2s_20_21({(~ (data_rsci_idat[647:630]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1534_nl);
  assign MultLoop_acc_1535_nl = nl_MultLoop_acc_1535_nl[20:0];
  assign nl_MultLoop_acc_1324_nl = conv_s2u_21_23(MultLoop_acc_1535_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[647:630])) , 4'b0100});
  assign MultLoop_acc_1324_nl = nl_MultLoop_acc_1324_nl[22:0];
  assign MultLoop_acc_1324_itm_22_7 = readslicef_23_16_7((MultLoop_acc_1324_nl));
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      res_rsci_d_431_414 <= 18'b000000000000000000;
      res_rsci_d_17_0 <= 18'b000000000000000000;
      res_rsci_d_413_396 <= 18'b000000000000000000;
      res_rsci_d_35_18 <= 18'b000000000000000000;
      res_rsci_d_395_378 <= 18'b000000000000000000;
      res_rsci_d_53_36 <= 18'b000000000000000000;
      res_rsci_d_377_360 <= 18'b000000000000000000;
      res_rsci_d_71_54 <= 18'b000000000000000000;
      res_rsci_d_359_342 <= 18'b000000000000000000;
      res_rsci_d_89_72 <= 18'b000000000000000000;
      res_rsci_d_341_324 <= 18'b000000000000000000;
      res_rsci_d_107_90 <= 18'b000000000000000000;
      res_rsci_d_323_306 <= 18'b000000000000000000;
      res_rsci_d_125_108 <= 18'b000000000000000000;
      res_rsci_d_305_288 <= 18'b000000000000000000;
      res_rsci_d_143_126 <= 18'b000000000000000000;
      res_rsci_d_287_270 <= 18'b000000000000000000;
      res_rsci_d_161_144 <= 18'b000000000000000000;
      res_rsci_d_269_252 <= 18'b000000000000000000;
      res_rsci_d_179_162 <= 18'b000000000000000000;
      res_rsci_d_251_234 <= 18'b000000000000000000;
      res_rsci_d_197_180 <= 18'b000000000000000000;
      res_rsci_d_233_216 <= 18'b000000000000000000;
      res_rsci_d_215_198 <= 18'b000000000000000000;
      MultLoop_acc_1588_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1578_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1562_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1561_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1576_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1575_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1585_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1590_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1582_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1581_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3913_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3881_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3880_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3896_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3895_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3894_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3911_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3910_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1683_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1673_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1659_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1658_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1671_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1670_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1669_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1668_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1685_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1677_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1676_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1800_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1772_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1771_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1783_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1782_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1781_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1780_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1779_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1791_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1797_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3720_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3719_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3718_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3717_itm_1_16_0 <= 17'b00000000000000000;
      MultLoop_acc_3716_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3715_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3725_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3724_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3710_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3709_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3722_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3706_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3705_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1911_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1910_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1918_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1917_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1916_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1889_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1888_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_1902_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_1914_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_1920_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3614_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3598_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3584_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3583_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3596_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3595_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3594_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3593_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3605_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3611_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3495_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3494_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3469_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3468_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3482_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3481_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3480_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3479_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3478_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3490_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3496_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2120_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2119_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2118_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2091_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2090_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2105_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2104_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2103_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2115_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2121_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3378_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3368_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3367_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3366_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3365_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3375_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3362_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3361_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3373_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3379_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_23_7_itm_1
          <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3264_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3258_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3233_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3232_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3245_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3256_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3255_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3254_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3238_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3237_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0 <=
          17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_26_10_itm_1
          <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_acc_1215_22_6_itm_1
          <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1 <= 15'b000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1 <= 15'b000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2470_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2469_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2458_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2457_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2438_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2437_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2455_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2466_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2452_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2451_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2464_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2463_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3018_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3008_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2984_itm_1 <= 15'b000000000000000;
      MultLoop_acc_2983_itm_1 <= 15'b000000000000000;
      MultLoop_acc_2993_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_3006_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3005_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3004_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3003_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_3020_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3012_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_3011_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0 <=
          17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1 <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_25_10_itm_1
          <= 16'b0000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1 <= 17'b00000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1 <= 18'b000000000000000000;
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2888_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2887_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2886_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2871_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2870_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2884_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2883_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2893_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2898_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2897_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2658_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2657_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2656_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2631_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2630_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2643_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2642_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2641_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2653_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2659_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2773_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2750_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2749_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2748_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2747_itm_1 <= 16'b0000000000000000;
      MultLoop_acc_2761_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2760_itm_1 <= 17'b00000000000000000;
      MultLoop_acc_2770_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2775_itm_1 <= 18'b000000000000000000;
      MultLoop_acc_2774_itm_1 <= 18'b000000000000000000;
    end
    else if ( ccs_ccore_en ) begin
      res_rsci_d_431_414 <= nl_res_rsci_d_431_414[17:0];
      res_rsci_d_17_0 <= nl_res_rsci_d_17_0[17:0];
      res_rsci_d_413_396 <= nl_res_rsci_d_413_396[17:0];
      res_rsci_d_35_18 <= nl_res_rsci_d_35_18[17:0];
      res_rsci_d_395_378 <= nl_res_rsci_d_395_378[17:0];
      res_rsci_d_53_36 <= nl_res_rsci_d_53_36[17:0];
      res_rsci_d_377_360 <= nl_res_rsci_d_377_360[17:0];
      res_rsci_d_71_54 <= nl_res_rsci_d_71_54[17:0];
      res_rsci_d_359_342 <= nl_res_rsci_d_359_342[17:0];
      res_rsci_d_89_72 <= nl_res_rsci_d_89_72[17:0];
      res_rsci_d_341_324 <= nl_res_rsci_d_341_324[17:0];
      res_rsci_d_107_90 <= nl_res_rsci_d_107_90[17:0];
      res_rsci_d_323_306 <= nl_res_rsci_d_323_306[17:0];
      res_rsci_d_125_108 <= nl_res_rsci_d_125_108[17:0];
      res_rsci_d_305_288 <= nl_res_rsci_d_305_288[17:0];
      res_rsci_d_143_126 <= nl_res_rsci_d_143_126[17:0];
      res_rsci_d_287_270 <= nl_res_rsci_d_287_270[17:0];
      res_rsci_d_161_144 <= nl_res_rsci_d_161_144[17:0];
      res_rsci_d_269_252 <= nl_res_rsci_d_269_252[17:0];
      res_rsci_d_179_162 <= nl_res_rsci_d_179_162[17:0];
      res_rsci_d_251_234 <= nl_res_rsci_d_251_234[17:0];
      res_rsci_d_197_180 <= nl_res_rsci_d_197_180[17:0];
      res_rsci_d_233_216 <= nl_res_rsci_d_233_216[17:0];
      res_rsci_d_215_198 <= nl_res_rsci_d_215_198[17:0];
      MultLoop_acc_1588_itm_1 <= nl_MultLoop_acc_1588_itm_1[17:0];
      MultLoop_acc_1578_itm_1 <= nl_MultLoop_acc_1578_itm_1[17:0];
      MultLoop_acc_1562_itm_1 <= nl_MultLoop_acc_1562_itm_1[15:0];
      MultLoop_acc_1561_itm_1 <= nl_MultLoop_acc_1561_itm_1[15:0];
      MultLoop_acc_1576_itm_1 <= nl_MultLoop_acc_1576_itm_1[16:0];
      MultLoop_acc_1575_itm_1 <= nl_MultLoop_acc_1575_itm_1[16:0];
      MultLoop_acc_1585_itm_1 <= nl_MultLoop_acc_1585_itm_1[17:0];
      MultLoop_acc_1590_itm_1 <= nl_MultLoop_acc_1590_itm_1[17:0];
      MultLoop_acc_1582_itm_1 <= nl_MultLoop_acc_1582_itm_1[17:0];
      MultLoop_acc_1581_itm_1 <= nl_MultLoop_acc_1581_itm_1[17:0];
      MultLoop_acc_3913_itm_1 <= nl_MultLoop_acc_3913_itm_1[17:0];
      MultLoop_acc_3881_itm_1 <= nl_MultLoop_acc_3881_itm_1[15:0];
      MultLoop_acc_3880_itm_1 <= nl_MultLoop_acc_3880_itm_1[15:0];
      MultLoop_acc_3896_itm_1 <= nl_MultLoop_acc_3896_itm_1[16:0];
      MultLoop_acc_3895_itm_1 <= nl_MultLoop_acc_3895_itm_1[16:0];
      MultLoop_acc_3894_itm_1 <= nl_MultLoop_acc_3894_itm_1[16:0];
      MultLoop_acc_3911_itm_1 <= nl_MultLoop_acc_3911_itm_1[17:0];
      MultLoop_acc_3910_itm_1 <= nl_MultLoop_acc_3910_itm_1[17:0];
      MultLoop_acc_1683_itm_1 <= nl_MultLoop_acc_1683_itm_1[17:0];
      MultLoop_acc_1673_itm_1 <= nl_MultLoop_acc_1673_itm_1[17:0];
      MultLoop_acc_1659_itm_1 <= nl_MultLoop_acc_1659_itm_1[15:0];
      MultLoop_acc_1658_itm_1 <= nl_MultLoop_acc_1658_itm_1[15:0];
      MultLoop_acc_1671_itm_1 <= nl_MultLoop_acc_1671_itm_1[16:0];
      MultLoop_acc_1670_itm_1 <= nl_MultLoop_acc_1670_itm_1[16:0];
      MultLoop_acc_1669_itm_1 <= nl_MultLoop_acc_1669_itm_1[16:0];
      MultLoop_acc_1668_itm_1 <= nl_MultLoop_acc_1668_itm_1[16:0];
      MultLoop_acc_1685_itm_1 <= nl_MultLoop_acc_1685_itm_1[17:0];
      MultLoop_acc_1677_itm_1 <= nl_MultLoop_acc_1677_itm_1[17:0];
      MultLoop_acc_1676_itm_1 <= nl_MultLoop_acc_1676_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1[17:0];
      MultLoop_acc_1800_itm_1 <= nl_MultLoop_acc_1800_itm_1[17:0];
      MultLoop_acc_1772_itm_1 <= nl_MultLoop_acc_1772_itm_1[15:0];
      MultLoop_acc_1771_itm_1 <= nl_MultLoop_acc_1771_itm_1[15:0];
      MultLoop_acc_1783_itm_1 <= nl_MultLoop_acc_1783_itm_1[16:0];
      MultLoop_acc_1782_itm_1 <= nl_MultLoop_acc_1782_itm_1[16:0];
      MultLoop_acc_1781_itm_1 <= nl_MultLoop_acc_1781_itm_1[16:0];
      MultLoop_acc_1780_itm_1 <= nl_MultLoop_acc_1780_itm_1[16:0];
      MultLoop_acc_1779_itm_1 <= nl_MultLoop_acc_1779_itm_1[16:0];
      MultLoop_acc_1791_itm_1 <= nl_MultLoop_acc_1791_itm_1[17:0];
      MultLoop_acc_1797_itm_1 <= nl_MultLoop_acc_1797_itm_1[17:0];
      MultLoop_acc_3720_itm_1 <= nl_MultLoop_acc_3720_itm_1[17:0];
      MultLoop_acc_3719_itm_1 <= nl_MultLoop_acc_3719_itm_1[17:0];
      MultLoop_acc_3718_itm_1 <= nl_MultLoop_acc_3718_itm_1[17:0];
      MultLoop_acc_3717_itm_1_16_0 <= nl_MultLoop_acc_3717_itm_1_16_0[16:0];
      MultLoop_acc_3716_itm_1 <= nl_MultLoop_acc_3716_itm_1[16:0];
      MultLoop_acc_3715_itm_1 <= nl_MultLoop_acc_3715_itm_1[16:0];
      MultLoop_acc_3725_itm_1 <= nl_MultLoop_acc_3725_itm_1[17:0];
      MultLoop_acc_3724_itm_1 <= nl_MultLoop_acc_3724_itm_1[17:0];
      MultLoop_acc_3710_itm_1 <= nl_MultLoop_acc_3710_itm_1[16:0];
      MultLoop_acc_3709_itm_1 <= nl_MultLoop_acc_3709_itm_1[16:0];
      MultLoop_acc_3722_itm_1 <= nl_MultLoop_acc_3722_itm_1[17:0];
      MultLoop_acc_3706_itm_1 <= nl_MultLoop_acc_3706_itm_1[16:0];
      MultLoop_acc_3705_itm_1 <= nl_MultLoop_acc_3705_itm_1[16:0];
      MultLoop_acc_1911_itm_1 <= nl_MultLoop_acc_1911_itm_1[17:0];
      MultLoop_acc_1910_itm_1 <= nl_MultLoop_acc_1910_itm_1[17:0];
      MultLoop_acc_1918_itm_1 <= nl_MultLoop_acc_1918_itm_1[17:0];
      MultLoop_acc_1917_itm_1 <= nl_MultLoop_acc_1917_itm_1[17:0];
      MultLoop_acc_1916_itm_1 <= nl_MultLoop_acc_1916_itm_1[17:0];
      MultLoop_acc_1889_itm_1 <= nl_MultLoop_acc_1889_itm_1[15:0];
      MultLoop_acc_1888_itm_1 <= nl_MultLoop_acc_1888_itm_1[15:0];
      MultLoop_acc_1902_itm_1 <= nl_MultLoop_acc_1902_itm_1[16:0];
      MultLoop_acc_1914_itm_1 <= nl_MultLoop_acc_1914_itm_1[17:0];
      MultLoop_acc_1920_itm_1 <= nl_MultLoop_acc_1920_itm_1[17:0];
      MultLoop_acc_3614_itm_1 <= nl_MultLoop_acc_3614_itm_1[17:0];
      MultLoop_acc_3598_itm_1 <= nl_MultLoop_acc_3598_itm_1[17:0];
      MultLoop_acc_3584_itm_1 <= nl_MultLoop_acc_3584_itm_1[15:0];
      MultLoop_acc_3583_itm_1 <= nl_MultLoop_acc_3583_itm_1[15:0];
      MultLoop_acc_3596_itm_1 <= nl_MultLoop_acc_3596_itm_1[16:0];
      MultLoop_acc_3595_itm_1 <= nl_MultLoop_acc_3595_itm_1[16:0];
      MultLoop_acc_3594_itm_1 <= nl_MultLoop_acc_3594_itm_1[16:0];
      MultLoop_acc_3593_itm_1 <= nl_MultLoop_acc_3593_itm_1[16:0];
      MultLoop_acc_3605_itm_1 <= nl_MultLoop_acc_3605_itm_1[17:0];
      MultLoop_acc_3611_itm_1 <= nl_MultLoop_acc_3611_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1[17:0];
      MultLoop_acc_3495_itm_1 <= nl_MultLoop_acc_3495_itm_1[17:0];
      MultLoop_acc_3494_itm_1 <= nl_MultLoop_acc_3494_itm_1[17:0];
      MultLoop_acc_3469_itm_1 <= nl_MultLoop_acc_3469_itm_1[15:0];
      MultLoop_acc_3468_itm_1 <= nl_MultLoop_acc_3468_itm_1[15:0];
      MultLoop_acc_3482_itm_1 <= nl_MultLoop_acc_3482_itm_1[16:0];
      MultLoop_acc_3481_itm_1 <= nl_MultLoop_acc_3481_itm_1[16:0];
      MultLoop_acc_3480_itm_1 <= nl_MultLoop_acc_3480_itm_1[16:0];
      MultLoop_acc_3479_itm_1 <= nl_MultLoop_acc_3479_itm_1[16:0];
      MultLoop_acc_3478_itm_1 <= nl_MultLoop_acc_3478_itm_1[16:0];
      MultLoop_acc_3490_itm_1 <= nl_MultLoop_acc_3490_itm_1[17:0];
      MultLoop_acc_3496_itm_1 <= nl_MultLoop_acc_3496_itm_1[17:0];
      MultLoop_acc_2120_itm_1 <= nl_MultLoop_acc_2120_itm_1[17:0];
      MultLoop_acc_2119_itm_1 <= nl_MultLoop_acc_2119_itm_1[17:0];
      MultLoop_acc_2118_itm_1 <= nl_MultLoop_acc_2118_itm_1[17:0];
      MultLoop_acc_2091_itm_1 <= nl_MultLoop_acc_2091_itm_1[15:0];
      MultLoop_acc_2090_itm_1 <= nl_MultLoop_acc_2090_itm_1[15:0];
      MultLoop_acc_2105_itm_1 <= nl_MultLoop_acc_2105_itm_1[16:0];
      MultLoop_acc_2104_itm_1 <= nl_MultLoop_acc_2104_itm_1[16:0];
      MultLoop_acc_2103_itm_1 <= nl_MultLoop_acc_2103_itm_1[16:0];
      MultLoop_acc_2115_itm_1 <= nl_MultLoop_acc_2115_itm_1[17:0];
      MultLoop_acc_2121_itm_1 <= nl_MultLoop_acc_2121_itm_1[17:0];
      MultLoop_acc_3378_itm_1 <= nl_MultLoop_acc_3378_itm_1[17:0];
      MultLoop_acc_3368_itm_1 <= nl_MultLoop_acc_3368_itm_1[17:0];
      MultLoop_acc_3367_itm_1 <= nl_MultLoop_acc_3367_itm_1[16:0];
      MultLoop_acc_3366_itm_1 <= nl_MultLoop_acc_3366_itm_1[16:0];
      MultLoop_acc_3365_itm_1 <= nl_MultLoop_acc_3365_itm_1[16:0];
      MultLoop_acc_3375_itm_1 <= nl_MultLoop_acc_3375_itm_1[17:0];
      MultLoop_acc_3362_itm_1 <= nl_MultLoop_acc_3362_itm_1[16:0];
      MultLoop_acc_3361_itm_1 <= nl_MultLoop_acc_3361_itm_1[16:0];
      MultLoop_acc_3373_itm_1 <= nl_MultLoop_acc_3373_itm_1[17:0];
      MultLoop_acc_3379_itm_1 <= nl_MultLoop_acc_3379_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_23_7_itm_1
          <= readslicef_24_17_7((MultLoop_acc_815_nl));
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1[17:0];
      MultLoop_acc_3264_itm_1 <= nl_MultLoop_acc_3264_itm_1[17:0];
      MultLoop_acc_3258_itm_1 <= nl_MultLoop_acc_3258_itm_1[17:0];
      MultLoop_acc_3233_itm_1 <= nl_MultLoop_acc_3233_itm_1[15:0];
      MultLoop_acc_3232_itm_1 <= nl_MultLoop_acc_3232_itm_1[15:0];
      MultLoop_acc_3245_itm_1 <= nl_MultLoop_acc_3245_itm_1[16:0];
      MultLoop_acc_3256_itm_1 <= nl_MultLoop_acc_3256_itm_1[17:0];
      MultLoop_acc_3255_itm_1 <= nl_MultLoop_acc_3255_itm_1[17:0];
      MultLoop_acc_3254_itm_1 <= nl_MultLoop_acc_3254_itm_1[17:0];
      MultLoop_acc_3238_itm_1 <= nl_MultLoop_acc_3238_itm_1[16:0];
      MultLoop_acc_3237_itm_1 <= nl_MultLoop_acc_3237_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0 <=
          nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_26_10_itm_1
          <= readslicef_27_17_10((MultLoop_acc_720_nl));
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_acc_1215_22_6_itm_1
          <= readslicef_23_17_6((MultLoop_acc_1215_nl));
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1[14:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1[14:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1[17:0];
      MultLoop_acc_2470_itm_1 <= nl_MultLoop_acc_2470_itm_1[17:0];
      MultLoop_acc_2469_itm_1 <= nl_MultLoop_acc_2469_itm_1[17:0];
      MultLoop_acc_2458_itm_1 <= nl_MultLoop_acc_2458_itm_1[16:0];
      MultLoop_acc_2457_itm_1 <= nl_MultLoop_acc_2457_itm_1[16:0];
      MultLoop_acc_2438_itm_1 <= nl_MultLoop_acc_2438_itm_1[15:0];
      MultLoop_acc_2437_itm_1 <= nl_MultLoop_acc_2437_itm_1[15:0];
      MultLoop_acc_2455_itm_1 <= nl_MultLoop_acc_2455_itm_1[16:0];
      MultLoop_acc_2466_itm_1 <= nl_MultLoop_acc_2466_itm_1[17:0];
      MultLoop_acc_2452_itm_1 <= nl_MultLoop_acc_2452_itm_1[16:0];
      MultLoop_acc_2451_itm_1 <= nl_MultLoop_acc_2451_itm_1[16:0];
      MultLoop_acc_2464_itm_1 <= nl_MultLoop_acc_2464_itm_1[17:0];
      MultLoop_acc_2463_itm_1 <= nl_MultLoop_acc_2463_itm_1[17:0];
      MultLoop_acc_3018_itm_1 <= nl_MultLoop_acc_3018_itm_1[17:0];
      MultLoop_acc_3008_itm_1 <= nl_MultLoop_acc_3008_itm_1[17:0];
      MultLoop_acc_2984_itm_1 <= nl_MultLoop_acc_2984_itm_1[14:0];
      MultLoop_acc_2983_itm_1 <= nl_MultLoop_acc_2983_itm_1[14:0];
      MultLoop_acc_2993_itm_1 <= nl_MultLoop_acc_2993_itm_1[15:0];
      MultLoop_acc_3006_itm_1 <= nl_MultLoop_acc_3006_itm_1[16:0];
      MultLoop_acc_3005_itm_1 <= nl_MultLoop_acc_3005_itm_1[16:0];
      MultLoop_acc_3004_itm_1 <= nl_MultLoop_acc_3004_itm_1[16:0];
      MultLoop_acc_3003_itm_1 <= nl_MultLoop_acc_3003_itm_1[16:0];
      MultLoop_acc_3020_itm_1 <= nl_MultLoop_acc_3020_itm_1[17:0];
      MultLoop_acc_3012_itm_1 <= nl_MultLoop_acc_3012_itm_1[17:0];
      MultLoop_acc_3011_itm_1 <= nl_MultLoop_acc_3011_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0 <=
          nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1[15:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_25_10_itm_1
          <= readslicef_18_16_2((MultLoop_acc_4207_nl));
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1[16:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1[17:0];
      nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1 <= nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1[17:0];
      MultLoop_acc_2888_itm_1 <= nl_MultLoop_acc_2888_itm_1[17:0];
      MultLoop_acc_2887_itm_1 <= nl_MultLoop_acc_2887_itm_1[17:0];
      MultLoop_acc_2886_itm_1 <= nl_MultLoop_acc_2886_itm_1[17:0];
      MultLoop_acc_2871_itm_1 <= nl_MultLoop_acc_2871_itm_1[15:0];
      MultLoop_acc_2870_itm_1 <= nl_MultLoop_acc_2870_itm_1[15:0];
      MultLoop_acc_2884_itm_1 <= nl_MultLoop_acc_2884_itm_1[16:0];
      MultLoop_acc_2883_itm_1 <= nl_MultLoop_acc_2883_itm_1[16:0];
      MultLoop_acc_2893_itm_1 <= nl_MultLoop_acc_2893_itm_1[17:0];
      MultLoop_acc_2898_itm_1 <= nl_MultLoop_acc_2898_itm_1[17:0];
      MultLoop_acc_2897_itm_1 <= nl_MultLoop_acc_2897_itm_1[17:0];
      MultLoop_acc_2658_itm_1 <= nl_MultLoop_acc_2658_itm_1[17:0];
      MultLoop_acc_2657_itm_1 <= nl_MultLoop_acc_2657_itm_1[17:0];
      MultLoop_acc_2656_itm_1 <= nl_MultLoop_acc_2656_itm_1[17:0];
      MultLoop_acc_2631_itm_1 <= nl_MultLoop_acc_2631_itm_1[15:0];
      MultLoop_acc_2630_itm_1 <= nl_MultLoop_acc_2630_itm_1[15:0];
      MultLoop_acc_2643_itm_1 <= nl_MultLoop_acc_2643_itm_1[16:0];
      MultLoop_acc_2642_itm_1 <= nl_MultLoop_acc_2642_itm_1[16:0];
      MultLoop_acc_2641_itm_1 <= nl_MultLoop_acc_2641_itm_1[16:0];
      MultLoop_acc_2653_itm_1 <= nl_MultLoop_acc_2653_itm_1[17:0];
      MultLoop_acc_2659_itm_1 <= nl_MultLoop_acc_2659_itm_1[17:0];
      MultLoop_acc_2773_itm_1 <= nl_MultLoop_acc_2773_itm_1[17:0];
      MultLoop_acc_2750_itm_1 <= nl_MultLoop_acc_2750_itm_1[15:0];
      MultLoop_acc_2749_itm_1 <= nl_MultLoop_acc_2749_itm_1[15:0];
      MultLoop_acc_2748_itm_1 <= nl_MultLoop_acc_2748_itm_1[15:0];
      MultLoop_acc_2747_itm_1 <= nl_MultLoop_acc_2747_itm_1[15:0];
      MultLoop_acc_2761_itm_1 <= nl_MultLoop_acc_2761_itm_1[16:0];
      MultLoop_acc_2760_itm_1 <= nl_MultLoop_acc_2760_itm_1[16:0];
      MultLoop_acc_2770_itm_1 <= nl_MultLoop_acc_2770_itm_1[17:0];
      MultLoop_acc_2775_itm_1 <= nl_MultLoop_acc_2775_itm_1[17:0];
      MultLoop_acc_2774_itm_1 <= nl_MultLoop_acc_2774_itm_1[17:0];
    end
  end
  assign nl_MultLoop_acc_1591_nl = MultLoop_acc_1585_itm_1 + conv_s2s_17_18(MultLoop_acc_1576_itm_1)
      + conv_s2s_17_18(MultLoop_acc_1575_itm_1);
  assign MultLoop_acc_1591_nl = nl_MultLoop_acc_1591_nl[17:0];
  assign nl_MultLoop_acc_1587_nl = MultLoop_acc_1578_itm_1 + conv_s2s_16_18(MultLoop_acc_1562_itm_1)
      + conv_s2s_16_18(MultLoop_acc_1561_itm_1);
  assign MultLoop_acc_1587_nl = nl_MultLoop_acc_1587_nl[17:0];
  assign nl_res_rsci_d_431_414  = (MultLoop_acc_1591_nl) + MultLoop_acc_1590_itm_1
      + MultLoop_acc_1582_itm_1 + MultLoop_acc_1581_itm_1 + MultLoop_acc_1588_itm_1
      + (MultLoop_acc_1587_nl);
  assign nl_MultLoop_acc_3912_nl = conv_s2s_17_18(MultLoop_acc_3896_itm_1) + conv_s2s_17_18(MultLoop_acc_3895_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3894_itm_1) + conv_s2s_16_18(MultLoop_acc_3881_itm_1)
      + conv_s2s_16_18(MultLoop_acc_3880_itm_1);
  assign MultLoop_acc_3912_nl = nl_MultLoop_acc_3912_nl[17:0];
  assign nl_res_rsci_d_17_0  = MultLoop_acc_3913_itm_1 + (MultLoop_acc_3912_nl) +
      MultLoop_acc_3911_itm_1 + MultLoop_acc_3910_itm_1;
  assign nl_MultLoop_acc_1686_nl = conv_s2s_17_18(MultLoop_acc_1671_itm_1) + conv_s2s_17_18(MultLoop_acc_1670_itm_1)
      + conv_s2s_17_18(MultLoop_acc_1669_itm_1) + conv_s2s_17_18(MultLoop_acc_1668_itm_1);
  assign MultLoop_acc_1686_nl = nl_MultLoop_acc_1686_nl[17:0];
  assign nl_MultLoop_acc_1682_nl = MultLoop_acc_1673_itm_1 + conv_s2s_16_18(MultLoop_acc_1659_itm_1)
      + conv_s2s_16_18(MultLoop_acc_1658_itm_1);
  assign MultLoop_acc_1682_nl = nl_MultLoop_acc_1682_nl[17:0];
  assign nl_res_rsci_d_413_396  = (MultLoop_acc_1686_nl) + MultLoop_acc_1685_itm_1
      + MultLoop_acc_1677_itm_1 + MultLoop_acc_1676_itm_1 + MultLoop_acc_1683_itm_1
      + (MultLoop_acc_1682_nl);
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl[17:0];
  assign nl_res_rsci_d_35_18  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_370_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_369_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1;
  assign nl_MultLoop_acc_1799_nl = conv_s2s_17_18(MultLoop_acc_1783_itm_1) + conv_s2s_17_18(MultLoop_acc_1782_itm_1)
      + conv_s2s_17_18(MultLoop_acc_1781_itm_1) + conv_s2s_16_18(MultLoop_acc_1772_itm_1)
      + conv_s2s_16_18(MultLoop_acc_1771_itm_1);
  assign MultLoop_acc_1799_nl = nl_MultLoop_acc_1799_nl[17:0];
  assign nl_res_rsci_d_395_378  = MultLoop_acc_1800_itm_1 + (MultLoop_acc_1799_nl)
      + MultLoop_acc_1797_itm_1 + MultLoop_acc_1791_itm_1 + conv_s2s_17_18(MultLoop_acc_1780_itm_1)
      + conv_s2s_17_18(MultLoop_acc_1779_itm_1);
  assign nl_MultLoop_acc_3731_nl = MultLoop_acc_3725_itm_1 + conv_s2s_17_18(MultLoop_acc_3716_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3715_itm_1);
  assign MultLoop_acc_3731_nl = nl_MultLoop_acc_3731_nl[17:0];
  assign nl_MultLoop_acc_3729_nl = MultLoop_acc_3722_itm_1 + conv_s2s_17_18(MultLoop_acc_3706_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3705_itm_1);
  assign MultLoop_acc_3729_nl = nl_MultLoop_acc_3729_nl[17:0];
  assign nl_MultLoop_acc_3727_nl = MultLoop_acc_3718_itm_1 + conv_s2s_17_18(MultLoop_acc_3717_itm_1_16_0);
  assign MultLoop_acc_3727_nl = nl_MultLoop_acc_3727_nl[17:0];
  assign nl_res_rsci_d_53_36  = (MultLoop_acc_3731_nl) + (MultLoop_acc_3729_nl) +
      MultLoop_acc_3724_itm_1 + (MultLoop_acc_3727_nl) + MultLoop_acc_3720_itm_1
      + MultLoop_acc_3719_itm_1 + conv_s2s_17_18(MultLoop_acc_3710_itm_1) + conv_s2s_17_18(MultLoop_acc_3709_itm_1);
  assign nl_res_rsci_d_377_360  = MultLoop_acc_1920_itm_1 + MultLoop_acc_1914_itm_1
      + MultLoop_acc_1918_itm_1 + MultLoop_acc_1911_itm_1 + MultLoop_acc_1910_itm_1
      + MultLoop_acc_1917_itm_1 + MultLoop_acc_1916_itm_1 + conv_s2s_17_18(MultLoop_acc_1902_itm_1)
      + conv_s2s_16_18(MultLoop_acc_1889_itm_1) + conv_s2s_16_18(MultLoop_acc_1888_itm_1);
  assign nl_MultLoop_acc_3608_nl = MultLoop_acc_3598_itm_1 + conv_s2s_16_18(MultLoop_acc_3584_itm_1)
      + conv_s2s_16_18(MultLoop_acc_3583_itm_1);
  assign MultLoop_acc_3608_nl = nl_MultLoop_acc_3608_nl[17:0];
  assign nl_MultLoop_acc_3613_nl = (MultLoop_acc_3608_nl) + conv_s2s_17_18(MultLoop_acc_3596_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3595_itm_1);
  assign MultLoop_acc_3613_nl = nl_MultLoop_acc_3613_nl[17:0];
  assign nl_res_rsci_d_71_54  = MultLoop_acc_3614_itm_1 + (MultLoop_acc_3613_nl)
      + MultLoop_acc_3611_itm_1 + MultLoop_acc_3605_itm_1 + conv_s2s_17_18(MultLoop_acc_3594_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3593_itm_1);
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl[17:0];
  assign nl_res_rsci_d_359_342  = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1 + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_48_nl)
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1 + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1);
  assign nl_MultLoop_acc_3498_nl = conv_s2s_17_18(MultLoop_acc_3482_itm_1) + conv_s2s_17_18(MultLoop_acc_3481_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3480_itm_1) + conv_s2s_16_18(MultLoop_acc_3469_itm_1)
      + conv_s2s_16_18(MultLoop_acc_3468_itm_1);
  assign MultLoop_acc_3498_nl = nl_MultLoop_acc_3498_nl[17:0];
  assign nl_res_rsci_d_89_72  = (MultLoop_acc_3498_nl) + MultLoop_acc_3496_itm_1
      + MultLoop_acc_3490_itm_1 + MultLoop_acc_3495_itm_1 + MultLoop_acc_3494_itm_1
      + conv_s2s_17_18(MultLoop_acc_3479_itm_1) + conv_s2s_17_18(MultLoop_acc_3478_itm_1);
  assign nl_MultLoop_acc_2123_nl = MultLoop_acc_2118_itm_1 + conv_s2s_17_18(MultLoop_acc_2105_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2091_itm_1) + conv_s2s_16_18(MultLoop_acc_2090_itm_1);
  assign MultLoop_acc_2123_nl = nl_MultLoop_acc_2123_nl[17:0];
  assign nl_res_rsci_d_341_324  = (MultLoop_acc_2123_nl) + MultLoop_acc_2121_itm_1
      + MultLoop_acc_2115_itm_1 + MultLoop_acc_2120_itm_1 + MultLoop_acc_2119_itm_1
      + conv_s2s_17_18(MultLoop_acc_2104_itm_1) + conv_s2s_17_18(MultLoop_acc_2103_itm_1);
  assign nl_MultLoop_acc_3381_nl = MultLoop_acc_3375_itm_1 + conv_s2s_17_18(MultLoop_acc_3366_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3365_itm_1);
  assign MultLoop_acc_3381_nl = nl_MultLoop_acc_3381_nl[17:0];
  assign nl_MultLoop_acc_3377_nl = MultLoop_acc_3368_itm_1 + conv_s2s_17_18(MultLoop_acc_3367_itm_1);
  assign MultLoop_acc_3377_nl = nl_MultLoop_acc_3377_nl[17:0];
  assign nl_res_rsci_d_107_90  = (MultLoop_acc_3381_nl) + MultLoop_acc_3379_itm_1
      + MultLoop_acc_3373_itm_1 + MultLoop_acc_3378_itm_1 + (MultLoop_acc_3377_nl)
      + conv_s2s_17_18(MultLoop_acc_3362_itm_1) + conv_s2s_17_18(MultLoop_acc_3361_itm_1);
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl = conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_825_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_23_7_itm_1
      + conv_s2s_16_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_85_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl[17:0];
  assign nl_res_rsci_d_323_306  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_99_nl)
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1 + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_95_nl);
  assign nl_MultLoop_acc_3263_nl = MultLoop_acc_3258_itm_1 + conv_s2s_17_18(MultLoop_acc_3245_itm_1)
      + conv_s2s_16_18(MultLoop_acc_3233_itm_1) + conv_s2s_16_18(MultLoop_acc_3232_itm_1);
  assign MultLoop_acc_3263_nl = nl_MultLoop_acc_3263_nl[17:0];
  assign nl_MultLoop_acc_3261_nl = MultLoop_acc_3254_itm_1 + conv_s2s_17_18(MultLoop_acc_3238_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3237_itm_1);
  assign MultLoop_acc_3261_nl = nl_MultLoop_acc_3261_nl[17:0];
  assign nl_res_rsci_d_125_108  = MultLoop_acc_3264_itm_1 + (MultLoop_acc_3263_nl)
      + (MultLoop_acc_3261_nl) + MultLoop_acc_3256_itm_1 + MultLoop_acc_3255_itm_1;
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_139_nl)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl = conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl[17:0];
  assign nl_res_rsci_d_305_288  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_143_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_142_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1;
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl = conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl[17:0];
  assign nl_res_rsci_d_143_126  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_324_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_323_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1);
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_728_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_26_10_itm_1
      + conv_s2s_16_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_174_nl)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl[17:0];
  assign nl_res_rsci_d_287_270  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_188_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_187_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1;
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_acc_1215_22_6_itm_1
      + conv_s2s_15_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1)
      + conv_s2s_15_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl = conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_265_nl)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl[17:0];
  assign nl_res_rsci_d_161_144  = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_280_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1 + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1);
  assign nl_MultLoop_acc_2473_nl = conv_s2s_17_18(MultLoop_acc_2458_itm_1) + conv_s2s_17_18(MultLoop_acc_2457_itm_1)
      + conv_s2s_17_18(MultLoop_acc_2455_itm_1) + conv_s2s_16_18(MultLoop_acc_2438_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2437_itm_1);
  assign MultLoop_acc_2473_nl = nl_MultLoop_acc_2473_nl[17:0];
  assign nl_res_rsci_d_269_252  = (MultLoop_acc_2473_nl) + MultLoop_acc_2466_itm_1
      + MultLoop_acc_2470_itm_1 + MultLoop_acc_2469_itm_1 + MultLoop_acc_2464_itm_1
      + MultLoop_acc_2463_itm_1 + conv_s2s_17_18(MultLoop_acc_2452_itm_1) + conv_s2s_17_18(MultLoop_acc_2451_itm_1);
  assign nl_MultLoop_acc_3021_nl = conv_s2s_17_18(MultLoop_acc_3006_itm_1) + conv_s2s_17_18(MultLoop_acc_3005_itm_1)
      + conv_s2s_17_18(MultLoop_acc_3004_itm_1) + conv_s2s_17_18(MultLoop_acc_3003_itm_1);
  assign MultLoop_acc_3021_nl = nl_MultLoop_acc_3021_nl[17:0];
  assign nl_MultLoop_acc_3017_nl = MultLoop_acc_3008_itm_1 + conv_s2s_16_18(MultLoop_acc_2993_itm_1)
      + conv_s2s_15_18(MultLoop_acc_2984_itm_1) + conv_s2s_15_18(MultLoop_acc_2983_itm_1);
  assign MultLoop_acc_3017_nl = nl_MultLoop_acc_3017_nl[17:0];
  assign nl_res_rsci_d_179_162  = (MultLoop_acc_3021_nl) + MultLoop_acc_3020_itm_1
      + MultLoop_acc_3012_itm_1 + MultLoop_acc_3011_itm_1 + MultLoop_acc_3018_itm_1
      + (MultLoop_acc_3017_nl);
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl = nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_230_nl)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl = conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1)
      + conv_s2s_17_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1)
      + conv_s2s_16_18(nnet_product_input_t_config2_weight_t_config2_accum_t_slc_MultLoop_667_nnet_product_input_t_config2_weight_t_config2_accum_t_mul_25_10_itm_1);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl[17:0];
  assign nl_res_rsci_d_251_234  = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_234_nl)
      + (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_233_nl) + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1
      + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1 + nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1;
  assign nl_MultLoop_acc_2899_nl = MultLoop_acc_2893_itm_1 + conv_s2s_17_18(MultLoop_acc_2884_itm_1)
      + conv_s2s_17_18(MultLoop_acc_2883_itm_1);
  assign MultLoop_acc_2899_nl = nl_MultLoop_acc_2899_nl[17:0];
  assign nl_MultLoop_acc_2895_nl = MultLoop_acc_2886_itm_1 + conv_s2s_16_18(MultLoop_acc_2871_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2870_itm_1);
  assign MultLoop_acc_2895_nl = nl_MultLoop_acc_2895_nl[17:0];
  assign nl_res_rsci_d_197_180  = (MultLoop_acc_2899_nl) + MultLoop_acc_2898_itm_1
      + MultLoop_acc_2897_itm_1 + (MultLoop_acc_2895_nl) + MultLoop_acc_2888_itm_1
      + MultLoop_acc_2887_itm_1;
  assign nl_MultLoop_acc_2661_nl = MultLoop_acc_2656_itm_1 + conv_s2s_17_18(MultLoop_acc_2643_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2631_itm_1) + conv_s2s_16_18(MultLoop_acc_2630_itm_1);
  assign MultLoop_acc_2661_nl = nl_MultLoop_acc_2661_nl[17:0];
  assign nl_res_rsci_d_233_216  = (MultLoop_acc_2661_nl) + MultLoop_acc_2659_itm_1
      + MultLoop_acc_2653_itm_1 + MultLoop_acc_2658_itm_1 + MultLoop_acc_2657_itm_1
      + conv_s2s_17_18(MultLoop_acc_2642_itm_1) + conv_s2s_17_18(MultLoop_acc_2641_itm_1);
  assign nl_MultLoop_acc_2777_nl = MultLoop_acc_2773_itm_1 + conv_s2s_16_18(MultLoop_acc_2750_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2749_itm_1) + conv_s2s_16_18(MultLoop_acc_2748_itm_1)
      + conv_s2s_16_18(MultLoop_acc_2747_itm_1);
  assign MultLoop_acc_2777_nl = nl_MultLoop_acc_2777_nl[17:0];
  assign nl_MultLoop_acc_2776_nl = MultLoop_acc_2770_itm_1 + conv_s2s_17_18(MultLoop_acc_2761_itm_1)
      + conv_s2s_17_18(MultLoop_acc_2760_itm_1);
  assign MultLoop_acc_2776_nl = nl_MultLoop_acc_2776_nl[17:0];
  assign nl_res_rsci_d_215_198  = (MultLoop_acc_2777_nl) + (MultLoop_acc_2776_nl)
      + MultLoop_acc_2775_itm_1 + MultLoop_acc_2774_itm_1;
  assign nl_Result_acc_17_nl = conv_s2s_19_27({MultLoop_MultLoop_conc_780_18_8 ,
      (~ (data_rsci_idat[25:18]))}) + conv_s2s_26_27({(~ (data_rsci_idat[35:18]))
      , 8'b00000001});
  assign Result_acc_17_nl = nl_Result_acc_17_nl[26:0];
  assign nl_Result_acc_181_nl = conv_s2s_10_11(data_rsci_idat[71:62]) + 11'b00000000001;
  assign Result_acc_181_nl = nl_Result_acc_181_nl[10:0];
  assign nl_Result_acc_146_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_17_18({(Result_acc_181_nl)
      , (data_rsci_idat[61:56])});
  assign Result_acc_146_nl = nl_Result_acc_146_nl[17:0];
  assign nl_Result_acc_77_nl = conv_s2u_18_25(Result_acc_146_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[71:54])) , 6'b000001});
  assign Result_acc_77_nl = nl_Result_acc_77_nl[24:0];
  assign nl_Result_acc_142_nl = conv_s2s_18_19(data_rsci_idat[827:810]) + conv_s2s_15_19({Result_acc_178_cse_1
      , (data_rsci_idat[817:814])});
  assign Result_acc_142_nl = nl_Result_acc_142_nl[18:0];
  assign nl_Result_acc_59_nl = conv_s2u_19_22(Result_acc_142_nl) + ({(~ (data_rsci_idat[827:810]))
      , 4'b0000});
  assign Result_acc_59_nl = nl_Result_acc_59_nl[21:0];
  assign nl_Result_acc_75_nl = conv_s2u_18_22(Result_acc_143_cse_1) + ({(data_rsci_idat[845:828])
      , 4'b0001});
  assign Result_acc_75_nl = nl_Result_acc_75_nl[21:0];
  assign nl_Result_acc_23_nl = conv_s2s_18_22(~ (data_rsci_idat[143:126])) + ({(data_rsci_idat[143:126])
      , 4'b0001});
  assign Result_acc_23_nl = nl_Result_acc_23_nl[21:0];
  assign nl_Result_acc_179_nl =  -conv_s2s_15_16(data_rsci_idat[755:741]);
  assign Result_acc_179_nl = nl_Result_acc_179_nl[15:0];
  assign nl_Result_acc_55_nl = conv_s2s_19_22({(Result_acc_179_nl) , (~ (data_rsci_idat[740:738]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[755:738])) , 3'b001});
  assign Result_acc_55_nl = nl_Result_acc_55_nl[21:0];
  assign nl_Result_acc_57_nl = conv_s2s_18_21(~ (data_rsci_idat[791:774])) + ({(data_rsci_idat[791:774])
      , 3'b001});
  assign Result_acc_57_nl = nl_Result_acc_57_nl[20:0];
  assign nl_MultLoop_acc_1588_itm_1  = conv_s2s_17_18(readslicef_27_17_10((Result_acc_17_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((Result_acc_77_nl))) + conv_s2s_16_18(readslicef_22_16_6((Result_acc_59_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((Result_acc_75_nl))) + conv_s2s_16_18(MultLoop_acc_1315_itm_19_4)
      + conv_s2s_14_18(readslicef_22_14_8((Result_acc_23_nl))) + conv_s2s_13_18(readslicef_22_13_9((Result_acc_55_nl)))
      + conv_s2s_13_18(readslicef_21_13_8((Result_acc_57_nl)));
  assign nl_Result_acc_149_nl = ({(~ (data_rsci_idat[395:378])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[395:378])
      + conv_s2s_17_20({MultLoop_MultLoop_conc_790_16_4 , (data_rsci_idat[383:380])});
  assign Result_acc_149_nl = nl_Result_acc_149_nl[19:0];
  assign nl_Result_acc_78_nl = conv_s2u_20_23(Result_acc_149_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[395:378])) , 4'b0100});
  assign Result_acc_78_nl = nl_Result_acc_78_nl[22:0];
  assign nl_Result_acc_151_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_16_18({Result_acc_183_cse_1
      , (data_rsci_idat[690:687])});
  assign Result_acc_151_nl = nl_Result_acc_151_nl[17:0];
  assign nl_Result_acc_79_nl = conv_s2u_18_23(Result_acc_151_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[701:684])) , 4'b0001});
  assign Result_acc_79_nl = nl_Result_acc_79_nl[22:0];
  assign nl_MultLoop_acc_1578_itm_1  = conv_s2s_17_18(readslicef_23_17_6((Result_acc_78_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((Result_acc_79_nl)));
  assign nl_Result_acc_184_nl =  -conv_s2s_13_14(data_rsci_idat[251:239]);
  assign Result_acc_184_nl = nl_Result_acc_184_nl[13:0];
  assign nl_Result_acc_29_nl = conv_s2s_23_24({(~ (data_rsci_idat[251:234])) , 5'b01000})
      + conv_s2s_21_24({(~ (data_rsci_idat[251:234])) , 3'b001}) + conv_s2s_19_24({(Result_acc_184_nl)
      , (~ (data_rsci_idat[238:234]))});
  assign Result_acc_29_nl = nl_Result_acc_29_nl[23:0];
  assign nl_Result_acc_63_nl = conv_s2u_15_19(data_rsci_idat[323:309]) + conv_s2u_18_19(data_rsci_idat[323:306]);
  assign Result_acc_63_nl = nl_Result_acc_63_nl[18:0];
  assign nl_Result_acc_217_nl = conv_s2u_19_20(MultLoop_acc_1520_cse_1[20:2]) + ({(data_rsci_idat[359:342])
      , 2'b01});
  assign Result_acc_217_nl = nl_Result_acc_217_nl[19:0];
  assign nl_Result_acc_88_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_15_18(data_rsci_idat[377:363]);
  assign Result_acc_88_nl = nl_Result_acc_88_nl[17:0];
  assign nl_Result_acc_64_nl = conv_s2u_18_21(Result_acc_88_nl) + ({(data_rsci_idat[377:360])
      , 3'b001});
  assign Result_acc_64_nl = nl_Result_acc_64_nl[20:0];
  assign nl_MultLoop_acc_1562_itm_1  = conv_s2s_14_16(readslicef_24_14_10((Result_acc_29_nl)))
      + conv_s2s_14_16(readslicef_19_14_5((Result_acc_63_nl))) + conv_s2s_14_16(readslicef_20_14_6((Result_acc_217_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((Result_acc_64_nl)));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl = ({(data_rsci_idat[17:0])
      , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_708_18_6 , (~ (data_rsci_idat[5:0]))});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = conv_s2u_15_18(readslicef_21_15_6((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_11_nl)))
      + (~ (data_rsci_idat[17:0]));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl[17:0];
  assign nl_Result_acc_89_nl = conv_s2s_21_22({(~ (data_rsci_idat[431:414])) , 3'b001})
      + conv_s2s_18_22(~ (data_rsci_idat[431:414]));
  assign Result_acc_89_nl = nl_Result_acc_89_nl[21:0];
  assign nl_Result_acc_38_nl = conv_s2s_22_24(Result_acc_89_nl) + ({(data_rsci_idat[431:414])
      , 6'b001000});
  assign Result_acc_38_nl = nl_Result_acc_38_nl[23:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_9_nl = ~((data_rsci_idat[271:270]!=2'b00));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_10_nl = ~((data_rsci_idat[437:432]!=6'b000000));
  assign nl_MultLoop_acc_1548_nl = conv_s2s_12_13(~ (data_rsci_idat[449:438])) +
      conv_u2s_9_13({8'b10100101 , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_9_nl)})
      + conv_u2s_1_13(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_10_nl);
  assign MultLoop_acc_1548_nl = nl_MultLoop_acc_1548_nl[12:0];
  assign nl_MultLoop_acc_1561_itm_1  = conv_s2s_15_16(readslicef_18_15_3((nnet_product_input_t_config2_weight_t_config2_accum_t_acc_nl)))
      + conv_s2s_14_16(readslicef_24_14_10((Result_acc_38_nl))) + conv_s2s_13_16(MultLoop_acc_1548_nl);
  assign nl_Result_acc_185_nl =  -conv_s2s_11_12(data_rsci_idat[53:43]);
  assign Result_acc_185_nl = nl_Result_acc_185_nl[11:0];
  assign nl_Result_acc_92_nl = ({(data_rsci_idat[53:36]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[53:36])) , 3'b001}) + conv_s2s_19_23({(Result_acc_185_nl) ,
      (~ (data_rsci_idat[42:36]))});
  assign Result_acc_92_nl = nl_Result_acc_92_nl[22:0];
  assign nl_Result_acc_186_nl = conv_s2u_16_18(readslicef_23_16_7((Result_acc_92_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign Result_acc_186_nl = nl_Result_acc_186_nl[17:0];
  assign nl_Result_acc_93_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_16_18(data_rsci_idat[89:74]);
  assign Result_acc_93_nl = nl_Result_acc_93_nl[17:0];
  assign nl_Result_acc_65_nl = conv_s2u_18_20(Result_acc_93_nl) + ({(data_rsci_idat[89:72])
      , 2'b01});
  assign Result_acc_65_nl = nl_Result_acc_65_nl[19:0];
  assign nl_Result_acc_96_nl = conv_s2s_20_21({(data_rsci_idat[125:108]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[125:108]) + conv_s2s_16_21({Result_acc_187_cse_1
      , (data_rsci_idat[114:111])});
  assign Result_acc_96_nl = nl_Result_acc_96_nl[20:0];
  assign nl_Result_acc_22_nl = conv_s2u_21_22(Result_acc_96_nl) + ({(~ (data_rsci_idat[125:108]))
      , 4'b0000});
  assign Result_acc_22_nl = nl_Result_acc_22_nl[21:0];
  assign nl_Result_acc_99_nl = ({(data_rsci_idat[233:216]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[233:216])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_730_18_7
      , (~ (data_rsci_idat[222:216]))});
  assign Result_acc_99_nl = nl_Result_acc_99_nl[21:0];
  assign nl_Result_acc_189_nl = conv_s2u_15_18(readslicef_22_15_7((Result_acc_99_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign Result_acc_189_nl = nl_Result_acc_189_nl[17:0];
  assign nl_MultLoop_acc_1576_itm_1  = conv_s2s_15_17(readslicef_18_15_3((Result_acc_186_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((Result_acc_65_nl))) + conv_s2s_15_17(readslicef_22_15_7((Result_acc_22_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((Result_acc_189_nl)));
  assign nl_Result_acc_101_nl = (~ (data_rsci_idat[503:486])) + conv_s2s_15_18({Result_acc_190_cse_1
      , (data_rsci_idat[491:490])});
  assign Result_acc_101_nl = nl_Result_acc_101_nl[17:0];
  assign nl_Result_acc_66_nl = conv_s2u_18_21(Result_acc_101_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[503:486])) , 2'b01});
  assign Result_acc_66_nl = nl_Result_acc_66_nl[20:0];
  assign nl_Result_acc_219_nl = conv_s2u_19_21(Result_acc_102_itm_20_2_1) + ({(data_rsci_idat[521:504])
      , 3'b001});
  assign Result_acc_219_nl = nl_Result_acc_219_nl[20:0];
  assign nl_Result_acc_103_nl = conv_s2s_18_19(data_rsci_idat[557:540]) + conv_s2s_16_19(data_rsci_idat[557:542]);
  assign Result_acc_103_nl = nl_Result_acc_103_nl[18:0];
  assign nl_Result_acc_67_nl = conv_s2u_19_23(Result_acc_103_nl) + conv_s2u_22_23({(data_rsci_idat[557:540])
      , 4'b0000});
  assign Result_acc_67_nl = nl_Result_acc_67_nl[22:0];
  assign nl_Result_acc_104_nl = (~ (data_rsci_idat[647:630])) + conv_s2s_15_18(data_rsci_idat[647:633]);
  assign Result_acc_104_nl = nl_Result_acc_104_nl[17:0];
  assign nl_Result_acc_68_nl = conv_s2u_18_22(Result_acc_104_nl) + ({(data_rsci_idat[647:630])
      , 4'b0001});
  assign Result_acc_68_nl = nl_Result_acc_68_nl[21:0];
  assign nl_MultLoop_acc_1575_itm_1  = conv_s2s_15_17(readslicef_21_15_6((Result_acc_66_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((Result_acc_219_nl))) + conv_s2s_15_17(readslicef_23_15_8((Result_acc_67_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((Result_acc_68_nl)));
  assign nl_Result_acc_112_nl = ({(~ (data_rsci_idat[107:90])) , 4'b0000}) + conv_s2s_19_22(Result_acc_111_cse_1);
  assign Result_acc_112_nl = nl_Result_acc_112_nl[21:0];
  assign nl_Result_acc_70_nl = conv_s2u_22_24(Result_acc_112_nl) + ({(data_rsci_idat[107:90])
      , 6'b010000});
  assign Result_acc_70_nl = nl_Result_acc_70_nl[23:0];
  assign nl_Result_acc_114_nl = conv_s2s_20_21({(data_rsci_idat[161:144]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[161:144]) + conv_s2s_16_21(data_rsci_idat[161:146]);
  assign Result_acc_114_nl = nl_Result_acc_114_nl[20:0];
  assign nl_Result_acc_71_nl = conv_s2u_21_23(Result_acc_114_nl) + conv_s2u_22_23({(data_rsci_idat[161:144])
      , 4'b0000});
  assign Result_acc_71_nl = nl_Result_acc_71_nl[22:0];
  assign nl_Result_acc_106_nl = conv_s2s_18_19(data_rsci_idat[737:720]) + conv_s2s_16_19({MultLoop_MultLoop_conc_714_15_2
      , (data_rsci_idat[724:723])});
  assign Result_acc_106_nl = nl_Result_acc_106_nl[18:0];
  assign nl_Result_acc_54_nl = conv_s2u_19_20(Result_acc_106_nl) + ({(~ (data_rsci_idat[737:720]))
      , 2'b00});
  assign Result_acc_54_nl = nl_Result_acc_54_nl[19:0];
  assign nl_Result_acc_108_nl = (~ (data_rsci_idat[773:756])) + conv_s2s_15_18({Result_acc_192_cse_1
      , (data_rsci_idat[761:760])});
  assign Result_acc_108_nl = nl_Result_acc_108_nl[17:0];
  assign nl_Result_acc_69_nl = conv_s2u_18_21(Result_acc_108_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[773:756])) , 2'b01});
  assign Result_acc_69_nl = nl_Result_acc_69_nl[20:0];
  assign nl_Result_acc_193_nl = conv_s2s_12_13(data_rsci_idat[809:798]) + 13'b0000000000001;
  assign Result_acc_193_nl = nl_Result_acc_193_nl[12:0];
  assign nl_Result_acc_110_nl = conv_s2s_18_19(data_rsci_idat[809:792]) + conv_s2s_16_19({(Result_acc_193_nl)
      , (data_rsci_idat[797:795])});
  assign Result_acc_110_nl = nl_Result_acc_110_nl[18:0];
  assign nl_Result_acc_58_nl = conv_s2u_19_21(Result_acc_110_nl) + ({(~ (data_rsci_idat[809:792]))
      , 3'b000});
  assign Result_acc_58_nl = nl_Result_acc_58_nl[20:0];
  assign nl_Result_acc_30_nl = conv_s2s_18_21(~ (data_rsci_idat[269:252])) + ({(data_rsci_idat[269:252])
      , 3'b001});
  assign Result_acc_30_nl = nl_Result_acc_30_nl[20:0];
  assign nl_Result_acc_83_nl = (~ (data_rsci_idat[593:576])) + conv_s2s_17_18({MultLoop_MultLoop_conc_772_16_2
      , (data_rsci_idat[579:578])});
  assign Result_acc_83_nl = nl_Result_acc_83_nl[17:0];
  assign nl_Result_acc_62_nl = conv_s2u_18_21(Result_acc_83_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[593:576])) , 2'b01});
  assign Result_acc_62_nl = nl_Result_acc_62_nl[20:0];
  assign nl_MultLoop_acc_1585_itm_1  = conv_s2s_16_18(readslicef_24_16_8((Result_acc_70_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_71_nl))) + conv_s2s_15_18(readslicef_20_15_5((Result_acc_54_nl)))
      + conv_s2s_15_18(readslicef_21_15_6((Result_acc_69_nl))) + conv_s2s_15_18(readslicef_21_15_6((Result_acc_58_nl)))
      + conv_s2s_13_18(readslicef_21_13_8((Result_acc_30_nl))) + conv_s2s_13_18(readslicef_21_13_8((Result_acc_62_nl)));
  assign nl_Result_acc_120_nl = conv_s2s_18_19(data_rsci_idat[341:324]) + conv_s2s_14_19(data_rsci_idat[341:328]);
  assign Result_acc_120_nl = nl_Result_acc_120_nl[18:0];
  assign nl_Result_acc_72_nl = conv_s2u_19_22(Result_acc_120_nl) + conv_s2u_21_22({(data_rsci_idat[341:324])
      , 3'b000});
  assign Result_acc_72_nl = nl_Result_acc_72_nl[21:0];
  assign nl_Result_acc_116_nl = ({(data_rsci_idat[179:162]) , 6'b000001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_718_18_8
      , (~ (data_rsci_idat[169:162]))});
  assign Result_acc_116_nl = nl_Result_acc_116_nl[23:0];
  assign nl_Result_acc_196_nl = conv_s2u_16_18(readslicef_24_16_8((Result_acc_116_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign Result_acc_196_nl = nl_Result_acc_196_nl[17:0];
  assign nl_Result_acc_26_nl = conv_s2u_15_18(data_rsci_idat[197:183]) - (data_rsci_idat[197:180]);
  assign Result_acc_26_nl = nl_Result_acc_26_nl[17:0];
  assign nl_Result_acc_118_nl = ({(data_rsci_idat[215:198]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_746_18_8
      , (~ (data_rsci_idat[205:198]))});
  assign Result_acc_118_nl = nl_Result_acc_118_nl[19:0];
  assign nl_Result_acc_119_nl = conv_s2s_23_24({(data_rsci_idat[215:198]) , 5'b00000})
      + conv_s2s_20_24(Result_acc_118_nl);
  assign Result_acc_119_nl = nl_Result_acc_119_nl[23:0];
  assign nl_Result_acc_198_nl = conv_s2u_16_18(readslicef_24_16_8((Result_acc_119_nl)))
      + (~ (data_rsci_idat[215:198]));
  assign Result_acc_198_nl = nl_Result_acc_198_nl[17:0];
  assign nl_Result_acc_122_nl = ({(data_rsci_idat[413:396]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_722_18_8
      , (~ (data_rsci_idat[403:396]))});
  assign Result_acc_122_nl = nl_Result_acc_122_nl[19:0];
  assign nl_Result_acc_123_nl = conv_s2s_22_23({(data_rsci_idat[413:396]) , 4'b0000})
      + conv_s2s_20_23(Result_acc_122_nl);
  assign Result_acc_123_nl = nl_Result_acc_123_nl[22:0];
  assign nl_Result_acc_200_nl = conv_s2u_15_18(readslicef_23_15_8((Result_acc_123_nl)))
      + (~ (data_rsci_idat[413:396]));
  assign Result_acc_200_nl = nl_Result_acc_200_nl[17:0];
  assign nl_MultLoop_acc_1590_itm_1  = conv_s2s_16_18(MultLoop_acc_4589_itm_19_4)
      + conv_s2s_16_18(readslicef_22_16_6((Result_acc_72_nl))) + conv_s2s_16_18(readslicef_18_16_2((Result_acc_196_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((Result_acc_26_nl))) + conv_s2s_16_18(readslicef_18_16_2((Result_acc_198_nl)))
      + conv_s2s_16_18(~ (data_rsci_idat[287:272])) + conv_s2s_16_18(readslicef_18_16_2((Result_acc_200_nl)))
      + conv_s2s_16_18(MultLoop_acc_3918_itm_17_2);
  assign nl_Result_acc_125_nl = conv_s2s_18_19(data_rsci_idat[485:468]) + conv_s2s_17_19({MultLoop_MultLoop_conc_860_16_4
      , (data_rsci_idat[473:470])});
  assign Result_acc_125_nl = nl_Result_acc_125_nl[18:0];
  assign nl_Result_acc_40_nl = conv_s2u_19_22(Result_acc_125_nl) + ({(~ (data_rsci_idat[485:468]))
      , 4'b0000});
  assign Result_acc_40_nl = nl_Result_acc_40_nl[21:0];
  assign nl_Result_acc_126_nl = conv_s2s_23_24({(~ (data_rsci_idat[539:522])) , 5'b00001})
      + conv_s2s_18_24(~ (data_rsci_idat[539:522]));
  assign Result_acc_126_nl = nl_Result_acc_126_nl[23:0];
  assign nl_Result_acc_43_nl = conv_s2s_24_26(Result_acc_126_nl) + ({(data_rsci_idat[539:522])
      , 8'b00100000});
  assign Result_acc_43_nl = nl_Result_acc_43_nl[25:0];
  assign nl_Result_acc_218_nl = conv_s2u_16_19(Result_acc_127_cse_1[18:3]) + conv_s2u_18_19(data_rsci_idat[575:558]);
  assign Result_acc_218_nl = nl_Result_acc_218_nl[18:0];
  assign nl_Result_acc_220_nl = ({(data_rsci_idat[611:594]) , 4'b0001}) + conv_s2u_19_22(Result_acc_129_cse_1[20:2]);
  assign Result_acc_220_nl = nl_Result_acc_220_nl[21:0];
  assign nl_Result_acc_203_nl = conv_s2u_16_18(readslicef_22_16_6((Result_acc_220_nl)))
      + (~ (data_rsci_idat[611:594]));
  assign Result_acc_203_nl = nl_Result_acc_203_nl[17:0];
  assign nl_MultLoop_acc_1582_itm_1  = conv_s2s_16_18(readslicef_22_16_6((Result_acc_40_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((Result_acc_43_nl))) + conv_s2s_16_18(readslicef_19_16_3((Result_acc_218_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((Result_acc_203_nl)));
  assign nl_Result_acc_48_nl = conv_s2s_25_26({(~ (data_rsci_idat[629:612])) , 7'b0010000})
      + conv_s2s_22_26({(~ (data_rsci_idat[629:612])) , 4'b0100}) + conv_s2s_20_26({(~
      (data_rsci_idat[629:612])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_766_18_7
      , (~ (data_rsci_idat[618:612]))});
  assign Result_acc_48_nl = nl_Result_acc_48_nl[25:0];
  assign nl_Result_acc_205_nl = conv_s2s_11_12(data_rsci_idat[665:655]) + 12'b000000000001;
  assign Result_acc_205_nl = nl_Result_acc_205_nl[11:0];
  assign nl_Result_acc_136_nl = ({(~ (data_rsci_idat[665:648])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[665:648])
      + conv_s2s_17_20({(Result_acc_205_nl) , (data_rsci_idat[654:650])});
  assign Result_acc_136_nl = nl_Result_acc_136_nl[19:0];
  assign nl_Result_acc_74_nl = conv_s2u_20_24(Result_acc_136_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[665:648])) , 5'b00100});
  assign Result_acc_74_nl = nl_Result_acc_74_nl[23:0];
  assign nl_Result_acc_137_nl = conv_s2s_21_22({(~ (data_rsci_idat[683:666])) , 3'b001})
      + conv_s2s_18_22(~ (data_rsci_idat[683:666]));
  assign Result_acc_137_nl = nl_Result_acc_137_nl[21:0];
  assign nl_Result_acc_51_nl = conv_s2s_22_24(Result_acc_137_nl) + ({(data_rsci_idat[683:666])
      , 6'b001000});
  assign Result_acc_51_nl = nl_Result_acc_51_nl[23:0];
  assign nl_Result_acc_140_nl = conv_s2s_21_22({(data_rsci_idat[719:702]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[719:702]) + conv_s2s_16_22({Result_acc_206_cse_1
      , (data_rsci_idat[709:705])});
  assign Result_acc_140_nl = nl_Result_acc_140_nl[21:0];
  assign nl_Result_acc_53_nl = conv_s2u_22_23(Result_acc_140_nl) + ({(~ (data_rsci_idat[719:702]))
      , 5'b00000});
  assign Result_acc_53_nl = nl_Result_acc_53_nl[22:0];
  assign nl_MultLoop_acc_1581_itm_1  = conv_s2s_16_18(readslicef_26_16_10((Result_acc_48_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((Result_acc_74_nl))) + conv_s2s_16_18(readslicef_24_16_8((Result_acc_51_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_53_nl)));
  assign nl_MultLoop_acc_3864_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_15_18(data_rsci_idat[359:345]);
  assign MultLoop_acc_3864_nl = nl_MultLoop_acc_3864_nl[17:0];
  assign nl_MultLoop_acc_3865_nl = ({(data_rsci_idat[359:342]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_3864_nl);
  assign MultLoop_acc_3865_nl = nl_MultLoop_acc_3865_nl[20:0];
  assign nl_MultLoop_acc_1080_nl = conv_s2u_21_24(MultLoop_acc_3865_nl) + conv_s2u_23_24({(data_rsci_idat[359:342])
      , 5'b00000});
  assign MultLoop_acc_1080_nl = nl_MultLoop_acc_1080_nl[23:0];
  assign nl_MultLoop_acc_4565_nl =  -conv_s2s_14_15(data_rsci_idat[287:274]);
  assign MultLoop_acc_4565_nl = nl_MultLoop_acc_4565_nl[14:0];
  assign nl_MultLoop_acc_18_nl = conv_s2s_19_23({(MultLoop_acc_4565_nl) , (~ (data_rsci_idat[273:270]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[287:270])) , 4'b0001});
  assign MultLoop_acc_18_nl = nl_MultLoop_acc_18_nl[22:0];
  assign nl_MultLoop_acc_13_nl = conv_s2s_19_26({MultLoop_MultLoop_conc_698_18_7
      , (~ (data_rsci_idat[186:180]))}) + conv_s2s_25_26({(~ (data_rsci_idat[197:180]))
      , 7'b0000001});
  assign MultLoop_acc_13_nl = nl_MultLoop_acc_13_nl[25:0];
  assign nl_MultLoop_acc_4567_nl = conv_s2u_13_19(MultLoop_acc_3761_itm_19_6[13:1])
      + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_4567_nl = nl_MultLoop_acc_4567_nl[18:0];
  assign nl_MultLoop_acc_3908_nl = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1080_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_18_nl))) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_13_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4567_nl)));
  assign MultLoop_acc_3908_nl = nl_MultLoop_acc_3908_nl[17:0];
  assign nl_MultLoop_acc_15_nl = conv_s2u_10_18(data_rsci_idat[233:224]) - (data_rsci_idat[233:216]);
  assign MultLoop_acc_15_nl = nl_MultLoop_acc_15_nl[17:0];
  assign nl_MultLoop_acc_3854_nl = ({(data_rsci_idat[143:126]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_848_18_7
      , (~ (data_rsci_idat[132:126]))});
  assign MultLoop_acc_3854_nl = nl_MultLoop_acc_3854_nl[22:0];
  assign nl_MultLoop_acc_4559_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3854_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_4559_nl = nl_MultLoop_acc_4559_nl[17:0];
  assign nl_MultLoop_acc_4658_nl = conv_s2u_19_24(MultLoop_acc_3338_itm_20_2_1) +
      ({(data_rsci_idat[35:18]) , 6'b000001});
  assign MultLoop_acc_4658_nl = nl_MultLoop_acc_4658_nl[23:0];
  assign nl_MultLoop_acc_4563_nl = conv_s2u_13_19(MultLoop_acc_1753_itm_19_4[15:3])
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_4563_nl = nl_MultLoop_acc_4563_nl[18:0];
  assign nl_MultLoop_acc_3863_nl = conv_s2s_24_25({(~ (data_rsci_idat[17:0])) , 6'b000100})
      + conv_s2s_21_25(MultLoop_acc_1722_cse_1);
  assign MultLoop_acc_3863_nl = nl_MultLoop_acc_3863_nl[24:0];
  assign nl_MultLoop_acc_2_nl = conv_s2s_25_26(MultLoop_acc_3863_nl) + ({(data_rsci_idat[17:0])
      , 8'b01000000});
  assign MultLoop_acc_2_nl = nl_MultLoop_acc_2_nl[25:0];
  assign nl_MultLoop_acc_4564_nl = conv_s2s_11_12(MultLoop_acc_25_itm_17_5[12:2])
      + 12'b111111011101;
  assign MultLoop_acc_4564_nl = nl_MultLoop_acc_4564_nl[11:0];
  assign nl_MultLoop_acc_4560_nl =  -conv_s2s_12_13(data_rsci_idat[125:114]);
  assign MultLoop_acc_4560_nl = nl_MultLoop_acc_4560_nl[12:0];
  assign nl_MultLoop_acc_3856_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4560_nl)
      , (~ (data_rsci_idat[113:108]))});
  assign MultLoop_acc_3856_nl = nl_MultLoop_acc_3856_nl[20:0];
  assign nl_MultLoop_acc_4561_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_3856_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_4561_nl = nl_MultLoop_acc_4561_nl[17:0];
  assign nl_MultLoop_acc_4562_nl = conv_s2s_10_11(data_rsci_idat[89:80]) + 11'b00000000001;
  assign MultLoop_acc_4562_nl = nl_MultLoop_acc_4562_nl[10:0];
  assign nl_MultLoop_acc_3858_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_15_18({(MultLoop_acc_4562_nl)
      , (data_rsci_idat[79:76])});
  assign MultLoop_acc_3858_nl = nl_MultLoop_acc_3858_nl[17:0];
  assign nl_MultLoop_acc_3859_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3858_nl);
  assign MultLoop_acc_3859_nl = nl_MultLoop_acc_3859_nl[19:0];
  assign nl_MultLoop_acc_7_nl = conv_s2u_20_22(MultLoop_acc_3859_nl) + ({(~ (data_rsci_idat[89:72]))
      , 4'b0000});
  assign MultLoop_acc_7_nl = nl_MultLoop_acc_7_nl[21:0];
  assign nl_MultLoop_acc_38_nl = conv_s2u_14_18(data_rsci_idat[665:652]) - (data_rsci_idat[665:648]);
  assign MultLoop_acc_38_nl = nl_MultLoop_acc_38_nl[17:0];
  assign nl_MultLoop_acc_27_nl = conv_s2u_14_18(data_rsci_idat[449:436]) - (data_rsci_idat[449:432]);
  assign MultLoop_acc_27_nl = nl_MultLoop_acc_27_nl[17:0];
  assign nl_MultLoop_acc_3913_itm_1  = (MultLoop_acc_3908_nl) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_15_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4559_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_4658_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4563_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_2_nl)))
      + conv_s2s_14_18({(MultLoop_acc_4564_nl) , (MultLoop_acc_25_itm_17_5[1:0])})
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4561_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_7_nl)))
      + conv_s2s_13_18(readslicef_18_13_5((MultLoop_acc_38_nl))) + conv_s2s_13_18(readslicef_18_13_5((MultLoop_acc_27_nl)));
  assign nl_MultLoop_acc_3799_nl = ({(data_rsci_idat[827:810]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[827:810]));
  assign MultLoop_acc_3799_nl = nl_MultLoop_acc_3799_nl[19:0];
  assign nl_MultLoop_acc_3800_nl = ({(~ (data_rsci_idat[827:810])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3799_nl);
  assign MultLoop_acc_3800_nl = nl_MultLoop_acc_3800_nl[21:0];
  assign nl_MultLoop_acc_46_nl = conv_s2s_22_24(MultLoop_acc_3800_nl) + ({(data_rsci_idat[827:810])
      , 6'b010000});
  assign MultLoop_acc_46_nl = nl_MultLoop_acc_46_nl[23:0];
  assign nl_MultLoop_acc_45_nl = conv_s2u_12_18(data_rsci_idat[809:798]) - (data_rsci_idat[809:792]);
  assign MultLoop_acc_45_nl = nl_MultLoop_acc_45_nl[17:0];
  assign nl_MultLoop_acc_4568_nl = conv_s2s_12_13(data_rsci_idat[341:330]) + 13'b0000000000001;
  assign MultLoop_acc_4568_nl = nl_MultLoop_acc_4568_nl[12:0];
  assign nl_MultLoop_acc_3803_nl = conv_s2s_18_19(data_rsci_idat[341:324]) + conv_s2s_16_19({(MultLoop_acc_4568_nl)
      , (data_rsci_idat[329:327])});
  assign MultLoop_acc_3803_nl = nl_MultLoop_acc_3803_nl[18:0];
  assign nl_MultLoop_acc_21_nl = conv_s2u_19_21(MultLoop_acc_3803_nl) + ({(~ (data_rsci_idat[341:324]))
      , 3'b000});
  assign MultLoop_acc_21_nl = nl_MultLoop_acc_21_nl[20:0];
  assign nl_MultLoop_acc_3881_itm_1  = conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_46_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_45_nl))) + conv_s2s_14_16(MultLoop_acc_3190_itm_19_4[15:2])
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_21_nl)));
  assign nl_MultLoop_acc_4569_nl =  -conv_s2s_13_14(data_rsci_idat[845:833]);
  assign MultLoop_acc_4569_nl = nl_MultLoop_acc_4569_nl[13:0];
  assign nl_MultLoop_acc_3805_nl = ({(data_rsci_idat[845:828]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4569_nl)
      , (~ (data_rsci_idat[832:828]))});
  assign MultLoop_acc_3805_nl = nl_MultLoop_acc_3805_nl[20:0];
  assign nl_MultLoop_acc_47_nl = conv_s2s_21_23(MultLoop_acc_3805_nl) + ({(~ (data_rsci_idat[845:828]))
      , 5'b00000});
  assign MultLoop_acc_47_nl = nl_MultLoop_acc_47_nl[22:0];
  assign nl_MultLoop_acc_4659_nl = conv_s2u_14_18(MultLoop_acc_2220_cse_1[18:5])
      + (~ (data_rsci_idat[719:702]));
  assign MultLoop_acc_4659_nl = nl_MultLoop_acc_4659_nl[17:0];
  assign nl_MultLoop_acc_3880_itm_1  = conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_47_nl)))
      + conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4659_nl)));
  assign nl_MultLoop_acc_3810_nl = ({(data_rsci_idat[683:666]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[683:666])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_816_18_7
      , (~ (data_rsci_idat[672:666]))});
  assign MultLoop_acc_3810_nl = nl_MultLoop_acc_3810_nl[21:0];
  assign nl_MultLoop_acc_4572_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_3810_nl)))
      + (~ (data_rsci_idat[683:666]));
  assign MultLoop_acc_4572_nl = nl_MultLoop_acc_4572_nl[17:0];
  assign nl_MultLoop_acc_3813_nl = ({(data_rsci_idat[611:594]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[611:594])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_750_18_7
      , (~ (data_rsci_idat[600:594]))});
  assign MultLoop_acc_3813_nl = nl_MultLoop_acc_3813_nl[22:0];
  assign nl_MultLoop_acc_4574_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3813_nl)))
      + (~ (data_rsci_idat[611:594]));
  assign MultLoop_acc_4574_nl = nl_MultLoop_acc_4574_nl[17:0];
  assign nl_MultLoop_acc_33_nl = conv_s2u_12_18(data_rsci_idat[575:564]) - (data_rsci_idat[575:558]);
  assign MultLoop_acc_33_nl = nl_MultLoop_acc_33_nl[17:0];
  assign nl_MultLoop_acc_3896_itm_1  = conv_s2s_15_17(data_rsci_idat[737:723]) +
      conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4572_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4574_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_33_nl)));
  assign nl_MultLoop_acc_4660_nl = conv_s2u_19_21(MultLoop_acc_2387_cse_1[20:2])
      + ({(data_rsci_idat[593:576]) , 3'b001});
  assign MultLoop_acc_4660_nl = nl_MultLoop_acc_4660_nl[20:0];
  assign nl_MultLoop_acc_4661_nl = conv_s2u_19_20(MultLoop_acc_1811_itm_20_2_1) +
      ({(data_rsci_idat[557:540]) , 2'b01});
  assign MultLoop_acc_4661_nl = nl_MultLoop_acc_4661_nl[19:0];
  assign nl_MultLoop_acc_3818_nl = ({(data_rsci_idat[503:486]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_716_18_7
      , (~ (data_rsci_idat[492:486]))});
  assign MultLoop_acc_3818_nl = nl_MultLoop_acc_3818_nl[21:0];
  assign nl_MultLoop_acc_4576_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_3818_nl)))
      + (~ (data_rsci_idat[503:486]));
  assign MultLoop_acc_4576_nl = nl_MultLoop_acc_4576_nl[17:0];
  assign nl_MultLoop_acc_3895_itm_1  = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_4660_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_4661_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4576_nl)))
      + conv_s2s_15_17(MultLoop_acc_4587_itm_18_3[15:1]);
  assign nl_MultLoop_acc_3820_nl = ({(~ (data_rsci_idat[323:306])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_3661_cse_1);
  assign MultLoop_acc_3820_nl = nl_MultLoop_acc_3820_nl[19:0];
  assign nl_MultLoop_acc_1079_nl = conv_s2u_20_22(MultLoop_acc_3820_nl) + ({(data_rsci_idat[323:306])
      , 4'b0100});
  assign MultLoop_acc_1079_nl = nl_MultLoop_acc_1079_nl[21:0];
  assign nl_MultLoop_acc_3823_nl = ({(~ (data_rsci_idat[179:162])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[179:162])
      + conv_s2s_17_20({MultLoop_MultLoop_conc_798_16_4 , (data_rsci_idat[167:164])});
  assign MultLoop_acc_3823_nl = nl_MultLoop_acc_3823_nl[19:0];
  assign nl_MultLoop_acc_1076_nl = conv_s2u_20_23(MultLoop_acc_3823_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[179:162])) , 4'b0100});
  assign MultLoop_acc_1076_nl = nl_MultLoop_acc_1076_nl[22:0];
  assign nl_MultLoop_acc_3825_nl = conv_s2s_23_24({(~ (data_rsci_idat[161:144]))
      , 5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[161:144])) , 2'b01}) + conv_s2s_18_24(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_3825_nl = nl_MultLoop_acc_3825_nl[23:0];
  assign nl_MultLoop_acc_11_nl = conv_s2s_24_25(MultLoop_acc_3825_nl) + ({(data_rsci_idat[161:144])
      , 7'b0100000});
  assign MultLoop_acc_11_nl = nl_MultLoop_acc_11_nl[24:0];
  assign nl_MultLoop_acc_3827_nl = ({(~ (data_rsci_idat[71:54])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[71:54])
      + conv_s2s_15_20(data_rsci_idat[71:57]);
  assign MultLoop_acc_3827_nl = nl_MultLoop_acc_3827_nl[19:0];
  assign nl_MultLoop_acc_1075_nl = conv_s2u_20_22(MultLoop_acc_3827_nl) + ({(data_rsci_idat[71:54])
      , 4'b0100});
  assign MultLoop_acc_1075_nl = nl_MultLoop_acc_1075_nl[21:0];
  assign nl_MultLoop_acc_3894_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1079_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1076_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_11_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1075_nl)));
  assign nl_MultLoop_acc_3832_nl = conv_s2s_18_19(data_rsci_idat[773:756]) + conv_s2s_17_19({Result_acc_192_cse_1
      , (data_rsci_idat[761:758])});
  assign MultLoop_acc_3832_nl = nl_MultLoop_acc_3832_nl[18:0];
  assign nl_MultLoop_acc_43_nl = conv_s2u_19_22(MultLoop_acc_3832_nl) + ({(~ (data_rsci_idat[773:756]))
      , 4'b0000});
  assign MultLoop_acc_43_nl = nl_MultLoop_acc_43_nl[21:0];
  assign nl_MultLoop_acc_4580_nl = conv_s2s_12_13(data_rsci_idat[701:690]) + 13'b0000000000001;
  assign MultLoop_acc_4580_nl = nl_MultLoop_acc_4580_nl[12:0];
  assign nl_MultLoop_acc_3834_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_17_18({(MultLoop_acc_4580_nl)
      , (data_rsci_idat[689:686])});
  assign MultLoop_acc_3834_nl = nl_MultLoop_acc_3834_nl[17:0];
  assign nl_MultLoop_acc_3835_nl = ({(data_rsci_idat[701:684]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3834_nl);
  assign MultLoop_acc_3835_nl = nl_MultLoop_acc_3835_nl[19:0];
  assign nl_MultLoop_acc_40_nl = conv_s2u_20_22(MultLoop_acc_3835_nl) + ({(~ (data_rsci_idat[701:684]))
      , 4'b0000});
  assign MultLoop_acc_40_nl = nl_MultLoop_acc_40_nl[21:0];
  assign nl_MultLoop_acc_1087_nl = conv_s2u_18_21(MultLoop_acc_1946_cse_1) + ({(data_rsci_idat[791:774])
      , 3'b001});
  assign MultLoop_acc_1087_nl = nl_MultLoop_acc_1087_nl[20:0];
  assign nl_MultLoop_acc_3830_nl = (~ (data_rsci_idat[863:846])) + conv_s2s_15_18({MultLoop_acc_3961_cse_1
      , (data_rsci_idat[851:850])});
  assign MultLoop_acc_3830_nl = nl_MultLoop_acc_3830_nl[17:0];
  assign nl_MultLoop_acc_1088_nl = conv_s2u_18_21(MultLoop_acc_3830_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[863:846])) , 2'b01});
  assign MultLoop_acc_1088_nl = nl_MultLoop_acc_1088_nl[20:0];
  assign nl_MultLoop_acc_42_nl = conv_s2u_14_18(data_rsci_idat[755:742]) - (data_rsci_idat[755:738]);
  assign MultLoop_acc_42_nl = nl_MultLoop_acc_42_nl[17:0];
  assign nl_MultLoop_acc_4581_nl = (~ (data_rsci_idat[647:630])) + conv_s2s_15_18(MultLoop_acc_3281_itm_20_6);
  assign MultLoop_acc_4581_nl = nl_MultLoop_acc_4581_nl[17:0];
  assign nl_MultLoop_acc_4582_nl = conv_s2u_18_20(MultLoop_acc_4581_nl) + ({(data_rsci_idat[647:630])
      , 2'b01});
  assign MultLoop_acc_4582_nl = nl_MultLoop_acc_4582_nl[19:0];
  assign nl_MultLoop_acc_3911_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_43_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_40_nl))) + conv_s2s_16_18(data_rsci_idat[467:452])
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1087_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1088_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_42_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_4582_nl)))
      + conv_s2s_16_18(MultLoop_acc_1943_itm_18_2[16:1]);
  assign nl_MultLoop_acc_4586_nl = conv_s2s_11_12(data_rsci_idat[305:295]) + 12'b000000000001;
  assign MultLoop_acc_4586_nl = nl_MultLoop_acc_4586_nl[11:0];
  assign nl_MultLoop_acc_3847_nl = ({(~ (data_rsci_idat[305:288])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[305:288])
      + conv_s2s_17_21({(MultLoop_acc_4586_nl) , (data_rsci_idat[294:290])});
  assign MultLoop_acc_3847_nl = nl_MultLoop_acc_3847_nl[20:0];
  assign nl_MultLoop_acc_1078_nl = conv_s2u_21_24(MultLoop_acc_3847_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[305:288])) , 5'b01000});
  assign MultLoop_acc_1078_nl = nl_MultLoop_acc_1078_nl[23:0];
  assign nl_MultLoop_acc_3849_nl = ({(~ (data_rsci_idat[251:234])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2591_cse_1);
  assign MultLoop_acc_3849_nl = nl_MultLoop_acc_3849_nl[19:0];
  assign nl_MultLoop_acc_3850_nl = conv_s2s_22_23({(~ (data_rsci_idat[251:234]))
      , 4'b0100}) + conv_s2s_20_23(MultLoop_acc_3849_nl);
  assign MultLoop_acc_3850_nl = nl_MultLoop_acc_3850_nl[22:0];
  assign nl_MultLoop_acc_1077_nl = conv_s2u_23_24(MultLoop_acc_3850_nl) + ({(data_rsci_idat[251:234])
      , 6'b010000});
  assign MultLoop_acc_1077_nl = nl_MultLoop_acc_1077_nl[23:0];
  assign nl_MultLoop_acc_4583_nl =  -conv_s2s_15_16(data_rsci_idat[539:525]);
  assign MultLoop_acc_4583_nl = nl_MultLoop_acc_4583_nl[15:0];
  assign nl_MultLoop_acc_31_nl = conv_s2s_19_22({(MultLoop_acc_4583_nl) , (~ (data_rsci_idat[524:522]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[539:522])) , 3'b001});
  assign MultLoop_acc_31_nl = nl_MultLoop_acc_31_nl[21:0];
  assign nl_MultLoop_acc_1084_nl = conv_s2u_18_22(MultLoop_acc_2133_cse_1) + ({(data_rsci_idat[521:504])
      , 4'b0001});
  assign MultLoop_acc_1084_nl = nl_MultLoop_acc_1084_nl[21:0];
  assign nl_MultLoop_acc_3841_nl = conv_s2s_20_21({(~ (data_rsci_idat[485:468]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2535_cse_1);
  assign MultLoop_acc_3841_nl = nl_MultLoop_acc_3841_nl[20:0];
  assign nl_MultLoop_acc_1083_nl = conv_s2u_21_22(MultLoop_acc_3841_nl) + ({(data_rsci_idat[485:468])
      , 4'b0100});
  assign MultLoop_acc_1083_nl = nl_MultLoop_acc_1083_nl[21:0];
  assign nl_MultLoop_acc_3844_nl = conv_s2s_20_21({(data_rsci_idat[377:360]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[377:360]) + conv_s2s_17_21({MultLoop_acc_4229_cse_1
      , (data_rsci_idat[367:362])});
  assign MultLoop_acc_3844_nl = nl_MultLoop_acc_3844_nl[20:0];
  assign nl_MultLoop_acc_4585_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_3844_nl)))
      + (~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_4585_nl = nl_MultLoop_acc_4585_nl[17:0];
  assign nl_MultLoop_acc_17_nl = conv_s2s_18_24(~ (data_rsci_idat[269:252])) + ({(data_rsci_idat[269:252])
      , 6'b000001});
  assign MultLoop_acc_17_nl = nl_MultLoop_acc_17_nl[23:0];
  assign nl_MultLoop_acc_3852_nl = conv_s2s_24_25({(~ (data_rsci_idat[215:198]))
      , 6'b001000}) + conv_s2s_22_25(MultLoop_acc_3099_cse_1);
  assign MultLoop_acc_3852_nl = nl_MultLoop_acc_3852_nl[24:0];
  assign nl_MultLoop_acc_14_nl = conv_s2s_25_26(MultLoop_acc_3852_nl) + ({(data_rsci_idat[215:198])
      , 8'b01000000});
  assign MultLoop_acc_14_nl = nl_MultLoop_acc_14_nl[25:0];
  assign nl_MultLoop_acc_3910_itm_1  = conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1078_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1077_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_31_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1084_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1083_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4585_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_17_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_14_nl)));
  assign nl_MultLoop_acc_3940_nl = conv_s2s_11_12(data_rsci_idat[539:529]) + 12'b000000000001;
  assign MultLoop_acc_3940_nl = nl_MultLoop_acc_3940_nl[11:0];
  assign nl_MultLoop_acc_1640_nl = ({(~ (data_rsci_idat[539:522])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[539:522])
      + conv_s2s_17_21({(MultLoop_acc_3940_nl) , (data_rsci_idat[528:524])});
  assign MultLoop_acc_1640_nl = nl_MultLoop_acc_1640_nl[20:0];
  assign nl_MultLoop_acc_1443_nl = conv_s2u_21_24(MultLoop_acc_1640_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[539:522])) , 5'b01000});
  assign MultLoop_acc_1443_nl = nl_MultLoop_acc_1443_nl[23:0];
  assign nl_MultLoop_acc_1642_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_16_18({MultLoop_acc_3941_cse_1
      , (data_rsci_idat[240:237])});
  assign MultLoop_acc_1642_nl = nl_MultLoop_acc_1642_nl[17:0];
  assign nl_MultLoop_acc_1435_nl = conv_s2u_18_23(MultLoop_acc_1642_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[251:234])) , 4'b0001});
  assign MultLoop_acc_1435_nl = nl_MultLoop_acc_1435_nl[22:0];
  assign nl_Result_acc_207_nl = conv_s2s_13_14(data_rsci_idat[647:635]) + 14'b00000000000001;
  assign Result_acc_207_nl = nl_Result_acc_207_nl[13:0];
  assign nl_Result_acc_171_nl = (~ (data_rsci_idat[647:630])) + conv_s2s_17_18({(Result_acc_207_nl)
      , (data_rsci_idat[634:632])});
  assign Result_acc_171_nl = nl_Result_acc_171_nl[17:0];
  assign nl_Result_acc_80_nl = conv_s2u_18_22(Result_acc_171_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[647:630])) , 3'b001});
  assign Result_acc_80_nl = nl_Result_acc_80_nl[21:0];
  assign nl_Result_acc_8_nl = conv_s2s_25_26({(~ (data_rsci_idat[719:702])) , 7'b0000100})
      + conv_s2s_20_26({(~ (data_rsci_idat[719:702])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_840_18_7
      , (~ (data_rsci_idat[708:702]))});
  assign Result_acc_8_nl = nl_Result_acc_8_nl[25:0];
  assign nl_MultLoop_acc_1683_itm_1  = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1443_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1435_nl))) + conv_s2s_17_18(readslicef_22_17_5((Result_acc_80_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((Result_acc_8_nl)));
  assign nl_Result_acc_11_nl = conv_s2s_26_27({(~ (data_rsci_idat[773:756])) , 8'b00000100})
      + conv_s2s_20_27({(~ (data_rsci_idat[773:756])) , 2'b01}) + conv_s2s_19_27({MultLoop_MultLoop_conc_846_18_8
      , (~ (data_rsci_idat[763:756]))});
  assign Result_acc_11_nl = nl_Result_acc_11_nl[26:0];
  assign nl_Result_acc_16_nl = conv_s2s_25_26({(~ (data_rsci_idat[863:846])) , 7'b0000100})
      + conv_s2s_20_26({(~ (data_rsci_idat[863:846])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_720_18_7
      , (~ (data_rsci_idat[852:846]))});
  assign Result_acc_16_nl = nl_Result_acc_16_nl[25:0];
  assign nl_MultLoop_acc_1673_itm_1  = conv_s2s_17_18(readslicef_27_17_10((Result_acc_11_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((Result_acc_16_nl)));
  assign nl_MultLoop_acc_3942_nl =  -conv_s2s_12_13(data_rsci_idat[557:546]);
  assign MultLoop_acc_3942_nl = nl_MultLoop_acc_3942_nl[12:0];
  assign nl_MultLoop_acc_1596_nl = ({(data_rsci_idat[557:540]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_3942_nl)
      , (~ (data_rsci_idat[545:540]))});
  assign MultLoop_acc_1596_nl = nl_MultLoop_acc_1596_nl[19:0];
  assign nl_MultLoop_acc_3943_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_1596_nl)))
      + (~ (data_rsci_idat[557:540]));
  assign MultLoop_acc_3943_nl = nl_MultLoop_acc_3943_nl[17:0];
  assign nl_MultLoop_acc_1597_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_14_18(data_rsci_idat[395:382]);
  assign MultLoop_acc_1597_nl = nl_MultLoop_acc_1597_nl[17:0];
  assign nl_MultLoop_acc_1439_nl = conv_s2u_18_20(MultLoop_acc_1597_nl) + ({(data_rsci_idat[395:378])
      , 2'b01});
  assign MultLoop_acc_1439_nl = nl_MultLoop_acc_1439_nl[19:0];
  assign nl_MultLoop_acc_1599_nl = (~ (data_rsci_idat[305:288])) + conv_s2s_17_18({MultLoop_MultLoop_conc_706_16_4
      , (data_rsci_idat[293:290])});
  assign MultLoop_acc_1599_nl = nl_MultLoop_acc_1599_nl[17:0];
  assign nl_MultLoop_acc_1600_nl = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1599_nl);
  assign MultLoop_acc_1600_nl = nl_MultLoop_acc_1600_nl[19:0];
  assign nl_MultLoop_acc_1059_nl = conv_s2u_20_22(MultLoop_acc_1600_nl) + ({(~ (data_rsci_idat[305:288]))
      , 4'b0000});
  assign MultLoop_acc_1059_nl = nl_MultLoop_acc_1059_nl[21:0];
  assign nl_MultLoop_acc_1659_itm_1  = conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_3943_nl)))
      + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_1439_nl))) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_1059_nl)))
      + conv_s2s_14_16(data_rsci_idat[323:310]);
  assign nl_MultLoop_acc_3945_nl =  -conv_s2s_13_14(data_rsci_idat[125:113]);
  assign MultLoop_acc_3945_nl = nl_MultLoop_acc_3945_nl[13:0];
  assign nl_MultLoop_acc_1049_nl = conv_s2s_23_24({(~ (data_rsci_idat[125:108]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[125:108])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_3945_nl)
      , (~ (data_rsci_idat[112:108]))});
  assign MultLoop_acc_1049_nl = nl_MultLoop_acc_1049_nl[23:0];
  assign nl_Result_acc_153_nl = ({(data_rsci_idat[665:648]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[665:648]));
  assign Result_acc_153_nl = nl_Result_acc_153_nl[19:0];
  assign nl_Result_acc_5_nl = conv_s2s_20_23(Result_acc_153_nl) + conv_s2s_22_23({(data_rsci_idat[665:648])
      , 4'b0000});
  assign Result_acc_5_nl = nl_Result_acc_5_nl[22:0];
  assign nl_Result_acc_222_nl = conv_s2u_18_20(MultLoop_asn_1479) + ({(data_rsci_idat[683:666])
      , 2'b01});
  assign Result_acc_222_nl = nl_Result_acc_222_nl[19:0];
  assign nl_Result_acc_7_nl = conv_s2u_12_18(data_rsci_idat[701:690]) - (data_rsci_idat[701:684]);
  assign Result_acc_7_nl = nl_Result_acc_7_nl[17:0];
  assign nl_MultLoop_acc_1658_itm_1  = conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_1049_nl)))
      + conv_s2s_14_16(readslicef_23_14_9((Result_acc_5_nl))) + conv_s2s_14_16(readslicef_20_14_6((Result_acc_222_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((Result_acc_7_nl)));
  assign nl_MultLoop_acc_1604_nl = conv_s2s_23_24({(~ (data_rsci_idat[521:504]))
      , 5'b01000}) + conv_s2s_22_24(MultLoop_acc_1603_cse_1);
  assign MultLoop_acc_1604_nl = nl_MultLoop_acc_1604_nl[23:0];
  assign nl_MultLoop_acc_1070_nl = conv_s2s_24_25(MultLoop_acc_1604_nl) + ({(data_rsci_idat[521:504])
      , 7'b0100000});
  assign MultLoop_acc_1070_nl = nl_MultLoop_acc_1070_nl[24:0];
  assign nl_MultLoop_acc_1068_nl = conv_s2s_18_23(~ (data_rsci_idat[485:468])) +
      ({(data_rsci_idat[485:468]) , 5'b00001});
  assign MultLoop_acc_1068_nl = nl_MultLoop_acc_1068_nl[22:0];
  assign nl_MultLoop_acc_1605_nl = (~ (data_rsci_idat[449:432])) + conv_s2s_16_18(data_rsci_idat[449:434]);
  assign MultLoop_acc_1605_nl = nl_MultLoop_acc_1605_nl[17:0];
  assign nl_MultLoop_acc_1606_nl = conv_s2s_20_21({(~ (data_rsci_idat[449:432]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1605_nl);
  assign MultLoop_acc_1606_nl = nl_MultLoop_acc_1606_nl[20:0];
  assign nl_MultLoop_acc_1441_nl = conv_s2u_21_22(MultLoop_acc_1606_nl) + ({(data_rsci_idat[449:432])
      , 4'b0100});
  assign MultLoop_acc_1441_nl = nl_MultLoop_acc_1441_nl[21:0];
  assign nl_Result_acc_211_nl = conv_s2s_14_15(data_rsci_idat[737:724]) + 15'b000000000000001;
  assign Result_acc_211_nl = nl_Result_acc_211_nl[14:0];
  assign nl_Result_acc_157_nl = conv_s2s_18_19(data_rsci_idat[737:720]) + conv_s2s_17_19({(Result_acc_211_nl)
      , (data_rsci_idat[723:722])});
  assign Result_acc_157_nl = nl_Result_acc_157_nl[18:0];
  assign nl_Result_acc_9_nl = conv_s2u_19_20(Result_acc_157_nl) + ({(~ (data_rsci_idat[737:720]))
      , 2'b00});
  assign Result_acc_9_nl = nl_Result_acc_9_nl[19:0];
  assign nl_MultLoop_acc_1442_nl = conv_s2u_15_19(data_rsci_idat[503:489]) + conv_s2u_18_19(data_rsci_idat[503:486]);
  assign MultLoop_acc_1442_nl = nl_MultLoop_acc_1442_nl[18:0];
  assign nl_MultLoop_acc_1671_itm_1  = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1070_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1068_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1441_nl)))
      + conv_s2s_14_17(readslicef_20_14_6((Result_acc_9_nl))) + conv_s2s_13_17(readslicef_19_13_6((MultLoop_acc_1442_nl)));
  assign nl_MultLoop_acc_1609_nl = ({(~ (data_rsci_idat[413:396])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[413:396])
      + conv_s2s_17_20({MultLoop_acc_3946_cse_1 , (data_rsci_idat[401:398])});
  assign MultLoop_acc_1609_nl = nl_MultLoop_acc_1609_nl[19:0];
  assign nl_MultLoop_acc_1440_nl = conv_s2u_20_23(MultLoop_acc_1609_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[413:396])) , 4'b0100});
  assign MultLoop_acc_1440_nl = nl_MultLoop_acc_1440_nl[22:0];
  assign nl_MultLoop_acc_1610_nl = ({(data_rsci_idat[377:360]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[377:360]));
  assign MultLoop_acc_1610_nl = nl_MultLoop_acc_1610_nl[19:0];
  assign nl_MultLoop_acc_1062_nl = conv_s2s_20_25(MultLoop_acc_1610_nl) + conv_s2s_24_25({(data_rsci_idat[377:360])
      , 6'b000000});
  assign MultLoop_acc_1062_nl = nl_MultLoop_acc_1062_nl[24:0];
  assign nl_MultLoop_acc_1612_nl = ({(~ (data_rsci_idat[269:252])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_1611_cse_1);
  assign MultLoop_acc_1612_nl = nl_MultLoop_acc_1612_nl[19:0];
  assign nl_MultLoop_acc_1436_nl = conv_s2u_20_22(MultLoop_acc_1612_nl) + ({(data_rsci_idat[269:252])
      , 4'b0100});
  assign MultLoop_acc_1436_nl = nl_MultLoop_acc_1436_nl[21:0];
  assign nl_MultLoop_acc_1053_nl = conv_s2s_24_25({(~ (data_rsci_idat[197:180]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[197:180])) , 4'b0001}) +
      conv_s2s_19_25({MultLoop_MultLoop_conc_862_18_6 , (~ (data_rsci_idat[185:180]))});
  assign MultLoop_acc_1053_nl = nl_MultLoop_acc_1053_nl[24:0];
  assign nl_MultLoop_acc_1670_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1440_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1062_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1436_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1053_nl)));
  assign nl_MultLoop_acc_1615_nl = ({(data_rsci_idat[215:198]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[215:198]));
  assign MultLoop_acc_1615_nl = nl_MultLoop_acc_1615_nl[19:0];
  assign nl_MultLoop_acc_1616_nl = ({(~ (data_rsci_idat[215:198])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_1615_nl);
  assign MultLoop_acc_1616_nl = nl_MultLoop_acc_1616_nl[22:0];
  assign nl_MultLoop_acc_1054_nl = conv_s2s_23_25(MultLoop_acc_1616_nl) + ({(data_rsci_idat[215:198])
      , 7'b0100000});
  assign MultLoop_acc_1054_nl = nl_MultLoop_acc_1054_nl[24:0];
  assign nl_MultLoop_acc_1051_nl = conv_s2s_18_21(~ (data_rsci_idat[161:144])) +
      ({(data_rsci_idat[161:144]) , 3'b001});
  assign MultLoop_acc_1051_nl = nl_MultLoop_acc_1051_nl[20:0];
  assign nl_MultLoop_acc_4662_nl = ({(data_rsci_idat[107:90]) , 3'b001}) + conv_s2u_19_21(MultLoop_acc_1618_cse_1[20:2]);
  assign MultLoop_acc_4662_nl = nl_MultLoop_acc_4662_nl[20:0];
  assign nl_MultLoop_acc_3949_nl = conv_s2u_16_18(readslicef_21_16_5((MultLoop_acc_4662_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_3949_nl = nl_MultLoop_acc_3949_nl[17:0];
  assign nl_Result_acc_160_nl = ({(data_rsci_idat[629:612]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[629:612])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_766_18_7
      , (~ (data_rsci_idat[618:612]))});
  assign Result_acc_160_nl = nl_Result_acc_160_nl[22:0];
  assign nl_Result_acc_213_nl = conv_s2u_16_18(readslicef_23_16_7((Result_acc_160_nl)))
      + (~ (data_rsci_idat[629:612]));
  assign Result_acc_213_nl = nl_Result_acc_213_nl[17:0];
  assign nl_MultLoop_acc_1669_itm_1  = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1054_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1051_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_3949_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((Result_acc_213_nl)));
  assign nl_MultLoop_acc_3950_nl = conv_s2s_11_12(data_rsci_idat[467:457]) + 12'b000000000001;
  assign MultLoop_acc_3950_nl = nl_MultLoop_acc_3950_nl[11:0];
  assign nl_MultLoop_acc_1621_nl = conv_s2s_18_19(data_rsci_idat[467:450]) + conv_s2s_16_19({(MultLoop_acc_3950_nl)
      , (data_rsci_idat[456:453])});
  assign MultLoop_acc_1621_nl = nl_MultLoop_acc_1621_nl[18:0];
  assign nl_MultLoop_acc_1067_nl = conv_s2u_19_22(MultLoop_acc_1621_nl) + ({(~ (data_rsci_idat[467:450]))
      , 4'b0000});
  assign MultLoop_acc_1067_nl = nl_MultLoop_acc_1067_nl[21:0];
  assign nl_Result_acc_161_nl = (~ (data_rsci_idat[791:774])) + conv_s2s_14_18(data_rsci_idat[791:778]);
  assign Result_acc_161_nl = nl_Result_acc_161_nl[17:0];
  assign nl_Result_acc_81_nl = conv_s2u_18_21(Result_acc_161_nl) + ({(data_rsci_idat[791:774])
      , 3'b001});
  assign Result_acc_81_nl = nl_Result_acc_81_nl[20:0];
  assign nl_Result_acc_nl = conv_s2u_18_20(Result_acc_152_cse_1) + ({(data_rsci_idat[593:576])
      , 2'b01});
  assign Result_acc_nl = nl_Result_acc_nl[19:0];
  assign nl_Result_acc_2_nl = conv_s2u_16_18(data_rsci_idat[611:596]) - (data_rsci_idat[611:594]);
  assign Result_acc_2_nl = nl_Result_acc_2_nl[17:0];
  assign nl_MultLoop_acc_1643_nl = conv_s2s_10_11(readslicef_18_10_8((Result_acc_2_nl)))
      + 11'b00010010011;
  assign MultLoop_acc_1643_nl = nl_MultLoop_acc_1643_nl[10:0];
  assign nl_MultLoop_acc_1073_nl = conv_s2u_16_18(data_rsci_idat[575:560]) - (data_rsci_idat[575:558]);
  assign MultLoop_acc_1073_nl = nl_MultLoop_acc_1073_nl[17:0];
  assign nl_MultLoop_acc_1668_itm_1  = conv_s2s_16_17(readslicef_22_16_6((MultLoop_acc_1067_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((Result_acc_81_nl))) + conv_s2s_13_17(readslicef_20_13_7((Result_acc_nl)))
      + conv_s2s_11_17(MultLoop_acc_1643_nl) + conv_s2s_11_17(readslicef_18_11_7((MultLoop_acc_1073_nl)));
  assign nl_MultLoop_acc_1627_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_13_18(data_rsci_idat[233:221]);
  assign MultLoop_acc_1627_nl = nl_MultLoop_acc_1627_nl[17:0];
  assign nl_MultLoop_acc_1434_nl = conv_s2u_18_20(MultLoop_acc_1627_nl) + ({(data_rsci_idat[233:216])
      , 2'b01});
  assign MultLoop_acc_1434_nl = nl_MultLoop_acc_1434_nl[19:0];
  assign nl_MultLoop_acc_3952_nl = conv_s2s_10_11(data_rsci_idat[179:170]) + 11'b00000000001;
  assign MultLoop_acc_3952_nl = nl_MultLoop_acc_3952_nl[10:0];
  assign nl_MultLoop_acc_1630_nl = conv_s2s_21_22({(data_rsci_idat[179:162]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[179:162]) + conv_s2s_16_22({(MultLoop_acc_3952_nl)
      , (data_rsci_idat[169:165])});
  assign MultLoop_acc_1630_nl = nl_MultLoop_acc_1630_nl[21:0];
  assign nl_MultLoop_acc_1052_nl = conv_s2u_22_23(MultLoop_acc_1630_nl) + ({(~ (data_rsci_idat[179:162]))
      , 5'b00000});
  assign MultLoop_acc_1052_nl = nl_MultLoop_acc_1052_nl[22:0];
  assign nl_MultLoop_acc_1065_nl = conv_s2s_25_26({(~ (data_rsci_idat[431:414]))
      , 7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[431:414])) , 5'b00001})
      + conv_s2s_19_26({MultLoop_MultLoop_conc_844_18_7 , (~ (data_rsci_idat[420:414]))});
  assign MultLoop_acc_1065_nl = nl_MultLoop_acc_1065_nl[25:0];
  assign nl_MultLoop_acc_1624_nl = (~ (data_rsci_idat[341:324])) + conv_s2s_15_18(data_rsci_idat[341:327]);
  assign MultLoop_acc_1624_nl = nl_MultLoop_acc_1624_nl[17:0];
  assign nl_MultLoop_acc_1625_nl = ({(data_rsci_idat[341:324]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1624_nl);
  assign MultLoop_acc_1625_nl = nl_MultLoop_acc_1625_nl[19:0];
  assign nl_MultLoop_acc_1438_nl = conv_s2u_20_23(MultLoop_acc_1625_nl) + conv_s2u_22_23({(data_rsci_idat[341:324])
      , 4'b0000});
  assign MultLoop_acc_1438_nl = nl_MultLoop_acc_1438_nl[22:0];
  assign nl_MultLoop_acc_1437_nl = conv_s2u_18_20(MultLoop_acc_1626_cse_1) + ({(data_rsci_idat[287:270])
      , 2'b01});
  assign MultLoop_acc_1437_nl = nl_MultLoop_acc_1437_nl[19:0];
  assign nl_MultLoop_acc_3953_nl = conv_s2s_11_12(data_rsci_idat[143:133]) + 12'b000000000001;
  assign MultLoop_acc_3953_nl = nl_MultLoop_acc_3953_nl[11:0];
  assign nl_MultLoop_acc_1632_nl = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_14_19({(MultLoop_acc_3953_nl)
      , (data_rsci_idat[132:131])});
  assign MultLoop_acc_1632_nl = nl_MultLoop_acc_1632_nl[18:0];
  assign nl_MultLoop_acc_1050_nl = conv_s2u_19_20(MultLoop_acc_1632_nl) + ({(~ (data_rsci_idat[143:126]))
      , 2'b00});
  assign MultLoop_acc_1050_nl = nl_MultLoop_acc_1050_nl[19:0];
  assign nl_MultLoop_acc_1685_itm_1  = conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1434_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1052_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_1065_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1438_nl))) + conv_s2s_16_18(MultLoop_acc_541_itm_23_8)
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1437_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1050_nl)))
      + conv_s2s_16_18(MultLoop_acc_1211_itm_23_8);
  assign nl_MultLoop_acc_3954_nl = conv_s2s_13_14(data_rsci_idat[53:41]) + 14'b00000000000001;
  assign MultLoop_acc_3954_nl = nl_MultLoop_acc_3954_nl[13:0];
  assign nl_MultLoop_acc_1634_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18({(MultLoop_acc_3954_nl)
      , (data_rsci_idat[40:39])});
  assign MultLoop_acc_1634_nl = nl_MultLoop_acc_1634_nl[17:0];
  assign nl_MultLoop_acc_1432_nl = conv_s2u_18_21(MultLoop_acc_1634_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[53:36])) , 2'b01});
  assign MultLoop_acc_1432_nl = nl_MultLoop_acc_1432_nl[20:0];
  assign nl_MultLoop_acc_1637_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1636_cse_1);
  assign MultLoop_acc_1637_nl = nl_MultLoop_acc_1637_nl[19:0];
  assign nl_MultLoop_acc_1046_nl = conv_s2u_20_23(MultLoop_acc_1637_nl) + ({(~ (data_rsci_idat[71:54]))
      , 5'b00000});
  assign MultLoop_acc_1046_nl = nl_MultLoop_acc_1046_nl[22:0];
  assign nl_MultLoop_acc_1677_itm_1  = conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1432_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1046_nl))) + conv_s2s_16_18(MultLoop_acc_1043_cse_1[19:4])
      + conv_s2s_16_18(MultLoop_acc_856_itm_22_7);
  assign nl_Result_acc_164_nl = conv_s2s_21_22({(data_rsci_idat[755:738]) , 3'b000})
      + conv_s2s_19_22(Result_acc_163_cse_1);
  assign Result_acc_164_nl = nl_Result_acc_164_nl[21:0];
  assign nl_Result_acc_10_nl = conv_s2u_22_23(Result_acc_164_nl) + ({(~ (data_rsci_idat[755:738]))
      , 5'b00000});
  assign Result_acc_10_nl = nl_Result_acc_10_nl[22:0];
  assign nl_Result_acc_215_nl = conv_s2s_14_15(data_rsci_idat[827:814]) + 15'b000000000000001;
  assign Result_acc_215_nl = nl_Result_acc_215_nl[14:0];
  assign nl_Result_acc_166_nl = conv_s2s_18_19(data_rsci_idat[827:810]) + conv_s2s_17_19({(Result_acc_215_nl)
      , (data_rsci_idat[813:812])});
  assign Result_acc_166_nl = nl_Result_acc_166_nl[18:0];
  assign nl_Result_acc_14_nl = conv_s2u_19_20(Result_acc_166_nl) + ({(~ (data_rsci_idat[827:810]))
      , 2'b00});
  assign Result_acc_14_nl = nl_Result_acc_14_nl[19:0];
  assign nl_Result_acc_169_nl = conv_s2s_21_22({(data_rsci_idat[845:828]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[845:828]) + conv_s2s_17_22({Result_acc_216_cse_1
      , (data_rsci_idat[834:830])});
  assign Result_acc_169_nl = nl_Result_acc_169_nl[21:0];
  assign nl_Result_acc_15_nl = conv_s2u_22_23(Result_acc_169_nl) + ({(~ (data_rsci_idat[845:828]))
      , 5'b00000});
  assign Result_acc_15_nl = nl_Result_acc_15_nl[22:0];
  assign nl_MultLoop_acc_1676_itm_1  = conv_s2s_16_18(readslicef_23_16_7((Result_acc_10_nl)))
      + conv_s2s_16_18(MultLoop_acc_3930_itm_17_2) + conv_s2s_16_18(readslicef_20_16_4((Result_acc_14_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((Result_acc_15_nl)));
  assign nl_MultLoop_acc_3794_nl = ({(data_rsci_idat[485:468]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_692_18_7
      , (~ (data_rsci_idat[474:468]))});
  assign MultLoop_acc_3794_nl = nl_MultLoop_acc_3794_nl[19:0];
  assign nl_MultLoop_acc_3795_nl = ({(~ (data_rsci_idat[485:468])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3794_nl);
  assign MultLoop_acc_3795_nl = nl_MultLoop_acc_3795_nl[21:0];
  assign nl_MultLoop_acc_74_nl = conv_s2s_22_26(MultLoop_acc_3795_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[485:468])) , 7'b0010000});
  assign MultLoop_acc_74_nl = nl_MultLoop_acc_74_nl[25:0];
  assign nl_MultLoop_acc_4529_nl =  -conv_s2s_14_15(data_rsci_idat[323:310]);
  assign MultLoop_acc_4529_nl = nl_MultLoop_acc_4529_nl[14:0];
  assign nl_MultLoop_acc_66_nl = conv_s2s_19_23({(MultLoop_acc_4529_nl) , (~ (data_rsci_idat[309:306]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[323:306])) , 4'b0001});
  assign MultLoop_acc_66_nl = nl_MultLoop_acc_66_nl[22:0];
  assign nl_MultLoop_acc_4530_nl = conv_s2s_12_13(data_rsci_idat[35:24]) + 13'b0000000000001;
  assign MultLoop_acc_4530_nl = nl_MultLoop_acc_4530_nl[12:0];
  assign nl_MultLoop_acc_3798_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_16_18({(MultLoop_acc_4530_nl)
      , (data_rsci_idat[23:21])});
  assign MultLoop_acc_3798_nl = nl_MultLoop_acc_3798_nl[17:0];
  assign nl_MultLoop_acc_1089_nl = conv_s2u_18_22(MultLoop_acc_3798_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[35:18])) , 3'b001});
  assign MultLoop_acc_1089_nl = nl_MultLoop_acc_1089_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_366_itm_1 
      = conv_s2s_17_18(MultLoop_acc_1095_itm_18_2) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_74_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_66_nl))) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1089_nl)));
  assign nl_MultLoop_acc_3740_nl = (~ (data_rsci_idat[791:774])) + conv_s2s_17_18({MultLoop_MultLoop_conc_740_16_4
      , (data_rsci_idat[779:776])});
  assign MultLoop_acc_3740_nl = nl_MultLoop_acc_3740_nl[17:0];
  assign nl_MultLoop_acc_3741_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3740_nl);
  assign MultLoop_acc_3741_nl = nl_MultLoop_acc_3741_nl[19:0];
  assign nl_MultLoop_acc_90_nl = conv_s2u_20_22(MultLoop_acc_3741_nl) + ({(~ (data_rsci_idat[791:774]))
      , 4'b0000});
  assign MultLoop_acc_90_nl = nl_MultLoop_acc_90_nl[21:0];
  assign nl_MultLoop_acc_4532_nl = conv_s2s_13_14(data_rsci_idat[665:653]) + 14'b00000000000001;
  assign MultLoop_acc_4532_nl = nl_MultLoop_acc_4532_nl[13:0];
  assign nl_MultLoop_acc_3743_nl = conv_s2s_18_19(data_rsci_idat[665:648]) + conv_s2s_17_19({(MultLoop_acc_4532_nl)
      , (data_rsci_idat[652:650])});
  assign MultLoop_acc_3743_nl = nl_MultLoop_acc_3743_nl[18:0];
  assign nl_MultLoop_acc_84_nl = conv_s2u_19_21(MultLoop_acc_3743_nl) + ({(~ (data_rsci_idat[665:648]))
      , 3'b000});
  assign MultLoop_acc_84_nl = nl_MultLoop_acc_84_nl[20:0];
  assign nl_MultLoop_acc_3744_nl = conv_s2s_18_19(data_rsci_idat[233:216]) + conv_s2s_16_19(data_rsci_idat[233:218]);
  assign MultLoop_acc_3744_nl = nl_MultLoop_acc_3744_nl[18:0];
  assign nl_MultLoop_acc_1091_nl = conv_s2u_19_21(MultLoop_acc_3744_nl) + conv_s2u_20_21({(data_rsci_idat[233:216])
      , 2'b00});
  assign MultLoop_acc_1091_nl = nl_MultLoop_acc_1091_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_344_itm_1 
      = conv_s2s_14_16(data_rsci_idat[467:454]) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_90_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_84_nl))) + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1091_nl)));
  assign nl_MultLoop_acc_59_nl = conv_s2u_12_18(data_rsci_idat[197:186]) - (data_rsci_idat[197:180]);
  assign MultLoop_acc_59_nl = nl_MultLoop_acc_59_nl[17:0];
  assign nl_MultLoop_acc_4533_nl = conv_s2s_13_14(data_rsci_idat[215:203]) + 14'b00000000000001;
  assign MultLoop_acc_4533_nl = nl_MultLoop_acc_4533_nl[13:0];
  assign nl_MultLoop_acc_3746_nl = conv_s2s_18_19(data_rsci_idat[215:198]) + conv_s2s_16_19({(MultLoop_acc_4533_nl)
      , (data_rsci_idat[202:201])});
  assign MultLoop_acc_3746_nl = nl_MultLoop_acc_3746_nl[18:0];
  assign nl_MultLoop_acc_60_nl = conv_s2u_19_20(MultLoop_acc_3746_nl) + ({(~ (data_rsci_idat[215:198]))
      , 2'b00});
  assign MultLoop_acc_60_nl = nl_MultLoop_acc_60_nl[19:0];
  assign nl_MultLoop_acc_1090_nl = conv_s2u_18_22(MultLoop_acc_2685_cse_1) + ({(data_rsci_idat[125:108])
      , 4'b0001});
  assign MultLoop_acc_1090_nl = nl_MultLoop_acc_1090_nl[21:0];
  assign nl_MultLoop_acc_4534_nl =  -conv_s2s_12_13(data_rsci_idat[89:78]);
  assign MultLoop_acc_4534_nl = nl_MultLoop_acc_4534_nl[12:0];
  assign nl_MultLoop_acc_3749_nl = ({(data_rsci_idat[89:72]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_4534_nl)
      , (~ (data_rsci_idat[77:72]))});
  assign MultLoop_acc_3749_nl = nl_MultLoop_acc_3749_nl[21:0];
  assign nl_MultLoop_acc_4535_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3749_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_4535_nl = nl_MultLoop_acc_4535_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_343_itm_1 
      = conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_59_nl))) + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_60_nl)))
      + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_1090_nl))) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4535_nl)));
  assign nl_MultLoop_acc_1099_nl = conv_s2u_18_22(MultLoop_acc_2307_cse_1) + ({(data_rsci_idat[773:756])
      , 4'b0001});
  assign MultLoop_acc_1099_nl = nl_MultLoop_acc_1099_nl[21:0];
  assign nl_MultLoop_acc_52_nl = conv_s2s_18_22(~ (data_rsci_idat[71:54])) + ({(data_rsci_idat[71:54])
      , 4'b0001});
  assign MultLoop_acc_52_nl = nl_MultLoop_acc_52_nl[21:0];
  assign nl_MultLoop_acc_4536_nl =  -conv_s2s_16_17(data_rsci_idat[377:362]);
  assign MultLoop_acc_4536_nl = nl_MultLoop_acc_4536_nl[16:0];
  assign nl_MultLoop_acc_69_nl = conv_s2s_19_21({(MultLoop_acc_4536_nl) , (~ (data_rsci_idat[361:360]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[377:360])) , 2'b01});
  assign MultLoop_acc_69_nl = nl_MultLoop_acc_69_nl[20:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl = ~((data_rsci_idat[727:720]!=8'b00000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl = (readslicef_21_12_9((MultLoop_acc_69_nl)))
      + conv_s2s_10_12(~ (data_rsci_idat[737:728])) + conv_u2s_1_12(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl[11:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_342_itm_1 
      = conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_1099_nl))) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_52_nl)))
      + conv_s2s_12_16(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_327_nl)
      + conv_s2s_12_16(MultLoop_acc_3182_cse_1[19:8]);
  assign nl_MultLoop_acc_4537_nl =  -conv_s2s_12_13(data_rsci_idat[683:672]);
  assign MultLoop_acc_4537_nl = nl_MultLoop_acc_4537_nl[12:0];
  assign nl_MultLoop_acc_3752_nl = ({(data_rsci_idat[683:666]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4537_nl)
      , (~ (data_rsci_idat[671:666]))});
  assign MultLoop_acc_3752_nl = nl_MultLoop_acc_3752_nl[19:0];
  assign nl_MultLoop_acc_3753_nl = ({(~ (data_rsci_idat[683:666])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3752_nl);
  assign MultLoop_acc_3753_nl = nl_MultLoop_acc_3753_nl[21:0];
  assign nl_MultLoop_acc_85_nl = conv_s2s_22_25(MultLoop_acc_3753_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[683:666])) , 6'b010000});
  assign MultLoop_acc_85_nl = nl_MultLoop_acc_85_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_341_itm_1 
      = conv_s2s_15_16(MultLoop_acc_87_itm_19_4[15:1]) + conv_s2s_15_16(readslicef_25_15_10((MultLoop_acc_85_nl)));
  assign nl_MultLoop_acc_3755_nl = ({(data_rsci_idat[449:432]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_806_18_5
      , (~ (data_rsci_idat[436:432]))});
  assign MultLoop_acc_3755_nl = nl_MultLoop_acc_3755_nl[20:0];
  assign nl_MultLoop_acc_73_nl = conv_s2s_21_23(MultLoop_acc_3755_nl) + ({(~ (data_rsci_idat[449:432]))
      , 5'b00000});
  assign MultLoop_acc_73_nl = nl_MultLoop_acc_73_nl[22:0];
  assign nl_MultLoop_acc_3756_nl = conv_s2s_21_22({(~ (data_rsci_idat[413:396]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[413:396]));
  assign MultLoop_acc_3756_nl = nl_MultLoop_acc_3756_nl[21:0];
  assign nl_MultLoop_acc_71_nl = conv_s2s_22_25(MultLoop_acc_3756_nl) + ({(data_rsci_idat[413:396])
      , 7'b0001000});
  assign MultLoop_acc_71_nl = nl_MultLoop_acc_71_nl[24:0];
  assign nl_MultLoop_acc_4539_nl =  -conv_s2s_12_13(data_rsci_idat[305:294]);
  assign MultLoop_acc_4539_nl = nl_MultLoop_acc_4539_nl[12:0];
  assign nl_MultLoop_acc_3758_nl = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4539_nl)
      , (~ (data_rsci_idat[293:288]))});
  assign MultLoop_acc_3758_nl = nl_MultLoop_acc_3758_nl[19:0];
  assign nl_MultLoop_acc_3759_nl = ({(~ (data_rsci_idat[305:288])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3758_nl);
  assign MultLoop_acc_3759_nl = nl_MultLoop_acc_3759_nl[21:0];
  assign nl_MultLoop_acc_65_nl = conv_s2s_22_25(MultLoop_acc_3759_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[305:288])) , 6'b010000});
  assign MultLoop_acc_65_nl = nl_MultLoop_acc_65_nl[24:0];
  assign nl_MultLoop_acc_4655_nl = conv_s2u_17_19(MultLoop_acc_2057_cse_1[18:2])
      + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_4655_nl = nl_MultLoop_acc_4655_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_354_itm_1 
      = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_73_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_71_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_65_nl))) + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4655_nl)));
  assign nl_MultLoop_acc_4656_nl = conv_s2u_14_19(MultLoop_acc_3761_itm_19_6) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_4656_nl = nl_MultLoop_acc_4656_nl[18:0];
  assign nl_MultLoop_acc_88_nl = conv_s2s_18_22(~ (data_rsci_idat[755:738])) + ({(data_rsci_idat[755:738])
      , 4'b0001});
  assign MultLoop_acc_88_nl = nl_MultLoop_acc_88_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl = conv_s2s_13_14(readslicef_22_13_9((MultLoop_acc_88_nl)))
      + conv_s2s_13_14(MultLoop_acc_1097_itm_18_4[14:2]);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl[13:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl = (readslicef_19_15_4((MultLoop_acc_4656_nl)))
      + conv_s2s_14_15(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_331_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl[14:0];
  assign nl_MultLoop_acc_3763_nl = conv_s2s_23_24({(~ (data_rsci_idat[845:828]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[845:828])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[845:828]));
  assign MultLoop_acc_3763_nl = nl_MultLoop_acc_3763_nl[23:0];
  assign nl_MultLoop_acc_93_nl = conv_s2s_24_25(MultLoop_acc_3763_nl) + ({(data_rsci_idat[845:828])
      , 7'b0100000});
  assign MultLoop_acc_93_nl = nl_MultLoop_acc_93_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_353_itm_1 
      = conv_s2s_15_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_338_nl)
      + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_93_nl)));
  assign nl_MultLoop_acc_4540_nl = conv_s2s_11_12(data_rsci_idat[827:817]) + 12'b000000000001;
  assign MultLoop_acc_4540_nl = nl_MultLoop_acc_4540_nl[11:0];
  assign nl_MultLoop_acc_3766_nl = conv_s2s_21_22({(data_rsci_idat[827:810]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[827:810]) + conv_s2s_17_22({(MultLoop_acc_4540_nl)
      , (data_rsci_idat[816:812])});
  assign MultLoop_acc_3766_nl = nl_MultLoop_acc_3766_nl[21:0];
  assign nl_MultLoop_acc_92_nl = conv_s2u_22_23(MultLoop_acc_3766_nl) + ({(~ (data_rsci_idat[827:810]))
      , 5'b00000});
  assign MultLoop_acc_92_nl = nl_MultLoop_acc_92_nl[22:0];
  assign nl_MultLoop_acc_3769_nl = ({(data_rsci_idat[701:684]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[701:684])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_828_18_7
      , (~ (data_rsci_idat[690:684]))});
  assign MultLoop_acc_3769_nl = nl_MultLoop_acc_3769_nl[22:0];
  assign nl_MultLoop_acc_4542_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3769_nl)))
      + (~ (data_rsci_idat[701:684]));
  assign MultLoop_acc_4542_nl = nl_MultLoop_acc_4542_nl[17:0];
  assign nl_MultLoop_acc_82_nl = conv_s2s_18_20(~ (data_rsci_idat[629:612])) + ({(data_rsci_idat[629:612])
      , 2'b01});
  assign MultLoop_acc_82_nl = nl_MultLoop_acc_82_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_363_itm_1 
      = conv_s2s_16_18(MultLoop_acc_3636_cse_1[19:4]) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_92_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4542_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_82_nl)));
  assign nl_MultLoop_acc_83_nl = conv_s2s_24_25({(~ (data_rsci_idat[647:630])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[647:630])) , 3'b001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_754_18_6
      , (~ (data_rsci_idat[635:630]))});
  assign MultLoop_acc_83_nl = nl_MultLoop_acc_83_nl[24:0];
  assign nl_MultLoop_acc_3774_nl = conv_s2s_22_23({(data_rsci_idat[539:522]) , 4'b0000})
      + conv_s2s_18_23(data_rsci_idat[539:522]) + conv_s2s_17_23({MultLoop_acc_4167_cse_1
      , (data_rsci_idat[529:524])});
  assign MultLoop_acc_3774_nl = nl_MultLoop_acc_3774_nl[22:0];
  assign nl_MultLoop_acc_4545_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3774_nl)))
      + (~ (data_rsci_idat[539:522]));
  assign MultLoop_acc_4545_nl = nl_MultLoop_acc_4545_nl[17:0];
  assign nl_MultLoop_acc_4657_nl = conv_s2u_18_19(data_rsci_idat[503:486]) + conv_s2u_16_19(MultLoop_acc_2317_itm_20_5);
  assign MultLoop_acc_4657_nl = nl_MultLoop_acc_4657_nl[18:0];
  assign nl_MultLoop_acc_4546_nl = conv_s2u_17_19(readslicef_19_17_2((MultLoop_acc_4657_nl)))
      + conv_s2u_18_19(data_rsci_idat[503:486]);
  assign MultLoop_acc_4546_nl = nl_MultLoop_acc_4546_nl[18:0];
  assign nl_MultLoop_acc_3779_nl = conv_s2s_20_21({(data_rsci_idat[431:414]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_2584_cse_1);
  assign MultLoop_acc_3779_nl = nl_MultLoop_acc_3779_nl[20:0];
  assign nl_MultLoop_acc_72_nl = conv_s2u_21_23(MultLoop_acc_3779_nl) + ({(~ (data_rsci_idat[431:414]))
      , 5'b00000});
  assign MultLoop_acc_72_nl = nl_MultLoop_acc_72_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_362_itm_1 
      = conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_83_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4545_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4546_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_72_nl)));
  assign nl_MultLoop_acc_4548_nl = conv_s2s_13_14(data_rsci_idat[359:347]) + 14'b00000000000001;
  assign MultLoop_acc_4548_nl = nl_MultLoop_acc_4548_nl[13:0];
  assign nl_MultLoop_acc_3781_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_17_18({(MultLoop_acc_4548_nl)
      , (data_rsci_idat[346:344])});
  assign MultLoop_acc_3781_nl = nl_MultLoop_acc_3781_nl[17:0];
  assign nl_MultLoop_acc_1094_nl = conv_s2u_18_22(MultLoop_acc_3781_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[359:342])) , 3'b001});
  assign MultLoop_acc_1094_nl = nl_MultLoop_acc_1094_nl[21:0];
  assign nl_MultLoop_acc_3783_nl = ({(data_rsci_idat[251:234]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_770_18_8
      , (~ (data_rsci_idat[241:234]))});
  assign MultLoop_acc_3783_nl = nl_MultLoop_acc_3783_nl[19:0];
  assign nl_MultLoop_acc_4550_nl = conv_s2u_12_18(readslicef_20_12_8((MultLoop_acc_3783_nl)))
      + (~ (data_rsci_idat[251:234]));
  assign MultLoop_acc_4550_nl = nl_MultLoop_acc_4550_nl[17:0];
  assign nl_MultLoop_acc_4551_nl =  -conv_s2s_10_11(data_rsci_idat[161:152]);
  assign MultLoop_acc_4551_nl = nl_MultLoop_acc_4551_nl[10:0];
  assign nl_MultLoop_acc_3785_nl = ({(data_rsci_idat[161:144]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4551_nl)
      , (~ (data_rsci_idat[151:144]))});
  assign MultLoop_acc_3785_nl = nl_MultLoop_acc_3785_nl[20:0];
  assign nl_MultLoop_acc_3786_nl = conv_s2s_23_24({(data_rsci_idat[161:144]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_3785_nl);
  assign MultLoop_acc_3786_nl = nl_MultLoop_acc_3786_nl[23:0];
  assign nl_MultLoop_acc_4552_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3786_nl)))
      + (~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_4552_nl = nl_MultLoop_acc_4552_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_361_itm_1 
      = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1094_nl))) + conv_s2s_16_18(MultLoop_acc_1611_cse_1[18:3])
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4550_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4552_nl)));
  assign nl_MultLoop_acc_3792_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_17_18({MultLoop_acc_4212_cse_1
      , (data_rsci_idat[565:560])});
  assign MultLoop_acc_3792_nl = nl_MultLoop_acc_3792_nl[17:0];
  assign nl_MultLoop_acc_1096_nl = conv_s2u_18_25(MultLoop_acc_3792_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[575:558])) , 6'b000001});
  assign MultLoop_acc_1096_nl = nl_MultLoop_acc_1096_nl[24:0];
  assign nl_MultLoop_acc_3788_nl = ({(data_rsci_idat[143:126]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_848_18_7
      , (~ (data_rsci_idat[132:126]))});
  assign MultLoop_acc_3788_nl = nl_MultLoop_acc_3788_nl[21:0];
  assign nl_MultLoop_acc_4554_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_3788_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_4554_nl = nl_MultLoop_acc_4554_nl[17:0];
  assign nl_MultLoop_acc_4555_nl =  -conv_s2s_13_14(data_rsci_idat[53:41]);
  assign MultLoop_acc_4555_nl = nl_MultLoop_acc_4555_nl[13:0];
  assign nl_MultLoop_acc_51_nl = conv_s2s_23_24({(~ (data_rsci_idat[53:36])) , 5'b00100})
      + conv_s2s_20_24({(~ (data_rsci_idat[53:36])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4555_nl)
      , (~ (data_rsci_idat[40:36]))});
  assign MultLoop_acc_51_nl = nl_MultLoop_acc_51_nl[23:0];
  assign nl_MultLoop_acc_49_nl = conv_s2u_14_18(data_rsci_idat[17:4]) - (data_rsci_idat[17:0]);
  assign MultLoop_acc_49_nl = nl_MultLoop_acc_49_nl[17:0];
  assign nl_MultLoop_49_MultLoop_acc_3_nl = (readslicef_18_16_2((MultLoop_acc_49_nl)))
      + 16'b0000001000010111;
  assign MultLoop_49_MultLoop_acc_3_nl = nl_MultLoop_49_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_78_nl = conv_s2s_18_23(~ (data_rsci_idat[557:540])) + ({(data_rsci_idat[557:540])
      , 5'b00001});
  assign MultLoop_acc_78_nl = nl_MultLoop_acc_78_nl[22:0];
  assign nl_MultLoop_acc_70_nl = conv_s2s_18_21(~ (data_rsci_idat[395:378])) + ({(data_rsci_idat[395:378])
      , 3'b001});
  assign MultLoop_acc_70_nl = nl_MultLoop_acc_70_nl[20:0];
  assign nl_MultLoop_acc_4556_nl =  -conv_s2s_14_15(data_rsci_idat[179:166]);
  assign MultLoop_acc_4556_nl = nl_MultLoop_acc_4556_nl[14:0];
  assign nl_MultLoop_acc_3738_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4556_nl)
      , (~ (data_rsci_idat[165:162]))});
  assign MultLoop_acc_3738_nl = nl_MultLoop_acc_3738_nl[19:0];
  assign nl_MultLoop_acc_58_nl = conv_s2s_20_22(MultLoop_acc_3738_nl) + ({(~ (data_rsci_idat[179:162]))
      , 4'b0000});
  assign MultLoop_acc_58_nl = nl_MultLoop_acc_58_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_367_itm_1 
      = conv_s2s_17_18(MultLoop_acc_4588_itm_18_2) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1096_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4554_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_51_nl)))
      + conv_s2s_16_18(MultLoop_49_MultLoop_acc_3_nl) + conv_s2s_13_18(readslicef_23_13_10((MultLoop_acc_78_nl)))
      + conv_s2s_13_18(readslicef_21_13_8((MultLoop_acc_70_nl))) + conv_s2s_13_18(MultLoop_acc_67_itm_17_3[14:2])
      + conv_s2s_13_18(readslicef_22_13_9((MultLoop_acc_58_nl)));
  assign nl_MultLoop_acc_1749_nl = ({(data_rsci_idat[323:306]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[323:306])) , 3'b001}) + conv_s2s_18_23(~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_1749_nl = nl_MultLoop_acc_1749_nl[22:0];
  assign nl_MultLoop_acc_3958_nl = conv_s2u_15_19(readslicef_23_15_8((MultLoop_acc_1749_nl)))
      + conv_s2u_18_19(data_rsci_idat[323:306]);
  assign MultLoop_acc_3958_nl = nl_MultLoop_acc_3958_nl[18:0];
  assign nl_MultLoop_acc_1750_nl = ({(data_rsci_idat[287:270]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[287:270]));
  assign MultLoop_acc_1750_nl = nl_MultLoop_acc_1750_nl[21:0];
  assign nl_MultLoop_acc_3959_nl = conv_s2u_14_19(readslicef_22_14_8((MultLoop_acc_1750_nl)))
      + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_3959_nl = nl_MultLoop_acc_3959_nl[18:0];
  assign nl_MultLoop_acc_1752_nl = conv_s2s_24_25({(~ (data_rsci_idat[161:144]))
      , 6'b010000}) + conv_s2s_23_25(MultLoop_acc_4690);
  assign MultLoop_acc_1752_nl = nl_MultLoop_acc_1752_nl[24:0];
  assign nl_MultLoop_acc_1004_nl = conv_s2s_25_27(MultLoop_acc_1752_nl) + ({(data_rsci_idat[161:144])
      , 9'b001000000});
  assign MultLoop_acc_1004_nl = nl_MultLoop_acc_1004_nl[26:0];
  assign nl_MultLoop_acc_4596_nl = conv_s2u_18_19(data_rsci_idat[53:36]) + conv_s2u_17_19(MultLoop_acc_4594_itm_18_2);
  assign MultLoop_acc_4596_nl = nl_MultLoop_acc_4596_nl[18:0];
  assign nl_MultLoop_acc_3960_nl = conv_s2u_17_19(readslicef_19_17_2((MultLoop_acc_4596_nl)))
      + conv_s2u_18_19(data_rsci_idat[53:36]);
  assign MultLoop_acc_3960_nl = nl_MultLoop_acc_3960_nl[18:0];
  assign nl_MultLoop_acc_1795_nl = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_3958_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_3959_nl))) + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_1004_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_3960_nl)));
  assign MultLoop_acc_1795_nl = nl_MultLoop_acc_1795_nl[17:0];
  assign nl_MultLoop_acc_1430_nl = conv_s2u_10_19(data_rsci_idat[737:728]) + conv_s2u_18_19(data_rsci_idat[737:720]);
  assign MultLoop_acc_1430_nl = nl_MultLoop_acc_1430_nl[18:0];
  assign nl_MultLoop_acc_4595_nl = conv_s2u_15_19(MultLoop_acc_1743_cse_1[20:6])
      + conv_s2u_18_19(data_rsci_idat[665:648]);
  assign MultLoop_acc_4595_nl = nl_MultLoop_acc_4595_nl[18:0];
  assign nl_MultLoop_acc_3956_nl = (~ (data_rsci_idat[449:432])) + conv_s2s_13_18(MultLoop_acc_4692[19:7]);
  assign MultLoop_acc_3956_nl = nl_MultLoop_acc_3956_nl[17:0];
  assign nl_MultLoop_acc_3957_nl = conv_s2u_18_20(MultLoop_acc_3956_nl) + ({(data_rsci_idat[449:432])
      , 2'b01});
  assign MultLoop_acc_3957_nl = nl_MultLoop_acc_3957_nl[19:0];
  assign nl_MultLoop_acc_1746_nl = (~ (data_rsci_idat[413:396])) + conv_s2s_15_18(data_rsci_idat[413:399]);
  assign MultLoop_acc_1746_nl = nl_MultLoop_acc_1746_nl[17:0];
  assign nl_MultLoop_acc_1747_nl = ({(data_rsci_idat[413:396]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1746_nl);
  assign MultLoop_acc_1747_nl = nl_MultLoop_acc_1747_nl[19:0];
  assign nl_MultLoop_acc_1422_nl = conv_s2u_20_24(MultLoop_acc_1747_nl) + conv_s2u_23_24({(data_rsci_idat[413:396])
      , 5'b00000});
  assign MultLoop_acc_1422_nl = nl_MultLoop_acc_1422_nl[23:0];
  assign nl_MultLoop_acc_1800_itm_1  = (MultLoop_acc_1795_nl) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_1430_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4595_nl))) + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_3957_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1422_nl)));
  assign nl_MultLoop_acc_1695_nl = (~ (data_rsci_idat[863:846])) + conv_s2s_17_18({MultLoop_acc_3961_cse_1
      , (data_rsci_idat[851:848])});
  assign MultLoop_acc_1695_nl = nl_MultLoop_acc_1695_nl[17:0];
  assign nl_MultLoop_acc_1696_nl = ({(data_rsci_idat[863:846]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1695_nl);
  assign MultLoop_acc_1696_nl = nl_MultLoop_acc_1696_nl[19:0];
  assign nl_MultLoop_acc_1042_nl = conv_s2u_20_22(MultLoop_acc_1696_nl) + ({(~ (data_rsci_idat[863:846]))
      , 4'b0000});
  assign MultLoop_acc_1042_nl = nl_MultLoop_acc_1042_nl[21:0];
  assign nl_MultLoop_acc_1431_nl = conv_s2u_16_19(data_rsci_idat[827:812]) + conv_s2u_18_19(data_rsci_idat[827:810]);
  assign MultLoop_acc_1431_nl = nl_MultLoop_acc_1431_nl[18:0];
  assign nl_MultLoop_acc_1698_nl = ({(data_rsci_idat[755:738]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_842_18_6
      , (~ (data_rsci_idat[743:738]))});
  assign MultLoop_acc_1698_nl = nl_MultLoop_acc_1698_nl[21:0];
  assign nl_MultLoop_acc_3963_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_1698_nl)))
      + (~ (data_rsci_idat[755:738]));
  assign MultLoop_acc_3963_nl = nl_MultLoop_acc_3963_nl[17:0];
  assign nl_MultLoop_acc_1002_nl = conv_s2s_18_22(~ (data_rsci_idat[125:108])) +
      ({(data_rsci_idat[125:108]) , 4'b0001});
  assign MultLoop_acc_1002_nl = nl_MultLoop_acc_1002_nl[21:0];
  assign nl_MultLoop_acc_1756_nl = conv_s2s_9_10(data_rsci_idat[269:261]) + 10'b0000111111;
  assign MultLoop_acc_1756_nl = nl_MultLoop_acc_1756_nl[9:0];
  assign nl_MultLoop_acc_1772_itm_1  = conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_1042_nl)))
      + conv_s2s_14_16(readslicef_19_14_5((MultLoop_acc_1431_nl))) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_3963_nl)))
      + conv_s2s_13_16(readslicef_22_13_9((MultLoop_acc_1002_nl))) + conv_s2s_10_16(MultLoop_acc_1756_nl);
  assign nl_MultLoop_acc_3964_nl = conv_s2s_14_15(data_rsci_idat[521:508]) + 15'b000000000000001;
  assign MultLoop_acc_3964_nl = nl_MultLoop_acc_3964_nl[14:0];
  assign nl_MultLoop_acc_1701_nl = (~ (data_rsci_idat[521:504])) + conv_s2s_17_18({(MultLoop_acc_3964_nl)
      , (data_rsci_idat[507:506])});
  assign MultLoop_acc_1701_nl = nl_MultLoop_acc_1701_nl[17:0];
  assign nl_MultLoop_acc_1423_nl = conv_s2u_18_21(MultLoop_acc_1701_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[521:504])) , 2'b01});
  assign MultLoop_acc_1423_nl = nl_MultLoop_acc_1423_nl[20:0];
  assign nl_MultLoop_acc_4597_nl = conv_s2u_19_20(MultLoop_acc_1702_cse_1[20:2])
      + ({(data_rsci_idat[431:414]) , 2'b01});
  assign MultLoop_acc_4597_nl = nl_MultLoop_acc_4597_nl[19:0];
  assign nl_MultLoop_acc_1771_itm_1  = conv_s2s_14_16(MultLoop_acc_4591_itm_18_2[16:3])
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1423_nl))) + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_4597_nl)))
      + conv_s2s_14_16(MultLoop_acc_355_itm_20_6[14:1]);
  assign nl_MultLoop_acc_1706_nl = ({(data_rsci_idat[809:792]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[809:792])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_858_18_7
      , (~ (data_rsci_idat[798:792]))});
  assign MultLoop_acc_1706_nl = nl_MultLoop_acc_1706_nl[22:0];
  assign nl_MultLoop_acc_3966_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_1706_nl)))
      + (~ (data_rsci_idat[809:792]));
  assign MultLoop_acc_3966_nl = nl_MultLoop_acc_3966_nl[17:0];
  assign nl_MultLoop_acc_1707_nl = conv_s2s_18_19(data_rsci_idat[719:702]) + conv_s2s_15_19(data_rsci_idat[719:705]);
  assign MultLoop_acc_1707_nl = nl_MultLoop_acc_1707_nl[18:0];
  assign nl_MultLoop_acc_1429_nl = conv_s2u_19_21(MultLoop_acc_1707_nl) + conv_s2u_20_21({(data_rsci_idat[719:702])
      , 2'b00});
  assign MultLoop_acc_1429_nl = nl_MultLoop_acc_1429_nl[20:0];
  assign nl_MultLoop_acc_1709_nl = conv_s2s_20_21({(data_rsci_idat[629:612]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_1708_cse_1);
  assign MultLoop_acc_1709_nl = nl_MultLoop_acc_1709_nl[20:0];
  assign nl_MultLoop_acc_1427_nl = conv_s2u_21_23(MultLoop_acc_1709_nl) + conv_s2u_22_23({(data_rsci_idat[629:612])
      , 4'b0000});
  assign MultLoop_acc_1427_nl = nl_MultLoop_acc_1427_nl[22:0];
  assign nl_MultLoop_acc_1703_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_15_18(data_rsci_idat[71:57]);
  assign MultLoop_acc_1703_nl = nl_MultLoop_acc_1703_nl[17:0];
  assign nl_MultLoop_acc_1418_nl = conv_s2u_18_20(MultLoop_acc_1703_nl) + ({(data_rsci_idat[71:54])
      , 2'b01});
  assign MultLoop_acc_1418_nl = nl_MultLoop_acc_1418_nl[19:0];
  assign nl_MultLoop_acc_1783_itm_1  = conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_3966_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1429_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1427_nl)))
      + conv_s2s_14_17(MultLoop_acc_1243_itm_19_6) + conv_s2s_14_17(readslicef_20_14_6((MultLoop_acc_1418_nl)));
  assign nl_MultLoop_acc_1027_nl = conv_s2s_24_25({(~ (data_rsci_idat[593:576]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[593:576])) , 4'b0001}) +
      conv_s2s_19_25({MultLoop_MultLoop_conc_704_18_6 , (~ (data_rsci_idat[581:576]))});
  assign MultLoop_acc_1027_nl = nl_MultLoop_acc_1027_nl[24:0];
  assign nl_MultLoop_acc_1712_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_15_18(data_rsci_idat[611:597]);
  assign MultLoop_acc_1712_nl = nl_MultLoop_acc_1712_nl[17:0];
  assign nl_MultLoop_acc_1426_nl = conv_s2u_18_21(MultLoop_acc_1712_nl) + ({(data_rsci_idat[611:594])
      , 3'b001});
  assign MultLoop_acc_1426_nl = nl_MultLoop_acc_1426_nl[20:0];
  assign nl_MultLoop_acc_3968_nl = conv_s2s_12_13(data_rsci_idat[557:546]) + 13'b0000000000001;
  assign MultLoop_acc_3968_nl = nl_MultLoop_acc_3968_nl[12:0];
  assign nl_MultLoop_acc_1714_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_16_18({(MultLoop_acc_3968_nl)
      , (data_rsci_idat[545:543])});
  assign MultLoop_acc_1714_nl = nl_MultLoop_acc_1714_nl[17:0];
  assign nl_MultLoop_acc_1424_nl = conv_s2u_18_22(MultLoop_acc_1714_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[557:540])) , 3'b001});
  assign MultLoop_acc_1424_nl = nl_MultLoop_acc_1424_nl[21:0];
  assign nl_MultLoop_acc_1782_itm_1  = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1027_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1426_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1424_nl)))
      + conv_s2s_15_17(MultLoop_acc_4663_itm_19_4[15:1]);
  assign nl_MultLoop_acc_3969_nl =  -conv_s2s_14_15(data_rsci_idat[503:490]);
  assign MultLoop_acc_3969_nl = nl_MultLoop_acc_3969_nl[14:0];
  assign nl_MultLoop_acc_1022_nl = conv_s2s_19_23({(MultLoop_acc_3969_nl) , (~ (data_rsci_idat[489:486]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[503:486])) , 4'b0001});
  assign MultLoop_acc_1022_nl = nl_MultLoop_acc_1022_nl[22:0];
  assign nl_MultLoop_acc_3970_nl =  -conv_s2s_12_13(data_rsci_idat[467:456]);
  assign MultLoop_acc_3970_nl = nl_MultLoop_acc_3970_nl[12:0];
  assign nl_MultLoop_acc_1020_nl = conv_s2s_24_25({(~ (data_rsci_idat[467:450]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[467:450])) , 4'b0001}) +
      conv_s2s_19_25({(MultLoop_acc_3970_nl) , (~ (data_rsci_idat[455:450]))});
  assign MultLoop_acc_1020_nl = nl_MultLoop_acc_1020_nl[24:0];
  assign nl_MultLoop_acc_1719_nl = conv_s2s_18_19(data_rsci_idat[197:180]) + conv_s2s_15_19(data_rsci_idat[197:183]);
  assign MultLoop_acc_1719_nl = nl_MultLoop_acc_1719_nl[18:0];
  assign nl_MultLoop_acc_1419_nl = conv_s2u_19_22(MultLoop_acc_1719_nl) + conv_s2u_21_22({(data_rsci_idat[197:180])
      , 3'b000});
  assign MultLoop_acc_1419_nl = nl_MultLoop_acc_1419_nl[21:0];
  assign nl_MultLoop_acc_1721_nl = ({(~ (data_rsci_idat[143:126])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_1720_cse_1);
  assign MultLoop_acc_1721_nl = nl_MultLoop_acc_1721_nl[22:0];
  assign nl_MultLoop_acc_1003_nl = conv_s2s_23_25(MultLoop_acc_1721_nl) + ({(data_rsci_idat[143:126])
      , 7'b0100000});
  assign MultLoop_acc_1003_nl = nl_MultLoop_acc_1003_nl[24:0];
  assign nl_MultLoop_acc_1781_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1022_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1020_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1419_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_1003_nl)));
  assign nl_MultLoop_acc_4598_nl = conv_s2u_19_21(MultLoop_acc_1722_cse_1[20:2])
      + ({(data_rsci_idat[17:0]) , 3'b001});
  assign MultLoop_acc_4598_nl = nl_MultLoop_acc_4598_nl[20:0];
  assign nl_MultLoop_acc_1038_nl = conv_s2s_22_23({(~ (data_rsci_idat[791:774]))
      , 4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[791:774])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_738_18_4
      , (~ (data_rsci_idat[777:774]))});
  assign MultLoop_acc_1038_nl = nl_MultLoop_acc_1038_nl[22:0];
  assign nl_MultLoop_acc_3972_nl = conv_s2s_13_14(data_rsci_idat[341:329]) + 14'b00000000000001;
  assign MultLoop_acc_3972_nl = nl_MultLoop_acc_3972_nl[13:0];
  assign nl_MultLoop_acc_1693_nl = conv_s2s_18_19(data_rsci_idat[341:324]) + conv_s2s_17_19({(MultLoop_acc_3972_nl)
      , (data_rsci_idat[328:326])});
  assign MultLoop_acc_1693_nl = nl_MultLoop_acc_1693_nl[18:0];
  assign nl_MultLoop_acc_1013_nl = conv_s2u_19_21(MultLoop_acc_1693_nl) + ({(~ (data_rsci_idat[341:324]))
      , 3'b000});
  assign MultLoop_acc_1013_nl = nl_MultLoop_acc_1013_nl[20:0];
  assign nl_MultLoop_acc_1780_itm_1  = conv_s2s_16_17(MultLoop_acc_4590_itm_20_5)
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_4598_nl))) + conv_s2s_13_17(readslicef_23_13_10((MultLoop_acc_1038_nl)))
      + conv_s2s_13_17(readslicef_21_13_8((MultLoop_acc_1013_nl)));
  assign nl_MultLoop_acc_1724_nl = ({(~ (data_rsci_idat[773:756])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_1723_cse_1);
  assign MultLoop_acc_1724_nl = nl_MultLoop_acc_1724_nl[21:0];
  assign nl_MultLoop_acc_1037_nl = conv_s2s_22_26(MultLoop_acc_1724_nl) + ({(data_rsci_idat[773:756])
      , 8'b00010000});
  assign MultLoop_acc_1037_nl = nl_MultLoop_acc_1037_nl[25:0];
  assign nl_MultLoop_acc_4599_nl = conv_s2u_16_19(Result_acc_154_itm_19_4) + conv_s2u_18_19(data_rsci_idat[683:666]);
  assign MultLoop_acc_4599_nl = nl_MultLoop_acc_4599_nl[18:0];
  assign nl_MultLoop_acc_1779_itm_1  = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_1037_nl)))
      + conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4599_nl)));
  assign nl_MultLoop_acc_1726_nl = conv_s2s_21_22({(~ (data_rsci_idat[647:630]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[647:630]));
  assign MultLoop_acc_1726_nl = nl_MultLoop_acc_1726_nl[21:0];
  assign nl_MultLoop_acc_1030_nl = conv_s2s_22_26(MultLoop_acc_1726_nl) + ({(data_rsci_idat[647:630])
      , 8'b00001000});
  assign MultLoop_acc_1030_nl = nl_MultLoop_acc_1030_nl[25:0];
  assign nl_MultLoop_acc_1728_nl = conv_s2s_20_21({(data_rsci_idat[575:558]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_1727_cse_1);
  assign MultLoop_acc_1728_nl = nl_MultLoop_acc_1728_nl[20:0];
  assign nl_MultLoop_acc_1425_nl = conv_s2u_21_23(MultLoop_acc_1728_nl) + conv_s2u_22_23({(data_rsci_idat[575:558])
      , 4'b0000});
  assign MultLoop_acc_1425_nl = nl_MultLoop_acc_1425_nl[22:0];
  assign nl_MultLoop_acc_1729_nl = conv_s2s_21_22({(~ (data_rsci_idat[539:522]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[539:522]));
  assign MultLoop_acc_1729_nl = nl_MultLoop_acc_1729_nl[21:0];
  assign nl_MultLoop_acc_1024_nl = conv_s2s_22_24(MultLoop_acc_1729_nl) + ({(data_rsci_idat[539:522])
      , 6'b001000});
  assign MultLoop_acc_1024_nl = nl_MultLoop_acc_1024_nl[23:0];
  assign nl_MultLoop_acc_1791_itm_1  = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_1030_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1425_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1024_nl)))
      + conv_s2s_16_18(MultLoop_acc_1350_itm_22_7);
  assign nl_MultLoop_acc_1736_nl = ({(data_rsci_idat[179:162]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[179:162]));
  assign MultLoop_acc_1736_nl = nl_MultLoop_acc_1736_nl[21:0];
  assign nl_MultLoop_acc_3975_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_1736_nl)))
      + conv_s2u_18_19(data_rsci_idat[179:162]);
  assign MultLoop_acc_3975_nl = nl_MultLoop_acc_3975_nl[18:0];
  assign nl_MultLoop_acc_1738_nl = conv_s2s_24_25({(~ (data_rsci_idat[89:72])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[89:72])) , 3'b001}) + conv_s2s_18_25(~
      (data_rsci_idat[89:72]));
  assign MultLoop_acc_1738_nl = nl_MultLoop_acc_1738_nl[24:0];
  assign nl_MultLoop_acc_1000_nl = conv_s2s_25_26(MultLoop_acc_1738_nl) + ({(data_rsci_idat[89:72])
      , 8'b01000000});
  assign MultLoop_acc_1000_nl = nl_MultLoop_acc_1000_nl[25:0];
  assign nl_MultLoop_acc_3973_nl = conv_s2u_16_19(MultLoop_acc_1730_itm_22_7) + conv_s2u_18_19(data_rsci_idat[395:378]);
  assign MultLoop_acc_3973_nl = nl_MultLoop_acc_3973_nl[18:0];
  assign nl_MultLoop_acc_1731_nl = conv_s2s_23_24({(~ (data_rsci_idat[305:288]))
      , 5'b00001}) + conv_s2s_18_24(~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_1731_nl = nl_MultLoop_acc_1731_nl[23:0];
  assign nl_MultLoop_acc_1011_nl = conv_s2s_24_25(MultLoop_acc_1731_nl) + ({(data_rsci_idat[305:288])
      , 7'b0100000});
  assign MultLoop_acc_1011_nl = nl_MultLoop_acc_1011_nl[24:0];
  assign nl_MultLoop_acc_1733_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_16_18({MultLoop_acc_3974_cse_1
      , (data_rsci_idat[223:219])});
  assign MultLoop_acc_1733_nl = nl_MultLoop_acc_1733_nl[17:0];
  assign nl_MultLoop_acc_1734_nl = ({(data_rsci_idat[233:216]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_1733_nl);
  assign MultLoop_acc_1734_nl = nl_MultLoop_acc_1734_nl[20:0];
  assign nl_MultLoop_acc_1008_nl = conv_s2u_21_23(MultLoop_acc_1734_nl) + ({(~ (data_rsci_idat[233:216]))
      , 5'b00000});
  assign MultLoop_acc_1008_nl = nl_MultLoop_acc_1008_nl[22:0];
  assign nl_MultLoop_acc_4600_nl = conv_s2u_19_24(MultLoop_acc_1735_cse_1[20:2])
      + ({(data_rsci_idat[251:234]) , 6'b000001});
  assign MultLoop_acc_4600_nl = nl_MultLoop_acc_4600_nl[23:0];
  assign nl_MultLoop_acc_1740_nl = ({(data_rsci_idat[107:90]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[107:90])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_1740_nl = nl_MultLoop_acc_1740_nl[21:0];
  assign nl_MultLoop_acc_1001_nl = conv_s2s_22_25(MultLoop_acc_1740_nl) + conv_s2s_24_25({(data_rsci_idat[107:90])
      , 6'b000000});
  assign MultLoop_acc_1001_nl = nl_MultLoop_acc_1001_nl[24:0];
  assign nl_MultLoop_acc_1742_nl = conv_s2s_20_21({(data_rsci_idat[35:18]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_1741_cse_1);
  assign MultLoop_acc_1742_nl = nl_MultLoop_acc_1742_nl[20:0];
  assign nl_MultLoop_acc_1417_nl = conv_s2u_21_23(MultLoop_acc_1742_nl) + conv_s2u_22_23({(data_rsci_idat[35:18])
      , 4'b0000});
  assign MultLoop_acc_1417_nl = nl_MultLoop_acc_1417_nl[22:0];
  assign nl_MultLoop_acc_1797_itm_1  = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_3975_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_1000_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_3973_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_1011_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1008_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_4600_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_1001_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1417_nl)));
  assign nl_MultLoop_acc_4500_nl =  -conv_s2s_14_15(data_rsci_idat[197:184]);
  assign MultLoop_acc_4500_nl = nl_MultLoop_acc_4500_nl[14:0];
  assign nl_MultLoop_acc_106_nl = conv_s2s_22_23({(~ (data_rsci_idat[197:180])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[197:180])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_4500_nl)
      , (~ (data_rsci_idat[183:180]))});
  assign MultLoop_acc_106_nl = nl_MultLoop_acc_106_nl[22:0];
  assign nl_MultLoop_acc_4501_nl =  -conv_s2s_11_12(data_rsci_idat[215:205]);
  assign MultLoop_acc_4501_nl = nl_MultLoop_acc_4501_nl[11:0];
  assign nl_MultLoop_acc_107_nl = conv_s2s_25_26({(~ (data_rsci_idat[215:198])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[215:198])) , 5'b00001}) +
      conv_s2s_19_26({(MultLoop_acc_4501_nl) , (~ (data_rsci_idat[204:198]))});
  assign MultLoop_acc_107_nl = nl_MultLoop_acc_107_nl[25:0];
  assign nl_MultLoop_acc_101_nl = conv_s2s_25_26({(~ (data_rsci_idat[107:90])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[107:90])) , 5'b00100}) +
      conv_s2s_21_26(MultLoop_acc_1618_cse_1);
  assign MultLoop_acc_101_nl = nl_MultLoop_acc_101_nl[25:0];
  assign nl_MultLoop_acc_3720_itm_1  = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_106_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_107_nl))) + conv_s2s_16_18(MultLoop_acc_1145_itm_22_7)
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_101_nl)));
  assign nl_MultLoop_acc_3676_nl = (~ (data_rsci_idat[827:810])) + conv_s2s_16_18({Result_acc_178_cse_1
      , (data_rsci_idat[817:813])});
  assign MultLoop_acc_3676_nl = nl_MultLoop_acc_3676_nl[17:0];
  assign nl_MultLoop_acc_3677_nl = conv_s2s_20_21({(~ (data_rsci_idat[827:810]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3676_nl);
  assign MultLoop_acc_3677_nl = nl_MultLoop_acc_3677_nl[20:0];
  assign nl_MultLoop_acc_1120_nl = conv_s2u_21_24(MultLoop_acc_3677_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[827:810])) , 5'b00100});
  assign MultLoop_acc_1120_nl = nl_MultLoop_acc_1120_nl[23:0];
  assign nl_MultLoop_acc_3679_nl = (~ (data_rsci_idat[773:756])) + conv_s2s_17_18({MultLoop_acc_4233_cse_1
      , (data_rsci_idat[762:758])});
  assign MultLoop_acc_3679_nl = nl_MultLoop_acc_3679_nl[17:0];
  assign nl_MultLoop_acc_3680_nl = conv_s2s_20_21({(~ (data_rsci_idat[773:756]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3679_nl);
  assign MultLoop_acc_3680_nl = nl_MultLoop_acc_3680_nl[20:0];
  assign nl_MultLoop_acc_1117_nl = conv_s2u_21_24(MultLoop_acc_3680_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[773:756])) , 5'b00100});
  assign MultLoop_acc_1117_nl = nl_MultLoop_acc_1117_nl[23:0];
  assign nl_MultLoop_acc_3719_itm_1  = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1120_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1117_nl)));
  assign nl_MultLoop_acc_4505_nl = conv_s2s_13_14(data_rsci_idat[125:113]) + 14'b00000000000001;
  assign MultLoop_acc_4505_nl = nl_MultLoop_acc_4505_nl[13:0];
  assign nl_MultLoop_acc_3682_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_17_18({(MultLoop_acc_4505_nl)
      , (data_rsci_idat[112:110])});
  assign MultLoop_acc_3682_nl = nl_MultLoop_acc_3682_nl[17:0];
  assign nl_MultLoop_acc_1104_nl = conv_s2u_18_22(MultLoop_acc_3682_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[125:108])) , 3'b001});
  assign MultLoop_acc_1104_nl = nl_MultLoop_acc_1104_nl[21:0];
  assign nl_MultLoop_acc_4506_nl = conv_s2s_11_12(data_rsci_idat[53:43]) + 12'b000000000001;
  assign MultLoop_acc_4506_nl = nl_MultLoop_acc_4506_nl[11:0];
  assign nl_MultLoop_acc_3687_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_14_18({(MultLoop_acc_4506_nl)
      , (data_rsci_idat[42:41])});
  assign MultLoop_acc_3687_nl = nl_MultLoop_acc_3687_nl[17:0];
  assign nl_MultLoop_acc_1102_nl = conv_s2u_18_21(MultLoop_acc_3687_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[53:36])) , 2'b01});
  assign MultLoop_acc_1102_nl = nl_MultLoop_acc_1102_nl[20:0];
  assign nl_MultLoop_acc_3688_nl = conv_s2s_18_19(data_rsci_idat[71:54]) + conv_s2s_16_19(data_rsci_idat[71:56]);
  assign MultLoop_acc_3688_nl = nl_MultLoop_acc_3688_nl[18:0];
  assign nl_MultLoop_acc_1103_nl = conv_s2u_19_21(MultLoop_acc_3688_nl) + conv_s2u_20_21({(data_rsci_idat[71:54])
      , 2'b00});
  assign MultLoop_acc_1103_nl = nl_MultLoop_acc_1103_nl[20:0];
  assign nl_MultLoop_acc_4653_nl = conv_s2u_18_20(MultLoop_acc_3556_itm_19_2_1) +
      ({(data_rsci_idat[35:18]) , 2'b01});
  assign MultLoop_acc_4653_nl = nl_MultLoop_acc_4653_nl[19:0];
  assign nl_MultLoop_acc_4696_nl = conv_s2u_16_19(MultLoop_acc_3683_itm_18_3_1) +
      conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_4696_nl = nl_MultLoop_acc_4696_nl[18:0];
  assign nl_MultLoop_97_MultLoop_acc_3_nl = (readslicef_19_14_5((MultLoop_acc_4696_nl)))
      + 14'b11111100011101;
  assign MultLoop_97_MultLoop_acc_3_nl = nl_MultLoop_97_MultLoop_acc_3_nl[13:0];
  assign nl_MultLoop_100_MultLoop_acc_3_nl = conv_s2s_16_17(readslicef_21_16_5((MultLoop_acc_1102_nl)))
      + conv_s2s_16_17(readslicef_21_16_5((MultLoop_acc_1103_nl))) + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_4653_nl)))
      + conv_s2s_14_17(MultLoop_97_MultLoop_acc_3_nl);
  assign MultLoop_100_MultLoop_acc_3_nl = nl_MultLoop_100_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_3718_itm_1  = conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1104_nl)))
      + conv_s2s_17_18(MultLoop_100_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_4507_nl =  -conv_s2s_15_16(data_rsci_idat[89:75]);
  assign MultLoop_acc_4507_nl = nl_MultLoop_acc_4507_nl[15:0];
  assign nl_MultLoop_acc_100_nl = conv_s2s_19_22({(MultLoop_acc_4507_nl) , (~ (data_rsci_idat[74:72]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[89:72])) , 3'b001});
  assign MultLoop_acc_100_nl = nl_MultLoop_acc_100_nl[21:0];
  assign nl_MultLoop_acc_4508_nl =  -conv_s2s_16_17(data_rsci_idat[143:128]);
  assign MultLoop_acc_4508_nl = nl_MultLoop_acc_4508_nl[16:0];
  assign nl_MultLoop_acc_103_nl = conv_s2s_19_21({(MultLoop_acc_4508_nl) , (~ (data_rsci_idat[127:126]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[143:126])) , 2'b01});
  assign MultLoop_acc_103_nl = nl_MultLoop_acc_103_nl[20:0];
  assign nl_MultLoop_acc_4509_nl =  -conv_s2s_14_15(data_rsci_idat[701:688]);
  assign MultLoop_acc_4509_nl = nl_MultLoop_acc_4509_nl[14:0];
  assign nl_MultLoop_acc_3618_nl = ({(data_rsci_idat[701:684]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4509_nl)
      , (~ (data_rsci_idat[687:684]))});
  assign MultLoop_acc_3618_nl = nl_MultLoop_acc_3618_nl[19:0];
  assign nl_MultLoop_acc_134_nl = conv_s2s_20_22(MultLoop_acc_3618_nl) + ({(~ (data_rsci_idat[701:684]))
      , 4'b0000});
  assign MultLoop_acc_134_nl = nl_MultLoop_acc_134_nl[21:0];
  assign nl_MultLoop_acc_3696_nl = (readslicef_21_15_6((MultLoop_acc_103_nl))) +
      conv_s2s_13_15(MultLoop_acc_2057_cse_1[18:6]) + conv_s2s_12_15(readslicef_22_12_10((MultLoop_acc_134_nl)));
  assign MultLoop_acc_3696_nl = nl_MultLoop_acc_3696_nl[14:0];
  assign nl_MultLoop_acc_3621_nl = conv_s2s_22_23({(~ (data_rsci_idat[629:612]))
      , 4'b0100}) + conv_s2s_21_23(MultLoop_acc_4688);
  assign MultLoop_acc_3621_nl = nl_MultLoop_acc_3621_nl[22:0];
  assign nl_MultLoop_acc_130_nl = conv_s2s_23_24(MultLoop_acc_3621_nl) + ({(data_rsci_idat[629:612])
      , 6'b010000});
  assign MultLoop_acc_130_nl = nl_MultLoop_acc_130_nl[23:0];
  assign nl_MultLoop_acc_3622_nl = conv_s2s_18_19(data_rsci_idat[593:576]) + conv_s2s_16_19(data_rsci_idat[593:578]);
  assign MultLoop_acc_3622_nl = nl_MultLoop_acc_3622_nl[18:0];
  assign nl_MultLoop_acc_1115_nl = conv_s2u_19_22(MultLoop_acc_3622_nl) + conv_s2u_21_22({(data_rsci_idat[593:576])
      , 3'b000});
  assign MultLoop_acc_1115_nl = nl_MultLoop_acc_1115_nl[21:0];
  assign nl_MultLoop_acc_3717_itm_1_16_0  = (readslicef_22_17_5((MultLoop_acc_100_nl)))
      + conv_s2s_15_17(MultLoop_acc_3696_nl) + conv_s2s_14_17(readslicef_24_14_10((MultLoop_acc_130_nl)))
      + conv_s2s_14_17(readslicef_22_14_8((MultLoop_acc_1115_nl)));
  assign nl_MultLoop_acc_3624_nl = (~ (data_rsci_idat[809:792])) + conv_s2s_15_18(data_rsci_idat[809:795]);
  assign MultLoop_acc_3624_nl = nl_MultLoop_acc_3624_nl[17:0];
  assign nl_MultLoop_acc_3625_nl = conv_s2s_20_21({(~ (data_rsci_idat[809:792]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3624_nl);
  assign MultLoop_acc_3625_nl = nl_MultLoop_acc_3625_nl[20:0];
  assign nl_MultLoop_acc_1119_nl = conv_s2u_21_22(MultLoop_acc_3625_nl) + ({(data_rsci_idat[809:792])
      , 4'b0100});
  assign MultLoop_acc_1119_nl = nl_MultLoop_acc_1119_nl[21:0];
  assign nl_MultLoop_acc_4510_nl =  -conv_s2s_11_12(data_rsci_idat[647:637]);
  assign MultLoop_acc_4510_nl = nl_MultLoop_acc_4510_nl[11:0];
  assign nl_MultLoop_acc_3628_nl = ({(data_rsci_idat[647:630]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[647:630])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_4510_nl)
      , (~ (data_rsci_idat[636:630]))});
  assign MultLoop_acc_3628_nl = nl_MultLoop_acc_3628_nl[22:0];
  assign nl_MultLoop_acc_4511_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3628_nl)))
      + (~ (data_rsci_idat[647:630]));
  assign MultLoop_acc_4511_nl = nl_MultLoop_acc_4511_nl[17:0];
  assign nl_MultLoop_acc_3623_nl = conv_s2s_22_23({(~ (data_rsci_idat[449:432]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[449:432]));
  assign MultLoop_acc_3623_nl = nl_MultLoop_acc_3623_nl[22:0];
  assign nl_MultLoop_acc_120_nl = conv_s2s_23_24(MultLoop_acc_3623_nl) + ({(data_rsci_idat[449:432])
      , 6'b010000});
  assign MultLoop_acc_120_nl = nl_MultLoop_acc_120_nl[23:0];
  assign nl_MultLoop_acc_1105_nl = conv_s2u_14_19(data_rsci_idat[161:148]) + conv_s2u_18_19(data_rsci_idat[161:144]);
  assign MultLoop_acc_1105_nl = nl_MultLoop_acc_1105_nl[18:0];
  assign nl_MultLoop_acc_1112_nl = conv_s2u_18_21(MultLoop_acc_2535_cse_1) + ({(data_rsci_idat[485:468])
      , 3'b001});
  assign MultLoop_acc_1112_nl = nl_MultLoop_acc_1112_nl[20:0];
  assign nl_MultLoop_acc_3716_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1119_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4511_nl))) + conv_s2s_14_17(readslicef_24_14_10((MultLoop_acc_120_nl)))
      + conv_s2s_14_17(MultLoop_acc_4589_itm_19_4[15:2]) + conv_s2s_14_17(readslicef_19_14_5((MultLoop_acc_1105_nl)))
      + conv_s2s_13_17(readslicef_21_13_8((MultLoop_acc_1112_nl)));
  assign nl_MultLoop_acc_4512_nl = conv_s2s_14_15(data_rsci_idat[611:598]) + 15'b000000000000001;
  assign MultLoop_acc_4512_nl = nl_MultLoop_acc_4512_nl[14:0];
  assign nl_MultLoop_acc_3630_nl = conv_s2s_18_19(data_rsci_idat[611:594]) + conv_s2s_17_19({(MultLoop_acc_4512_nl)
      , (data_rsci_idat[597:596])});
  assign MultLoop_acc_3630_nl = nl_MultLoop_acc_3630_nl[18:0];
  assign nl_MultLoop_acc_129_nl = conv_s2u_19_20(MultLoop_acc_3630_nl) + ({(~ (data_rsci_idat[611:594]))
      , 2'b00});
  assign MultLoop_acc_129_nl = nl_MultLoop_acc_129_nl[19:0];
  assign nl_MultLoop_acc_3631_nl = (~ (data_rsci_idat[539:522])) + conv_s2s_14_18(data_rsci_idat[539:526]);
  assign MultLoop_acc_3631_nl = nl_MultLoop_acc_3631_nl[17:0];
  assign nl_MultLoop_acc_1114_nl = conv_s2u_18_20(MultLoop_acc_3631_nl) + ({(data_rsci_idat[539:522])
      , 2'b01});
  assign MultLoop_acc_1114_nl = nl_MultLoop_acc_1114_nl[19:0];
  assign nl_MultLoop_acc_3633_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_16_19({MultLoop_acc_3946_cse_1
      , (data_rsci_idat[401:399])});
  assign MultLoop_acc_3633_nl = nl_MultLoop_acc_3633_nl[18:0];
  assign nl_MultLoop_acc_118_nl = conv_s2u_19_21(MultLoop_acc_3633_nl) + ({(~ (data_rsci_idat[413:396]))
      , 3'b000});
  assign MultLoop_acc_118_nl = nl_MultLoop_acc_118_nl[20:0];
  assign nl_MultLoop_acc_3715_itm_1  = conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_129_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1114_nl))) + conv_s2s_15_17(MultLoop_acc_123_itm_17_3)
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_118_nl)));
  assign nl_MultLoop_acc_3635_nl = ({(data_rsci_idat[845:828]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[845:828]));
  assign MultLoop_acc_3635_nl = nl_MultLoop_acc_3635_nl[21:0];
  assign nl_MultLoop_acc_4514_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_3635_nl)))
      + conv_s2u_18_19(data_rsci_idat[845:828]);
  assign MultLoop_acc_4514_nl = nl_MultLoop_acc_4514_nl[18:0];
  assign nl_MultLoop_acc_3637_nl = ({(~ (data_rsci_idat[863:846])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_3636_cse_1);
  assign MultLoop_acc_3637_nl = nl_MultLoop_acc_3637_nl[22:0];
  assign nl_MultLoop_acc_143_nl = conv_s2s_23_25(MultLoop_acc_3637_nl) + ({(data_rsci_idat[863:846])
      , 7'b0100000});
  assign MultLoop_acc_143_nl = nl_MultLoop_acc_143_nl[24:0];
  assign nl_MultLoop_acc_3639_nl = (~ (data_rsci_idat[791:774])) + conv_s2s_17_18({MultLoop_acc_4083_cse_1
      , (data_rsci_idat[780:776])});
  assign MultLoop_acc_3639_nl = nl_MultLoop_acc_3639_nl[17:0];
  assign nl_MultLoop_acc_3640_nl = conv_s2s_20_21({(~ (data_rsci_idat[791:774]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3639_nl);
  assign MultLoop_acc_3640_nl = nl_MultLoop_acc_3640_nl[20:0];
  assign nl_MultLoop_acc_1118_nl = conv_s2u_21_24(MultLoop_acc_3640_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[791:774])) , 5'b00100});
  assign MultLoop_acc_1118_nl = nl_MultLoop_acc_1118_nl[23:0];
  assign nl_MultLoop_acc_110_nl = conv_s2u_13_18(data_rsci_idat[269:257]) - (data_rsci_idat[269:252]);
  assign MultLoop_acc_110_nl = nl_MultLoop_acc_110_nl[17:0];
  assign nl_MultLoop_acc_3725_itm_1  = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4514_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_143_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1118_nl)))
      + conv_s2s_15_18(MultLoop_acc_119_itm_23_9) + conv_s2s_15_18(readslicef_18_15_3((MultLoop_acc_110_nl)));
  assign nl_MultLoop_acc_4686_nl = ({(data_rsci_idat[737:720]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_1949_cse_1[20:2]);
  assign MultLoop_acc_4686_nl = nl_MultLoop_acc_4686_nl[19:0];
  assign nl_MultLoop_acc_4517_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_4686_nl)))
      + (~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_4517_nl = nl_MultLoop_acc_4517_nl[17:0];
  assign nl_MultLoop_acc_3646_nl = conv_s2s_22_23({(data_rsci_idat[755:738]) , 4'b0000})
      + conv_s2s_18_23(data_rsci_idat[755:738]) + conv_s2s_17_23({Result_acc_214_cse_1
      , (data_rsci_idat[745:740])});
  assign MultLoop_acc_3646_nl = nl_MultLoop_acc_3646_nl[22:0];
  assign nl_MultLoop_acc_4519_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3646_nl)))
      + (~ (data_rsci_idat[755:738]));
  assign MultLoop_acc_4519_nl = nl_MultLoop_acc_4519_nl[17:0];
  assign nl_MultLoop_acc_4520_nl = conv_s2s_12_13(data_rsci_idat[665:654]) + 13'b0000000000001;
  assign MultLoop_acc_4520_nl = nl_MultLoop_acc_4520_nl[12:0];
  assign nl_MultLoop_acc_3648_nl = conv_s2s_18_19(data_rsci_idat[665:648]) + conv_s2s_17_19({(MultLoop_acc_4520_nl)
      , (data_rsci_idat[653:650])});
  assign MultLoop_acc_3648_nl = nl_MultLoop_acc_3648_nl[18:0];
  assign nl_MultLoop_acc_132_nl = conv_s2u_19_22(MultLoop_acc_3648_nl) + ({(~ (data_rsci_idat[665:648]))
      , 4'b0000});
  assign MultLoop_acc_132_nl = nl_MultLoop_acc_132_nl[21:0];
  assign nl_MultLoop_acc_3724_itm_1  = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4517_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4519_nl))) + conv_s2s_16_18(MultLoop_acc_87_itm_19_4)
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_132_nl)));
  assign nl_MultLoop_acc_3649_nl = (~ (data_rsci_idat[683:666])) + conv_s2s_15_18(data_rsci_idat[683:669]);
  assign MultLoop_acc_3649_nl = nl_MultLoop_acc_3649_nl[17:0];
  assign nl_MultLoop_acc_1116_nl = conv_s2u_18_20(MultLoop_acc_3649_nl) + ({(data_rsci_idat[683:666])
      , 2'b01});
  assign MultLoop_acc_1116_nl = nl_MultLoop_acc_1116_nl[19:0];
  assign nl_MultLoop_acc_126_nl = conv_s2s_25_26({(~ (data_rsci_idat[557:540])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[557:540])) , 5'b01000}) +
      conv_s2s_21_26({(~ (data_rsci_idat[557:540])) , 3'b001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_700_18_7
      , (~ (data_rsci_idat[546:540]))});
  assign MultLoop_acc_126_nl = nl_MultLoop_acc_126_nl[25:0];
  assign nl_MultLoop_acc_3710_itm_1  = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_1116_nl)))
      + conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_126_nl)));
  assign nl_MultLoop_acc_3654_nl = ({(data_rsci_idat[575:558]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_686_18_6
      , (~ (data_rsci_idat[563:558]))});
  assign MultLoop_acc_3654_nl = nl_MultLoop_acc_3654_nl[19:0];
  assign nl_MultLoop_acc_4523_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_3654_nl)))
      + (~ (data_rsci_idat[575:558]));
  assign MultLoop_acc_4523_nl = nl_MultLoop_acc_4523_nl[17:0];
  assign nl_MultLoop_acc_3709_itm_1  = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4523_nl)))
      + conv_s2s_16_17(MultLoop_acc_1095_itm_18_2[16:1]);
  assign nl_MultLoop_acc_3657_nl = ({(~ (data_rsci_idat[377:360])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[377:360])
      + conv_s2s_17_20({MultLoop_MultLoop_conc_736_16_5 , (data_rsci_idat[366:362])});
  assign MultLoop_acc_3657_nl = nl_MultLoop_acc_3657_nl[19:0];
  assign nl_MultLoop_acc_1110_nl = conv_s2u_20_24(MultLoop_acc_3657_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[377:360])) , 5'b00100});
  assign MultLoop_acc_1110_nl = nl_MultLoop_acc_1110_nl[23:0];
  assign nl_MultLoop_acc_1111_nl = conv_s2u_16_19(data_rsci_idat[395:380]) + conv_s2u_18_19(data_rsci_idat[395:378]);
  assign MultLoop_acc_1111_nl = nl_MultLoop_acc_1111_nl[18:0];
  assign nl_MultLoop_acc_4525_nl = conv_s2u_14_19(MultLoop_acc_447_itm_20_7) + conv_s2u_18_19(data_rsci_idat[341:324]);
  assign MultLoop_acc_4525_nl = nl_MultLoop_acc_4525_nl[18:0];
  assign nl_MultLoop_acc_3722_itm_1  = conv_s2s_16_18(MultLoop_acc_3918_itm_17_2)
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1110_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1111_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4525_nl)));
  assign nl_MultLoop_acc_3659_nl = ({(data_rsci_idat[359:342]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[359:342]));
  assign MultLoop_acc_3659_nl = nl_MultLoop_acc_3659_nl[19:0];
  assign nl_MultLoop_acc_3660_nl = ({(~ (data_rsci_idat[359:342])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3659_nl);
  assign MultLoop_acc_3660_nl = nl_MultLoop_acc_3660_nl[21:0];
  assign nl_MultLoop_acc_115_nl = conv_s2s_22_24(MultLoop_acc_3660_nl) + ({(data_rsci_idat[359:342])
      , 6'b010000});
  assign MultLoop_acc_115_nl = nl_MultLoop_acc_115_nl[23:0];
  assign nl_MultLoop_acc_4654_nl = conv_s2u_17_19(MultLoop_acc_3661_cse_1[18:2])
      + conv_s2u_18_19(data_rsci_idat[323:306]);
  assign MultLoop_acc_4654_nl = nl_MultLoop_acc_4654_nl[18:0];
  assign nl_MultLoop_acc_3706_itm_1  = conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_115_nl)))
      + conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4654_nl)));
  assign nl_MultLoop_acc_4526_nl =  -conv_s2s_10_11(data_rsci_idat[233:224]);
  assign MultLoop_acc_4526_nl = nl_MultLoop_acc_4526_nl[10:0];
  assign nl_MultLoop_acc_3665_nl = ({(data_rsci_idat[233:216]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[233:216])) , 4'b0100}) + conv_s2s_20_24({(~ (data_rsci_idat[233:216]))
      , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4526_nl) , (~ (data_rsci_idat[223:216]))});
  assign MultLoop_acc_3665_nl = nl_MultLoop_acc_3665_nl[23:0];
  assign nl_MultLoop_acc_4527_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3665_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_4527_nl = nl_MultLoop_acc_4527_nl[17:0];
  assign nl_MultLoop_acc_3667_nl = ({(~ (data_rsci_idat[251:234])) , 4'b0000}) +
      conv_s2s_19_22(MultLoop_acc_2591_cse_1);
  assign MultLoop_acc_3667_nl = nl_MultLoop_acc_3667_nl[21:0];
  assign nl_MultLoop_acc_1107_nl = conv_s2u_22_24(MultLoop_acc_3667_nl) + ({(data_rsci_idat[251:234])
      , 6'b010000});
  assign MultLoop_acc_1107_nl = nl_MultLoop_acc_1107_nl[23:0];
  assign nl_MultLoop_acc_3705_itm_1  = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4527_nl)))
      + conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_1107_nl)));
  assign nl_MultLoop_acc_1838_nl = (~ (data_rsci_idat[287:270])) + conv_s2s_16_18({MultLoop_acc_3976_cse_1
      , (data_rsci_idat[277:273])});
  assign MultLoop_acc_1838_nl = nl_MultLoop_acc_1838_nl[17:0];
  assign nl_MultLoop_acc_1839_nl = ({(data_rsci_idat[287:270]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1838_nl);
  assign MultLoop_acc_1839_nl = nl_MultLoop_acc_1839_nl[19:0];
  assign nl_MultLoop_acc_965_nl = conv_s2u_20_23(MultLoop_acc_1839_nl) + ({(~ (data_rsci_idat[287:270]))
      , 5'b00000});
  assign MultLoop_acc_965_nl = nl_MultLoop_acc_965_nl[22:0];
  assign nl_MultLoop_acc_3977_nl = conv_s2s_11_12(data_rsci_idat[233:223]) + 12'b000000000001;
  assign MultLoop_acc_3977_nl = nl_MultLoop_acc_3977_nl[11:0];
  assign nl_MultLoop_acc_1841_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_16_18({(MultLoop_acc_3977_nl)
      , (data_rsci_idat[222:219])});
  assign MultLoop_acc_1841_nl = nl_MultLoop_acc_1841_nl[17:0];
  assign nl_MultLoop_acc_1405_nl = conv_s2u_18_23(MultLoop_acc_1841_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[233:216])) , 4'b0001});
  assign MultLoop_acc_1405_nl = nl_MultLoop_acc_1405_nl[22:0];
  assign nl_MultLoop_acc_1843_nl = conv_s2s_24_25({(~ (data_rsci_idat[251:234]))
      , 6'b000100}) + conv_s2s_21_25(MultLoop_acc_1735_cse_1);
  assign MultLoop_acc_1843_nl = nl_MultLoop_acc_1843_nl[24:0];
  assign nl_MultLoop_acc_963_nl = conv_s2s_25_26(MultLoop_acc_1843_nl) + ({(data_rsci_idat[251:234])
      , 8'b01000000});
  assign MultLoop_acc_963_nl = nl_MultLoop_acc_963_nl[25:0];
  assign nl_MultLoop_acc_1911_itm_1  = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_965_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1405_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_963_nl)))
      + conv_s2s_16_18(MultLoop_acc_3920_itm_17_2);
  assign nl_MultLoop_acc_1403_nl = conv_s2u_18_22(MultLoop_acc_1844_cse_1) + ({(data_rsci_idat[161:144])
      , 4'b0001});
  assign MultLoop_acc_1403_nl = nl_MultLoop_acc_1403_nl[21:0];
  assign nl_MultLoop_acc_1846_nl = ({(~ (data_rsci_idat[179:162])) , 4'b0000}) +
      conv_s2s_18_22(data_rsci_idat[179:162]) + conv_s2s_16_22(data_rsci_idat[179:164]);
  assign MultLoop_acc_1846_nl = nl_MultLoop_acc_1846_nl[21:0];
  assign nl_MultLoop_acc_1404_nl = conv_s2u_22_24(MultLoop_acc_1846_nl) + ({(data_rsci_idat[179:162])
      , 6'b010000});
  assign MultLoop_acc_1404_nl = nl_MultLoop_acc_1404_nl[23:0];
  assign nl_MultLoop_acc_4664_nl = conv_s2u_16_19(MultLoop_acc_1848_itm_21_6) + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_4664_nl = nl_MultLoop_acc_4664_nl[18:0];
  assign nl_MultLoop_acc_954_nl = conv_s2s_25_26({(~ (data_rsci_idat[89:72])) , 7'b0100000})
      + conv_s2s_23_26({(~ (data_rsci_idat[89:72])) , 5'b00100}) + conv_s2s_20_26({(~
      (data_rsci_idat[89:72])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_804_18_7
      , (~ (data_rsci_idat[78:72]))});
  assign MultLoop_acc_954_nl = nl_MultLoop_acc_954_nl[25:0];
  assign nl_MultLoop_acc_1910_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1403_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1404_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4664_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_954_nl)));
  assign nl_MultLoop_acc_3981_nl =  -conv_s2s_10_11(data_rsci_idat[755:746]);
  assign MultLoop_acc_3981_nl = nl_MultLoop_acc_3981_nl[10:0];
  assign nl_MultLoop_acc_1856_nl = ({(data_rsci_idat[755:738]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_3981_nl)
      , (~ (data_rsci_idat[745:738]))});
  assign MultLoop_acc_1856_nl = nl_MultLoop_acc_1856_nl[19:0];
  assign nl_MultLoop_acc_3982_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_14_18(readslicef_20_14_6((MultLoop_acc_1856_nl)));
  assign MultLoop_acc_3982_nl = nl_MultLoop_acc_3982_nl[17:0];
  assign nl_MultLoop_acc_3983_nl = conv_s2u_18_21(MultLoop_acc_3982_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[755:738])) , 2'b01});
  assign MultLoop_acc_3983_nl = nl_MultLoop_acc_3983_nl[20:0];
  assign nl_MultLoop_acc_4601_nl = conv_s2u_15_19(MultLoop_acc_1541_itm_18_2[16:2])
      + conv_s2u_18_19(data_rsci_idat[701:684]);
  assign MultLoop_acc_4601_nl = nl_MultLoop_acc_4601_nl[18:0];
  assign nl_MultLoop_acc_3984_nl =  -conv_s2s_11_12(data_rsci_idat[665:655]);
  assign MultLoop_acc_3984_nl = nl_MultLoop_acc_3984_nl[11:0];
  assign nl_MultLoop_acc_1860_nl = ({(data_rsci_idat[665:648]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_3984_nl)
      , (~ (data_rsci_idat[654:648]))});
  assign MultLoop_acc_1860_nl = nl_MultLoop_acc_1860_nl[19:0];
  assign nl_MultLoop_acc_1861_nl = ({(~ (data_rsci_idat[665:648])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_1860_nl);
  assign MultLoop_acc_1861_nl = nl_MultLoop_acc_1861_nl[21:0];
  assign nl_MultLoop_acc_984_nl = conv_s2s_22_26(MultLoop_acc_1861_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[665:648])) , 7'b0010000});
  assign MultLoop_acc_984_nl = nl_MultLoop_acc_984_nl[25:0];
  assign nl_MultLoop_acc_1853_nl = ({(data_rsci_idat[53:36]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_802_18_8
      , (~ (data_rsci_idat[43:36]))});
  assign MultLoop_acc_1853_nl = nl_MultLoop_acc_1853_nl[19:0];
  assign nl_MultLoop_acc_1854_nl = conv_s2s_22_23({(data_rsci_idat[53:36]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_1853_nl);
  assign MultLoop_acc_1854_nl = nl_MultLoop_acc_1854_nl[22:0];
  assign nl_MultLoop_acc_3980_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_1854_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_3980_nl = nl_MultLoop_acc_3980_nl[17:0];
  assign nl_MultLoop_acc_953_nl = conv_s2s_18_20(~ (data_rsci_idat[71:54])) + ({(data_rsci_idat[71:54])
      , 2'b01});
  assign MultLoop_acc_953_nl = nl_MultLoop_acc_953_nl[19:0];
  assign nl_MultLoop_acc_1918_itm_1  = conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_3983_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4601_nl))) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_984_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_3980_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_953_nl)));
  assign nl_MultLoop_acc_1863_nl = ({(data_rsci_idat[629:612]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_766_18_7
      , (~ (data_rsci_idat[618:612]))});
  assign MultLoop_acc_1863_nl = nl_MultLoop_acc_1863_nl[19:0];
  assign nl_MultLoop_acc_1864_nl = ({(~ (data_rsci_idat[629:612])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_1863_nl);
  assign MultLoop_acc_1864_nl = nl_MultLoop_acc_1864_nl[22:0];
  assign nl_MultLoop_acc_982_nl = conv_s2s_23_26(MultLoop_acc_1864_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[629:612])) , 7'b0100000});
  assign MultLoop_acc_982_nl = nl_MultLoop_acc_982_nl[25:0];
  assign nl_MultLoop_acc_4665_nl = conv_s2u_19_24(MultLoop_acc_1866_itm_20_2_1) +
      conv_s2u_23_24({(~ (data_rsci_idat[593:576])) , 5'b00001});
  assign MultLoop_acc_4665_nl = nl_MultLoop_acc_4665_nl[23:0];
  assign nl_MultLoop_acc_1869_nl = ({(~ (data_rsci_idat[521:504])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[521:504])
      + conv_s2s_15_20({MultLoop_acc_3987_cse_1 , (data_rsci_idat[511:508])});
  assign MultLoop_acc_1869_nl = nl_MultLoop_acc_1869_nl[19:0];
  assign nl_MultLoop_acc_1410_nl = conv_s2u_20_23(MultLoop_acc_1869_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[521:504])) , 4'b0100});
  assign MultLoop_acc_1410_nl = nl_MultLoop_acc_1410_nl[22:0];
  assign nl_MultLoop_acc_974_nl = conv_s2s_25_26({(~ (data_rsci_idat[467:450])) ,
      7'b0000100}) + conv_s2s_20_26({(~ (data_rsci_idat[467:450])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_678_18_7
      , (~ (data_rsci_idat[456:450]))});
  assign MultLoop_acc_974_nl = nl_MultLoop_acc_974_nl[25:0];
  assign nl_MultLoop_acc_1917_itm_1  = conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_982_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_4665_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1410_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_974_nl)));
  assign nl_MultLoop_acc_3991_nl =  -conv_s2s_12_13(data_rsci_idat[35:24]);
  assign MultLoop_acc_3991_nl = nl_MultLoop_acc_3991_nl[12:0];
  assign nl_MultLoop_acc_951_nl = conv_s2s_19_25({(MultLoop_acc_3991_nl) , (~ (data_rsci_idat[23:18]))})
      + conv_s2s_24_25({(~ (data_rsci_idat[35:18])) , 6'b000001});
  assign MultLoop_acc_951_nl = nl_MultLoop_acc_951_nl[24:0];
  assign nl_MultLoop_acc_991_nl = conv_s2s_19_23({MultLoop_MultLoop_conc_738_18_4
      , (~ (data_rsci_idat[777:774]))}) + conv_s2s_22_23({(~ (data_rsci_idat[791:774]))
      , 4'b0001});
  assign MultLoop_acc_991_nl = nl_MultLoop_acc_991_nl[22:0];
  assign nl_MultLoop_acc_970_nl = conv_s2u_16_18(data_rsci_idat[377:362]) - (data_rsci_idat[377:360]);
  assign MultLoop_acc_970_nl = nl_MultLoop_acc_970_nl[17:0];
  assign nl_MultLoop_acc_1807_nl = (~ (data_rsci_idat[485:468])) + conv_s2s_16_18({MultLoop_MultLoop_conc_810_15_2
      , (data_rsci_idat[472:471])});
  assign MultLoop_acc_1807_nl = nl_MultLoop_acc_1807_nl[17:0];
  assign nl_MultLoop_acc_1409_nl = conv_s2u_18_21(MultLoop_acc_1807_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[485:468])) , 2'b01});
  assign MultLoop_acc_1409_nl = nl_MultLoop_acc_1409_nl[20:0];
  assign nl_MultLoop_acc_1808_nl = ({(data_rsci_idat[341:324]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[341:324]));
  assign MultLoop_acc_1808_nl = nl_MultLoop_acc_1808_nl[19:0];
  assign nl_MultLoop_acc_968_nl = conv_s2s_20_23(MultLoop_acc_1808_nl) + conv_s2s_22_23({(data_rsci_idat[341:324])
      , 4'b0000});
  assign MultLoop_acc_968_nl = nl_MultLoop_acc_968_nl[22:0];
  assign nl_MultLoop_acc_1904_nl = (readslicef_25_17_8((MultLoop_acc_951_nl))) +
      conv_s2s_14_17(readslicef_23_14_9((MultLoop_acc_991_nl))) + conv_s2s_13_17(readslicef_18_13_5((MultLoop_acc_970_nl)))
      + conv_s2s_8_17(data_rsci_idat[575:568]) + conv_s2s_14_17(readslicef_21_14_7((MultLoop_acc_1409_nl)))
      + conv_s2s_14_17(readslicef_23_14_9((MultLoop_acc_968_nl)));
  assign MultLoop_acc_1904_nl = nl_MultLoop_acc_1904_nl[16:0];
  assign nl_MultLoop_acc_1875_nl = ({(~ (data_rsci_idat[305:288])) , 4'b0000}) +
      conv_s2s_20_22({(data_rsci_idat[305:288]) , 2'b00}) + conv_s2s_18_22(data_rsci_idat[305:288])
      + conv_s2s_17_22({MultLoop_acc_3989_cse_1 , (data_rsci_idat[295:290])});
  assign MultLoop_acc_1875_nl = nl_MultLoop_acc_1875_nl[21:0];
  assign nl_MultLoop_acc_1406_nl = conv_s2u_22_25(MultLoop_acc_1875_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[305:288])) , 6'b010000});
  assign MultLoop_acc_1406_nl = nl_MultLoop_acc_1406_nl[24:0];
  assign nl_MultLoop_acc_3990_nl = conv_s2s_10_11(data_rsci_idat[107:98]) + 11'b00000000001;
  assign MultLoop_acc_3990_nl = nl_MultLoop_acc_3990_nl[10:0];
  assign nl_MultLoop_acc_1878_nl = ({(~ (data_rsci_idat[107:90])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[107:90])
      + conv_s2s_17_20({(MultLoop_acc_3990_nl) , (data_rsci_idat[97:92])});
  assign MultLoop_acc_1878_nl = nl_MultLoop_acc_1878_nl[19:0];
  assign nl_MultLoop_acc_1402_nl = conv_s2u_20_25(MultLoop_acc_1878_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[107:90])) , 6'b000100});
  assign MultLoop_acc_1402_nl = nl_MultLoop_acc_1402_nl[24:0];
  assign nl_MultLoop_acc_1916_itm_1  = conv_s2s_17_18(MultLoop_acc_1904_nl) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1406_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1402_nl)));
  assign nl_MultLoop_acc_1809_nl = conv_s2s_22_23({(~ (data_rsci_idat[737:720]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_1809_nl = nl_MultLoop_acc_1809_nl[22:0];
  assign nl_MultLoop_acc_988_nl = conv_s2s_23_25(MultLoop_acc_1809_nl) + ({(data_rsci_idat[737:720])
      , 7'b0010000});
  assign MultLoop_acc_988_nl = nl_MultLoop_acc_988_nl[24:0];
  assign nl_MultLoop_acc_3994_nl =  -conv_s2s_14_15(data_rsci_idat[773:760]);
  assign MultLoop_acc_3994_nl = nl_MultLoop_acc_3994_nl[14:0];
  assign nl_MultLoop_acc_990_nl = conv_s2s_22_23({(~ (data_rsci_idat[773:756])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[773:756])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_3994_nl)
      , (~ (data_rsci_idat[759:756]))});
  assign MultLoop_acc_990_nl = nl_MultLoop_acc_990_nl[22:0];
  assign nl_MultLoop_acc_1889_itm_1  = conv_s2s_15_16(readslicef_25_15_10((MultLoop_acc_988_nl)))
      + conv_s2s_14_16(MultLoop_acc_343_itm_19_5[14:1]) + conv_s2s_13_16(readslicef_23_13_10((MultLoop_acc_990_nl)));
  assign nl_MultLoop_acc_1888_itm_1  = conv_s2s_15_16(MultLoop_acc_4593_itm_18_3[15:1])
      + conv_s2s_15_16(data_rsci_idat[395:381]);
  assign nl_MultLoop_acc_4602_nl = conv_s2u_19_21(MultLoop_acc_1811_itm_20_2_1) +
      ({(data_rsci_idat[557:540]) , 3'b001});
  assign MultLoop_acc_4602_nl = nl_MultLoop_acc_4602_nl[20:0];
  assign nl_MultLoop_acc_3995_nl =  -conv_s2s_15_16(data_rsci_idat[503:489]);
  assign MultLoop_acc_3995_nl = nl_MultLoop_acc_3995_nl[15:0];
  assign nl_MultLoop_acc_976_nl = conv_s2s_19_22({(MultLoop_acc_3995_nl) , (~ (data_rsci_idat[488:486]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[503:486])) , 3'b001});
  assign MultLoop_acc_976_nl = nl_MultLoop_acc_976_nl[21:0];
  assign nl_MultLoop_acc_3996_nl =  -conv_s2s_11_12(data_rsci_idat[413:403]);
  assign MultLoop_acc_3996_nl = nl_MultLoop_acc_3996_nl[11:0];
  assign nl_MultLoop_acc_1814_nl = ({(data_rsci_idat[413:396]) , 5'b00001}) + conv_s2s_19_23({(MultLoop_acc_3996_nl)
      , (~ (data_rsci_idat[402:396]))});
  assign MultLoop_acc_1814_nl = nl_MultLoop_acc_1814_nl[22:0];
  assign nl_MultLoop_acc_3997_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_1814_nl)))
      + (~ (data_rsci_idat[413:396]));
  assign MultLoop_acc_3997_nl = nl_MultLoop_acc_3997_nl[17:0];
  assign nl_MultLoop_acc_4666_nl = conv_s2u_19_23(MultLoop_acc_1816_itm_20_2_1) +
      conv_s2u_22_23({(~ (data_rsci_idat[197:180])) , 4'b0001});
  assign MultLoop_acc_4666_nl = nl_MultLoop_acc_4666_nl[22:0];
  assign nl_MultLoop_acc_1902_itm_1  = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_4602_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_976_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_3997_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_4666_nl)));
  assign nl_MultLoop_acc_3999_nl = conv_s2s_10_11(data_rsci_idat[845:836]) + 11'b00000000001;
  assign MultLoop_acc_3999_nl = nl_MultLoop_acc_3999_nl[10:0];
  assign nl_MultLoop_acc_1820_nl = conv_s2s_20_21({(data_rsci_idat[845:828]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[845:828]) + conv_s2s_15_21({(MultLoop_acc_3999_nl)
      , (data_rsci_idat[835:832])});
  assign MultLoop_acc_1820_nl = nl_MultLoop_acc_1820_nl[20:0];
  assign nl_MultLoop_acc_994_nl = conv_s2u_21_22(MultLoop_acc_1820_nl) + ({(~ (data_rsci_idat[845:828]))
      , 4'b0000});
  assign MultLoop_acc_994_nl = nl_MultLoop_acc_994_nl[21:0];
  assign nl_MultLoop_acc_1823_nl = ({(~ (data_rsci_idat[863:846])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_1822_cse_1);
  assign MultLoop_acc_1823_nl = nl_MultLoop_acc_1823_nl[19:0];
  assign nl_MultLoop_acc_1416_nl = conv_s2u_20_23(MultLoop_acc_1823_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[863:846])) , 4'b0100});
  assign MultLoop_acc_1416_nl = nl_MultLoop_acc_1416_nl[22:0];
  assign nl_MultLoop_acc_1825_nl = ({(data_rsci_idat[809:792]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_682_18_8
      , (~ (data_rsci_idat[799:792]))});
  assign MultLoop_acc_1825_nl = nl_MultLoop_acc_1825_nl[22:0];
  assign nl_MultLoop_acc_4002_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_1825_nl)))
      + (~ (data_rsci_idat[809:792]));
  assign MultLoop_acc_4002_nl = nl_MultLoop_acc_4002_nl[17:0];
  assign nl_MultLoop_acc_1817_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_13_18(data_rsci_idat[17:5]);
  assign MultLoop_acc_1817_nl = nl_MultLoop_acc_1817_nl[17:0];
  assign nl_MultLoop_acc_950_nl = conv_s2u_18_20(MultLoop_acc_1817_nl) + ({(data_rsci_idat[17:0])
      , 2'b01});
  assign MultLoop_acc_950_nl = nl_MultLoop_acc_950_nl[19:0];
  assign nl_MultLoop_961_MultLoop_acc_3_nl = (readslicef_20_15_5((MultLoop_acc_950_nl)))
      + 15'b000000000010001;
  assign MultLoop_961_MultLoop_acc_3_nl = nl_MultLoop_961_MultLoop_acc_3_nl[14:0];
  assign nl_MultLoop_acc_985_nl = conv_s2s_18_23(~ (data_rsci_idat[683:666])) + ({(data_rsci_idat[683:666])
      , 5'b00001});
  assign MultLoop_acc_985_nl = nl_MultLoop_acc_985_nl[22:0];
  assign nl_MultLoop_acc_1914_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_994_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1416_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4002_nl)))
      + conv_s2s_15_18(MultLoop_961_MultLoop_acc_3_nl) + conv_s2s_13_18(readslicef_23_13_10((MultLoop_acc_985_nl)))
      + conv_s2s_13_18(MultLoop_acc_506_itm_17_5);
  assign nl_MultLoop_acc_1833_nl = conv_s2s_23_24({(~ (data_rsci_idat[431:414]))
      , 5'b00100}) + conv_s2s_21_24(MultLoop_acc_1702_cse_1);
  assign MultLoop_acc_1833_nl = nl_MultLoop_acc_1833_nl[23:0];
  assign nl_MultLoop_acc_972_nl = conv_s2s_24_26(MultLoop_acc_1833_nl) + ({(data_rsci_idat[431:414])
      , 8'b00100000});
  assign MultLoop_acc_972_nl = nl_MultLoop_acc_972_nl[25:0];
  assign nl_MultLoop_acc_1826_nl = (~ (data_rsci_idat[827:810])) + conv_s2s_16_18(data_rsci_idat[827:812]);
  assign MultLoop_acc_1826_nl = nl_MultLoop_acc_1826_nl[17:0];
  assign nl_MultLoop_acc_1828_nl = conv_s2s_22_23({(~ (data_rsci_idat[827:810]))
      , 4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[827:810])) , 2'b01}) + conv_s2s_18_23(MultLoop_acc_1826_nl);
  assign MultLoop_acc_1828_nl = nl_MultLoop_acc_1828_nl[22:0];
  assign nl_MultLoop_acc_1415_nl = conv_s2u_23_24(MultLoop_acc_1828_nl) + ({(data_rsci_idat[827:810])
      , 6'b010000});
  assign MultLoop_acc_1415_nl = nl_MultLoop_acc_1415_nl[23:0];
  assign nl_MultLoop_acc_4003_nl = conv_s2s_13_14(data_rsci_idat[611:599]) + 14'b00000000000001;
  assign MultLoop_acc_4003_nl = nl_MultLoop_acc_4003_nl[13:0];
  assign nl_MultLoop_acc_1830_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_17_18({(MultLoop_acc_4003_nl)
      , (data_rsci_idat[598:596])});
  assign MultLoop_acc_1830_nl = nl_MultLoop_acc_1830_nl[17:0];
  assign nl_MultLoop_acc_1412_nl = conv_s2u_18_22(MultLoop_acc_1830_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[611:594])) , 3'b001});
  assign MultLoop_acc_1412_nl = nl_MultLoop_acc_1412_nl[21:0];
  assign nl_MultLoop_acc_1831_nl = conv_s2s_18_19(data_rsci_idat[449:432]) + conv_s2s_14_19(data_rsci_idat[449:436]);
  assign MultLoop_acc_1831_nl = nl_MultLoop_acc_1831_nl[18:0];
  assign nl_MultLoop_acc_1408_nl = conv_s2u_19_22(MultLoop_acc_1831_nl) + conv_s2u_21_22({(data_rsci_idat[449:432])
      , 3'b000});
  assign MultLoop_acc_1408_nl = nl_MultLoop_acc_1408_nl[21:0];
  assign nl_MultLoop_acc_1834_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_15_18(data_rsci_idat[323:309]);
  assign MultLoop_acc_1834_nl = nl_MultLoop_acc_1834_nl[17:0];
  assign nl_MultLoop_acc_1407_nl = conv_s2u_18_21(MultLoop_acc_1834_nl) + ({(data_rsci_idat[323:306])
      , 3'b001});
  assign MultLoop_acc_1407_nl = nl_MultLoop_acc_1407_nl[20:0];
  assign nl_MultLoop_acc_1836_nl = conv_s2s_23_24({(~ (data_rsci_idat[269:252]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[269:252])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[269:252]));
  assign MultLoop_acc_1836_nl = nl_MultLoop_acc_1836_nl[23:0];
  assign nl_MultLoop_acc_964_nl = conv_s2s_24_26(MultLoop_acc_1836_nl) + ({(data_rsci_idat[269:252])
      , 8'b00100000});
  assign MultLoop_acc_964_nl = nl_MultLoop_acc_964_nl[25:0];
  assign nl_MultLoop_acc_1920_itm_1  = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_972_nl)))
      + conv_s2s_16_18(MultLoop_acc_826_itm_25_10) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1415_nl)))
      + conv_s2s_16_18(MultLoop_acc_1324_itm_22_7) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1412_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1408_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1407_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_964_nl)));
  assign nl_MultLoop_acc_3560_nl = conv_s2s_18_19(data_rsci_idat[719:702]) + conv_s2s_12_19(data_rsci_idat[719:708]);
  assign MultLoop_acc_3560_nl = nl_MultLoop_acc_3560_nl[18:0];
  assign nl_MultLoop_acc_1137_nl = conv_s2u_19_21(MultLoop_acc_3560_nl) + conv_s2u_20_21({(data_rsci_idat[719:702])
      , 2'b00});
  assign MultLoop_acc_1137_nl = nl_MultLoop_acc_1137_nl[20:0];
  assign nl_MultLoop_acc_4695_nl = ({(data_rsci_idat[629:612]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_4688[20:2]);
  assign MultLoop_acc_4695_nl = nl_MultLoop_acc_4695_nl[19:0];
  assign nl_MultLoop_acc_4473_nl = conv_s2u_15_19(readslicef_20_15_5((MultLoop_acc_4695_nl)))
      + conv_s2u_18_19(data_rsci_idat[629:612]);
  assign MultLoop_acc_4473_nl = nl_MultLoop_acc_4473_nl[18:0];
  assign nl_MultLoop_acc_3563_nl = conv_s2s_22_23({(~ (data_rsci_idat[521:504]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[521:504]));
  assign MultLoop_acc_3563_nl = nl_MultLoop_acc_3563_nl[22:0];
  assign nl_MultLoop_acc_173_nl = conv_s2s_23_24(MultLoop_acc_3563_nl) + ({(data_rsci_idat[521:504])
      , 6'b010000});
  assign MultLoop_acc_173_nl = nl_MultLoop_acc_173_nl[23:0];
  assign nl_MultLoop_acc_3565_nl = conv_s2s_22_23({(data_rsci_idat[467:450]) , 4'b0000})
      + conv_s2s_19_23(MultLoop_acc_3187_cse_1);
  assign MultLoop_acc_3565_nl = nl_MultLoop_acc_3565_nl[22:0];
  assign nl_MultLoop_acc_1132_nl = conv_s2u_23_25(MultLoop_acc_3565_nl) + conv_s2u_24_25({(data_rsci_idat[467:450])
      , 6'b000000});
  assign MultLoop_acc_1132_nl = nl_MultLoop_acc_1132_nl[24:0];
  assign nl_MultLoop_acc_3609_nl = conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1137_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4473_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_173_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1132_nl)));
  assign MultLoop_acc_3609_nl = nl_MultLoop_acc_3609_nl[17:0];
  assign nl_MultLoop_acc_3552_nl = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_15_19(data_rsci_idat[53:39]);
  assign MultLoop_acc_3552_nl = nl_MultLoop_acc_3552_nl[18:0];
  assign nl_MultLoop_acc_1122_nl = conv_s2u_19_21(MultLoop_acc_3552_nl) + conv_s2u_20_21({(data_rsci_idat[53:36])
      , 2'b00});
  assign MultLoop_acc_1122_nl = nl_MultLoop_acc_1122_nl[20:0];
  assign nl_MultLoop_acc_3557_nl = conv_s2s_18_19(data_rsci_idat[827:810]) + conv_s2s_13_19(data_rsci_idat[827:815]);
  assign MultLoop_acc_3557_nl = nl_MultLoop_acc_3557_nl[18:0];
  assign nl_MultLoop_acc_1140_nl = conv_s2u_19_22(MultLoop_acc_3557_nl) + conv_s2u_21_22({(data_rsci_idat[827:810])
      , 3'b000});
  assign MultLoop_acc_1140_nl = nl_MultLoop_acc_1140_nl[21:0];
  assign nl_MultLoop_acc_3558_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_14_18(data_rsci_idat[755:742]);
  assign MultLoop_acc_3558_nl = nl_MultLoop_acc_3558_nl[17:0];
  assign nl_MultLoop_acc_3559_nl = ({(data_rsci_idat[755:738]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3558_nl);
  assign MultLoop_acc_3559_nl = nl_MultLoop_acc_3559_nl[19:0];
  assign nl_MultLoop_acc_1138_nl = conv_s2u_20_23(MultLoop_acc_3559_nl) + conv_s2u_22_23({(data_rsci_idat[755:738])
      , 4'b0000});
  assign MultLoop_acc_1138_nl = nl_MultLoop_acc_1138_nl[22:0];
  assign nl_MultLoop_acc_4472_nl = conv_s2s_12_13(data_rsci_idat[71:60]) + 13'b0000000000001;
  assign MultLoop_acc_4472_nl = nl_MultLoop_acc_4472_nl[12:0];
  assign nl_MultLoop_acc_3554_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_16_18({(MultLoop_acc_4472_nl)
      , (data_rsci_idat[59:57])});
  assign MultLoop_acc_3554_nl = nl_MultLoop_acc_3554_nl[17:0];
  assign nl_MultLoop_acc_1123_nl = conv_s2u_18_22(MultLoop_acc_3554_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[71:54])) , 3'b001});
  assign MultLoop_acc_1123_nl = nl_MultLoop_acc_1123_nl[21:0];
  assign nl_MultLoop_acc_4651_nl = conv_s2u_18_21(MultLoop_acc_3556_itm_19_2_1) +
      ({(data_rsci_idat[35:18]) , 3'b001});
  assign MultLoop_acc_4651_nl = nl_MultLoop_acc_4651_nl[20:0];
  assign nl_MultLoop_acc_3614_itm_1  = (MultLoop_acc_3609_nl) + conv_s2s_16_18(MultLoop_acc_149_itm_23_8)
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1122_nl))) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1140_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1138_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1123_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_4651_nl)));
  assign nl_MultLoop_acc_3567_nl = ({(data_rsci_idat[269:252]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3063_cse_1);
  assign MultLoop_acc_3567_nl = nl_MultLoop_acc_3567_nl[19:0];
  assign nl_MultLoop_acc_1125_nl = conv_s2u_20_23(MultLoop_acc_3567_nl) + conv_s2u_22_23({(data_rsci_idat[269:252])
      , 4'b0000});
  assign MultLoop_acc_1125_nl = nl_MultLoop_acc_1125_nl[22:0];
  assign nl_MultLoop_acc_4474_nl = conv_s2u_15_19(MultLoop_acc_2026_itm_21_6[15:1])
      + conv_s2u_18_19(data_rsci_idat[233:216]);
  assign MultLoop_acc_4474_nl = nl_MultLoop_acc_4474_nl[18:0];
  assign nl_MultLoop_acc_3598_itm_1  = conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1125_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4474_nl)));
  assign nl_MultLoop_acc_188_nl = conv_s2u_13_18(data_rsci_idat[791:779]) - (data_rsci_idat[791:774]);
  assign MultLoop_acc_188_nl = nl_MultLoop_acc_188_nl[17:0];
  assign nl_MultLoop_acc_3504_nl = ({(data_rsci_idat[593:576]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_704_18_6
      , (~ (data_rsci_idat[581:576]))});
  assign MultLoop_acc_3504_nl = nl_MultLoop_acc_3504_nl[21:0];
  assign nl_MultLoop_acc_4476_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3504_nl)))
      + (~ (data_rsci_idat[593:576]));
  assign MultLoop_acc_4476_nl = nl_MultLoop_acc_4476_nl[17:0];
  assign nl_MultLoop_acc_1133_nl = conv_s2u_13_19(data_rsci_idat[485:473]) + conv_s2u_18_19(data_rsci_idat[485:468]);
  assign MultLoop_acc_1133_nl = nl_MultLoop_acc_1133_nl[18:0];
  assign nl_MultLoop_acc_3506_nl = (~ (data_rsci_idat[449:432])) + conv_s2s_16_18({MultLoop_MultLoop_conc_768_15_2
      , (data_rsci_idat[436:435])});
  assign MultLoop_acc_3506_nl = nl_MultLoop_acc_3506_nl[17:0];
  assign nl_MultLoop_acc_1131_nl = conv_s2u_18_21(MultLoop_acc_3506_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[449:432])) , 2'b01});
  assign MultLoop_acc_1131_nl = nl_MultLoop_acc_1131_nl[20:0];
  assign nl_MultLoop_acc_3584_itm_1  = conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_188_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4476_nl))) + conv_s2s_14_16(readslicef_19_14_5((MultLoop_acc_1133_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1131_nl)));
  assign nl_MultLoop_acc_3507_nl = (~ (data_rsci_idat[305:288])) + conv_s2s_14_18(data_rsci_idat[305:292]);
  assign MultLoop_acc_3507_nl = nl_MultLoop_acc_3507_nl[17:0];
  assign nl_MultLoop_acc_1127_nl = conv_s2u_18_20(MultLoop_acc_3507_nl) + ({(data_rsci_idat[305:288])
      , 2'b01});
  assign MultLoop_acc_1127_nl = nl_MultLoop_acc_1127_nl[19:0];
  assign nl_MultLoop_acc_4478_nl =  -conv_s2s_12_13(data_rsci_idat[251:240]);
  assign MultLoop_acc_4478_nl = nl_MultLoop_acc_4478_nl[12:0];
  assign nl_MultLoop_acc_3509_nl = ({(data_rsci_idat[251:234]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_4478_nl)
      , (~ (data_rsci_idat[239:234]))});
  assign MultLoop_acc_3509_nl = nl_MultLoop_acc_3509_nl[21:0];
  assign nl_MultLoop_acc_4479_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3509_nl)))
      + (~ (data_rsci_idat[251:234]));
  assign MultLoop_acc_4479_nl = nl_MultLoop_acc_4479_nl[17:0];
  assign nl_MultLoop_acc_4480_nl =  -conv_s2s_14_15(data_rsci_idat[161:148]);
  assign MultLoop_acc_4480_nl = nl_MultLoop_acc_4480_nl[14:0];
  assign nl_MultLoop_acc_153_nl = conv_s2s_19_23({(MultLoop_acc_4480_nl) , (~ (data_rsci_idat[147:144]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[161:144])) , 4'b0001});
  assign MultLoop_acc_153_nl = nl_MultLoop_acc_153_nl[22:0];
  assign nl_MultLoop_acc_3583_itm_1  = conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_1127_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4479_nl))) + conv_s2s_14_16(MultLoop_acc_3920_itm_17_2[15:2])
      + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_153_nl)));
  assign nl_MultLoop_acc_1141_nl = conv_s2u_18_23(MultLoop_acc_2375_cse_1) + conv_s2u_22_23({(~
      (data_rsci_idat[845:828])) , 4'b0001});
  assign MultLoop_acc_1141_nl = nl_MultLoop_acc_1141_nl[22:0];
  assign nl_MultLoop_acc_183_nl = conv_s2s_18_24(~ (data_rsci_idat[701:684])) + ({(data_rsci_idat[701:684])
      , 6'b000001});
  assign MultLoop_acc_183_nl = nl_MultLoop_acc_183_nl[23:0];
  assign nl_MultLoop_acc_4481_nl =  -conv_s2s_16_17(data_rsci_idat[395:380]);
  assign MultLoop_acc_4481_nl = nl_MultLoop_acc_4481_nl[16:0];
  assign nl_MultLoop_acc_166_nl = conv_s2s_19_21({(MultLoop_acc_4481_nl) , (~ (data_rsci_idat[379:378]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[395:378])) , 2'b01});
  assign MultLoop_acc_166_nl = nl_MultLoop_acc_166_nl[20:0];
  assign nl_MultLoop_acc_4482_nl = conv_s2s_9_10(MultLoop_acc_123_itm_17_3[14:6])
      + 10'b1111110001;
  assign MultLoop_acc_4482_nl = nl_MultLoop_acc_4482_nl[9:0];
  assign nl_MultLoop_acc_3571_nl = (readslicef_21_13_8((MultLoop_acc_166_nl))) +
      conv_s2s_12_13({(MultLoop_acc_4482_nl) , (MultLoop_acc_123_itm_17_3[5:4])});
  assign MultLoop_acc_3571_nl = nl_MultLoop_acc_3571_nl[12:0];
  assign nl_MultLoop_acc_3596_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1141_nl)))
      + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_183_nl))) + conv_s2s_15_17(MultLoop_acc_181_itm_22_8)
      + conv_s2s_14_17(MultLoop_acc_150_itm_17_4) + conv_s2s_13_17(MultLoop_acc_3571_nl);
  assign nl_MultLoop_acc_175_nl = conv_s2u_14_18(data_rsci_idat[557:544]) - (data_rsci_idat[557:540]);
  assign MultLoop_acc_175_nl = nl_MultLoop_acc_175_nl[17:0];
  assign nl_MultLoop_acc_4685_nl = conv_s2u_19_20(MultLoop_acc_2409_itm_20_2_1) +
      ({(data_rsci_idat[377:360]) , 2'b01});
  assign MultLoop_acc_4685_nl = nl_MultLoop_acc_4685_nl[19:0];
  assign nl_MultLoop_acc_3514_nl = (~ (data_rsci_idat[287:270])) + conv_s2s_13_18(data_rsci_idat[287:275]);
  assign MultLoop_acc_3514_nl = nl_MultLoop_acc_3514_nl[17:0];
  assign nl_MultLoop_acc_1126_nl = conv_s2u_18_20(MultLoop_acc_3514_nl) + ({(data_rsci_idat[287:270])
      , 2'b01});
  assign MultLoop_acc_1126_nl = nl_MultLoop_acc_1126_nl[19:0];
  assign nl_MultLoop_acc_3595_itm_1  = conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_175_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_4685_nl))) + conv_s2s_15_17(MultLoop_acc_1128_itm_21_7)
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1126_nl)));
  assign nl_MultLoop_acc_4652_nl = conv_s2u_19_20(MultLoop_acc_1722_cse_1[20:2])
      + ({(data_rsci_idat[17:0]) , 2'b01});
  assign MultLoop_acc_4652_nl = nl_MultLoop_acc_4652_nl[19:0];
  assign nl_MultLoop_acc_3577_nl = (readslicef_20_15_5((MultLoop_acc_4652_nl))) +
      conv_s2s_14_15(MultLoop_acc_4588_itm_18_2[16:3]);
  assign MultLoop_acc_3577_nl = nl_MultLoop_acc_3577_nl[14:0];
  assign nl_MultLoop_acc_3517_nl = ({(data_rsci_idat[197:180]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[197:180])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_698_18_7
      , (~ (data_rsci_idat[186:180]))});
  assign MultLoop_acc_3517_nl = nl_MultLoop_acc_3517_nl[22:0];
  assign nl_MultLoop_acc_4485_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3517_nl)))
      + (~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_4485_nl = nl_MultLoop_acc_4485_nl[17:0];
  assign nl_MultLoop_acc_3594_itm_1  = conv_s2s_15_17(MultLoop_acc_3577_nl) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4485_nl)))
      + conv_s2s_15_17(MultLoop_acc_1720_cse_1[20:6]);
  assign nl_MultLoop_acc_3519_nl = conv_s2s_21_22({(~ (data_rsci_idat[863:846]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_3519_nl = nl_MultLoop_acc_3519_nl[21:0];
  assign nl_MultLoop_acc_192_nl = conv_s2s_22_26(MultLoop_acc_3519_nl) + ({(data_rsci_idat[863:846])
      , 8'b00001000});
  assign MultLoop_acc_192_nl = nl_MultLoop_acc_192_nl[25:0];
  assign nl_MultLoop_acc_3523_nl = conv_s2s_24_25({(data_rsci_idat[773:756]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[773:756]) , 4'b0000}) + conv_s2s_20_25(MultLoop_acc_2520_cse_1);
  assign MultLoop_acc_3523_nl = nl_MultLoop_acc_3523_nl[24:0];
  assign nl_MultLoop_acc_4487_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_3523_nl)))
      + (~ (data_rsci_idat[773:756]));
  assign MultLoop_acc_4487_nl = nl_MultLoop_acc_4487_nl[17:0];
  assign nl_MultLoop_acc_3593_itm_1  = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_192_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4487_nl)));
  assign nl_MultLoop_acc_3525_nl = ({(data_rsci_idat[737:720]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_856_18_7
      , (~ (data_rsci_idat[726:720]))});
  assign MultLoop_acc_3525_nl = nl_MultLoop_acc_3525_nl[20:0];
  assign nl_MultLoop_acc_3526_nl = conv_s2s_23_24({(data_rsci_idat[737:720]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_3525_nl);
  assign MultLoop_acc_3526_nl = nl_MultLoop_acc_3526_nl[23:0];
  assign nl_MultLoop_acc_4489_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_3526_nl)))
      + (~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_4489_nl = nl_MultLoop_acc_4489_nl[17:0];
  assign nl_MultLoop_acc_3528_nl = (~ (data_rsci_idat[683:666])) + conv_s2s_17_18({MultLoop_MultLoop_conc_784_16_6
      , (data_rsci_idat[673:668])});
  assign MultLoop_acc_3528_nl = nl_MultLoop_acc_3528_nl[17:0];
  assign nl_MultLoop_acc_3529_nl = ({(data_rsci_idat[683:666]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3528_nl);
  assign MultLoop_acc_3529_nl = nl_MultLoop_acc_3529_nl[19:0];
  assign nl_MultLoop_acc_3530_nl = conv_s2s_22_23({(data_rsci_idat[683:666]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_3529_nl);
  assign MultLoop_acc_3530_nl = nl_MultLoop_acc_3530_nl[22:0];
  assign nl_MultLoop_acc_4491_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3530_nl)))
      + (~ (data_rsci_idat[683:666]));
  assign MultLoop_acc_4491_nl = nl_MultLoop_acc_4491_nl[17:0];
  assign nl_MultLoop_acc_4693_nl = conv_s2u_16_19(MultLoop_acc_3532_itm_20_5_1) +
      conv_s2u_18_19(data_rsci_idat[647:630]);
  assign MultLoop_acc_4693_nl = nl_MultLoop_acc_4693_nl[18:0];
  assign nl_MultLoop_acc_3534_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_16_18({MultLoop_MultLoop_conc_776_15_4
      , (data_rsci_idat[600:597])});
  assign MultLoop_acc_3534_nl = nl_MultLoop_acc_3534_nl[17:0];
  assign nl_MultLoop_acc_3535_nl = conv_s2s_20_21({(~ (data_rsci_idat[611:594]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3534_nl);
  assign MultLoop_acc_3535_nl = nl_MultLoop_acc_3535_nl[20:0];
  assign nl_MultLoop_acc_1135_nl = conv_s2u_21_23(MultLoop_acc_3535_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[611:594])) , 4'b0100});
  assign MultLoop_acc_1135_nl = nl_MultLoop_acc_1135_nl[22:0];
  assign nl_MultLoop_acc_3605_itm_1  = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4489_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4491_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4693_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1135_nl)));
  assign nl_MultLoop_acc_3546_nl = ({(data_rsci_idat[341:324]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_854_18_8
      , (~ (data_rsci_idat[331:324]))});
  assign MultLoop_acc_3546_nl = nl_MultLoop_acc_3546_nl[22:0];
  assign nl_MultLoop_acc_4496_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_3546_nl)))
      + (~ (data_rsci_idat[341:324]));
  assign MultLoop_acc_4496_nl = nl_MultLoop_acc_4496_nl[17:0];
  assign nl_MultLoop_acc_3548_nl = ({(data_rsci_idat[323:306]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_836_18_8
      , (~ (data_rsci_idat[313:306]))});
  assign MultLoop_acc_3548_nl = nl_MultLoop_acc_3548_nl[19:0];
  assign nl_MultLoop_acc_4498_nl = conv_s2u_12_18(readslicef_20_12_8((MultLoop_acc_3548_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_4498_nl = nl_MultLoop_acc_4498_nl[17:0];
  assign nl_MultLoop_acc_3536_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_13_18(data_rsci_idat[575:563]);
  assign MultLoop_acc_3536_nl = nl_MultLoop_acc_3536_nl[17:0];
  assign nl_MultLoop_acc_1134_nl = conv_s2u_18_20(MultLoop_acc_3536_nl) + ({(data_rsci_idat[575:558])
      , 2'b01});
  assign MultLoop_acc_1134_nl = nl_MultLoop_acc_1134_nl[19:0];
  assign nl_MultLoop_acc_3539_nl = conv_s2s_21_22({(data_rsci_idat[539:522]) , 3'b000})
      + conv_s2s_19_22(MultLoop_acc_2424_cse_1);
  assign MultLoop_acc_3539_nl = nl_MultLoop_acc_3539_nl[21:0];
  assign nl_MultLoop_acc_174_nl = conv_s2u_22_23(MultLoop_acc_3539_nl) + ({(~ (data_rsci_idat[539:522]))
      , 5'b00000});
  assign MultLoop_acc_174_nl = nl_MultLoop_acc_174_nl[22:0];
  assign nl_MultLoop_acc_3540_nl = (~ (data_rsci_idat[413:396])) + conv_s2s_14_18(data_rsci_idat[413:400]);
  assign MultLoop_acc_3540_nl = nl_MultLoop_acc_3540_nl[17:0];
  assign nl_MultLoop_acc_3541_nl = conv_s2s_20_21({(~ (data_rsci_idat[413:396]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3540_nl);
  assign MultLoop_acc_3541_nl = nl_MultLoop_acc_3541_nl[20:0];
  assign nl_MultLoop_acc_1129_nl = conv_s2u_21_22(MultLoop_acc_3541_nl) + ({(data_rsci_idat[413:396])
      , 4'b0100});
  assign MultLoop_acc_1129_nl = nl_MultLoop_acc_1129_nl[21:0];
  assign nl_MultLoop_acc_3543_nl = (~ (data_rsci_idat[431:414])) + conv_s2s_17_18({MultLoop_MultLoop_conc_794_16_5
      , (data_rsci_idat[420:416])});
  assign MultLoop_acc_3543_nl = nl_MultLoop_acc_3543_nl[17:0];
  assign nl_MultLoop_acc_3544_nl = conv_s2s_20_21({(~ (data_rsci_idat[431:414]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3543_nl);
  assign MultLoop_acc_3544_nl = nl_MultLoop_acc_3544_nl[20:0];
  assign nl_MultLoop_acc_1130_nl = conv_s2u_21_24(MultLoop_acc_3544_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[431:414])) , 5'b00100});
  assign MultLoop_acc_1130_nl = nl_MultLoop_acc_1130_nl[23:0];
  assign nl_MultLoop_acc_3550_nl = ({(data_rsci_idat[179:162]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_826_18_5
      , (~ (data_rsci_idat[166:162]))});
  assign MultLoop_acc_3550_nl = nl_MultLoop_acc_3550_nl[20:0];
  assign nl_MultLoop_acc_154_nl = conv_s2s_21_23(MultLoop_acc_3550_nl) + ({(~ (data_rsci_idat[179:162]))
      , 5'b00000});
  assign MultLoop_acc_154_nl = nl_MultLoop_acc_154_nl[22:0];
  assign nl_MultLoop_acc_1124_nl = conv_s2u_18_21(MultLoop_acc_2079_cse_1) + ({(data_rsci_idat[125:108])
      , 3'b001});
  assign MultLoop_acc_1124_nl = nl_MultLoop_acc_1124_nl[20:0];
  assign nl_MultLoop_acc_3611_itm_1  = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4496_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4498_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1134_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_174_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1129_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1130_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_154_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1124_nl)));
  assign nl_MultLoop_acc_1992_nl = ({(~ (data_rsci_idat[863:846])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[863:846])
      + conv_s2s_16_21({MultLoop_acc_4011_cse_1 , (data_rsci_idat[853:849])});
  assign MultLoop_acc_1992_nl = nl_MultLoop_acc_1992_nl[20:0];
  assign nl_MultLoop_acc_1401_nl = conv_s2u_21_24(MultLoop_acc_1992_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[863:846])) , 5'b01000});
  assign MultLoop_acc_1401_nl = nl_MultLoop_acc_1401_nl[23:0];
  assign nl_MultLoop_acc_4603_nl = conv_s2u_16_19(MultLoop_acc_1993_itm_18_2[16:1])
      + conv_s2u_18_19(data_rsci_idat[683:666]);
  assign MultLoop_acc_4603_nl = nl_MultLoop_acc_4603_nl[18:0];
  assign nl_MultLoop_acc_1983_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_13_18(data_rsci_idat[125:113]);
  assign MultLoop_acc_1983_nl = nl_MultLoop_acc_1983_nl[17:0];
  assign nl_MultLoop_acc_1385_nl = conv_s2u_18_20(MultLoop_acc_1983_nl) + ({(data_rsci_idat[125:108])
      , 2'b01});
  assign MultLoop_acc_1385_nl = nl_MultLoop_acc_1385_nl[19:0];
  assign nl_MultLoop_acc_4004_nl =  -conv_s2s_10_11(data_rsci_idat[107:98]);
  assign MultLoop_acc_4004_nl = nl_MultLoop_acc_4004_nl[10:0];
  assign nl_MultLoop_acc_1986_nl = ({(data_rsci_idat[107:90]) , 6'b001000}) + conv_s2s_21_24({(~
      (data_rsci_idat[107:90])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4004_nl)
      , (~ (data_rsci_idat[97:90]))});
  assign MultLoop_acc_1986_nl = nl_MultLoop_acc_1986_nl[23:0];
  assign nl_MultLoop_acc_4005_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_1986_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_4005_nl = nl_MultLoop_acc_4005_nl[17:0];
  assign nl_MultLoop_acc_4006_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_17_18(MultLoop_acc_4594_itm_18_2);
  assign MultLoop_acc_4006_nl = nl_MultLoop_acc_4006_nl[17:0];
  assign nl_MultLoop_acc_4007_nl = conv_s2u_18_20(MultLoop_acc_4006_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign MultLoop_acc_4007_nl = nl_MultLoop_acc_4007_nl[19:0];
  assign nl_MultLoop_acc_4009_nl =  -conv_s2s_12_13(data_rsci_idat[845:834]);
  assign MultLoop_acc_4009_nl = nl_MultLoop_acc_4009_nl[12:0];
  assign nl_MultLoop_acc_1929_nl = ({(data_rsci_idat[845:828]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4009_nl)
      , (~ (data_rsci_idat[833:828]))});
  assign MultLoop_acc_1929_nl = nl_MultLoop_acc_1929_nl[20:0];
  assign nl_MultLoop_acc_4010_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_1929_nl)))
      + (~ (data_rsci_idat[845:828]));
  assign MultLoop_acc_4010_nl = nl_MultLoop_acc_4010_nl[17:0];
  assign nl_MultLoop_acc_1927_nl = conv_s2s_18_19(data_rsci_idat[485:468]) + conv_s2s_16_19({MultLoop_MultLoop_conc_810_15_2
      , (data_rsci_idat[472:471])});
  assign MultLoop_acc_1927_nl = nl_MultLoop_acc_1927_nl[18:0];
  assign nl_MultLoop_acc_927_nl = conv_s2u_19_20(MultLoop_acc_1927_nl) + ({(~ (data_rsci_idat[485:468]))
      , 2'b00});
  assign MultLoop_acc_927_nl = nl_MultLoop_acc_927_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_50_itm_1  =
      conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1401_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4603_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1385_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4005_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_4007_nl))) + conv_s2s_14_18(readslicef_18_14_4((MultLoop_acc_4010_nl)))
      + conv_s2s_13_18(Result_acc_127_cse_1[18:6]) + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_927_nl)));
  assign nl_MultLoop_acc_4012_nl =  -conv_s2s_10_11(data_rsci_idat[593:584]);
  assign MultLoop_acc_4012_nl = nl_MultLoop_acc_4012_nl[10:0];
  assign nl_MultLoop_acc_933_nl = conv_s2s_26_27({(~ (data_rsci_idat[593:576])) ,
      8'b00001000}) + conv_s2s_21_27({(~ (data_rsci_idat[593:576])) , 3'b001}) +
      conv_s2s_19_27({(MultLoop_acc_4012_nl) , (~ (data_rsci_idat[583:576]))});
  assign MultLoop_acc_933_nl = nl_MultLoop_acc_933_nl[26:0];
  assign nl_MultLoop_acc_4013_nl =  -conv_s2s_13_14(data_rsci_idat[359:347]);
  assign MultLoop_acc_4013_nl = nl_MultLoop_acc_4013_nl[13:0];
  assign nl_MultLoop_acc_920_nl = conv_s2s_23_24({(~ (data_rsci_idat[359:342])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[359:342])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4013_nl)
      , (~ (data_rsci_idat[346:342]))});
  assign MultLoop_acc_920_nl = nl_MultLoop_acc_920_nl[23:0];
  assign nl_MultLoop_acc_1999_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1844_cse_1);
  assign MultLoop_acc_1999_nl = nl_MultLoop_acc_1999_nl[19:0];
  assign nl_MultLoop_acc_1386_nl = conv_s2u_20_23(MultLoop_acc_1999_nl) + conv_s2u_22_23({(data_rsci_idat[161:144])
      , 4'b0000});
  assign MultLoop_acc_1386_nl = nl_MultLoop_acc_1386_nl[22:0];
  assign nl_MultLoop_acc_910_nl = conv_s2s_26_27({(~ (data_rsci_idat[179:162])) ,
      8'b00010000}) + conv_s2s_22_27({(~ (data_rsci_idat[179:162])) , 4'b0100}) +
      conv_s2s_20_27({(~ (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_27({MultLoop_MultLoop_conc_718_18_8
      , (~ (data_rsci_idat[169:162]))});
  assign MultLoop_acc_910_nl = nl_MultLoop_acc_910_nl[26:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_49_itm_1  =
      conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_933_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_920_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1386_nl))) + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_910_nl)));
  assign nl_MultLoop_acc_2003_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[35:18]));
  assign MultLoop_acc_2003_nl = nl_MultLoop_acc_2003_nl[19:0];
  assign nl_MultLoop_acc_2004_nl = ({(~ (data_rsci_idat[35:18])) , 5'b00000}) + conv_s2s_20_23(MultLoop_acc_2003_nl);
  assign MultLoop_acc_2004_nl = nl_MultLoop_acc_2004_nl[22:0];
  assign nl_MultLoop_acc_903_nl = conv_s2s_23_25(MultLoop_acc_2004_nl) + ({(data_rsci_idat[35:18])
      , 7'b0100000});
  assign MultLoop_acc_903_nl = nl_MultLoop_acc_903_nl[24:0];
  assign nl_MultLoop_acc_2007_nl = (readslicef_25_15_10((MultLoop_acc_903_nl))) +
      15'b000000011101011;
  assign MultLoop_acc_2007_nl = nl_MultLoop_acc_2007_nl[14:0];
  assign nl_MultLoop_acc_2006_nl = (~ (data_rsci_idat[17:0])) + conv_s2s_13_18({MultLoop_acc_4015_cse_1
      , (data_rsci_idat[7:6])});
  assign MultLoop_acc_2006_nl = nl_MultLoop_acc_2006_nl[17:0];
  assign nl_MultLoop_acc_902_nl = conv_s2u_18_21(MultLoop_acc_2006_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[17:0])) , 2'b01});
  assign MultLoop_acc_902_nl = nl_MultLoop_acc_902_nl[20:0];
  assign nl_MultLoop_914_MultLoop_acc_3_nl = conv_s2s_15_17(MultLoop_acc_2007_nl)
      + (readslicef_21_17_4((MultLoop_acc_902_nl)));
  assign MultLoop_914_MultLoop_acc_3_nl = nl_MultLoop_914_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_4016_nl =  -conv_s2s_14_15(data_rsci_idat[611:598]);
  assign MultLoop_acc_4016_nl = nl_MultLoop_acc_4016_nl[14:0];
  assign nl_MultLoop_acc_934_nl = conv_s2s_19_23({(MultLoop_acc_4016_nl) , (~ (data_rsci_idat[597:594]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[611:594])) , 4'b0001});
  assign MultLoop_acc_934_nl = nl_MultLoop_acc_934_nl[22:0];
  assign nl_MultLoop_acc_1931_nl = conv_s2s_18_19(data_rsci_idat[449:432]) + conv_s2s_15_19(data_rsci_idat[449:435]);
  assign MultLoop_acc_1931_nl = nl_MultLoop_acc_1931_nl[18:0];
  assign nl_MultLoop_acc_1392_nl = conv_s2u_19_21(MultLoop_acc_1931_nl) + conv_s2u_20_21({(data_rsci_idat[449:432])
      , 2'b00});
  assign MultLoop_acc_1392_nl = nl_MultLoop_acc_1392_nl[20:0];
  assign nl_MultLoop_acc_4017_nl =  -conv_s2s_13_14(data_rsci_idat[377:365]);
  assign MultLoop_acc_4017_nl = nl_MultLoop_acc_4017_nl[13:0];
  assign nl_MultLoop_acc_921_nl = conv_s2s_23_24({(~ (data_rsci_idat[377:360])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[377:360])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4017_nl)
      , (~ (data_rsci_idat[364:360]))});
  assign MultLoop_acc_921_nl = nl_MultLoop_acc_921_nl[23:0];
  assign nl_MultLoop_acc_4018_nl =  -conv_s2s_16_17(data_rsci_idat[305:290]);
  assign MultLoop_acc_4018_nl = nl_MultLoop_acc_4018_nl[16:0];
  assign nl_MultLoop_acc_917_nl = conv_s2s_19_21({(MultLoop_acc_4018_nl) , (~ (data_rsci_idat[289:288]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[305:288])) , 2'b01});
  assign MultLoop_acc_917_nl = nl_MultLoop_acc_917_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_38_itm_1  =
      conv_s2s_17_18(MultLoop_914_MultLoop_acc_3_nl) + conv_s2s_14_18(readslicef_23_14_9((MultLoop_acc_934_nl)))
      + conv_s2s_14_18(readslicef_21_14_7((MultLoop_acc_1392_nl))) + conv_s2s_14_18(readslicef_24_14_10((MultLoop_acc_921_nl)))
      + conv_s2s_14_18(readslicef_21_14_7((MultLoop_acc_917_nl)));
  assign nl_MultLoop_acc_4604_nl = conv_s2u_15_19(MultLoop_acc_1940_cse_1[19:5])
      + conv_s2u_18_19(data_rsci_idat[701:684]);
  assign MultLoop_acc_4604_nl = nl_MultLoop_acc_4604_nl[18:0];
  assign nl_MultLoop_acc_1936_nl = ({(data_rsci_idat[233:216]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_702_18_6
      , (~ (data_rsci_idat[221:216]))});
  assign MultLoop_acc_1936_nl = nl_MultLoop_acc_1936_nl[19:0];
  assign nl_MultLoop_acc_1937_nl = conv_s2s_22_23({(data_rsci_idat[233:216]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_1936_nl);
  assign MultLoop_acc_1937_nl = nl_MultLoop_acc_1937_nl[22:0];
  assign nl_MultLoop_acc_4020_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_1937_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_4020_nl = nl_MultLoop_acc_4020_nl[17:0];
  assign nl_MultLoop_acc_1939_nl = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_15_19({MultLoop_acc_4021_cse_1
      , (data_rsci_idat[131:130])});
  assign MultLoop_acc_1939_nl = nl_MultLoop_acc_1939_nl[18:0];
  assign nl_MultLoop_acc_908_nl = conv_s2u_19_20(MultLoop_acc_1939_nl) + ({(~ (data_rsci_idat[143:126]))
      , 2'b00});
  assign MultLoop_acc_908_nl = nl_MultLoop_acc_908_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_23_itm_1  =
      conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_4604_nl))) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4020_nl)))
      + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_908_nl)));
  assign nl_MultLoop_acc_4022_nl =  -conv_s2s_14_15(data_rsci_idat[665:652]);
  assign MultLoop_acc_4022_nl = nl_MultLoop_acc_4022_nl[14:0];
  assign nl_MultLoop_acc_937_nl = conv_s2s_22_23({(~ (data_rsci_idat[665:648])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[665:648])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_4022_nl)
      , (~ (data_rsci_idat[651:648]))});
  assign MultLoop_acc_937_nl = nl_MultLoop_acc_937_nl[22:0];
  assign nl_MultLoop_acc_4605_nl = conv_s2u_17_19(MultLoop_acc_1943_itm_18_2) + conv_s2u_18_19(data_rsci_idat[629:612]);
  assign MultLoop_acc_4605_nl = nl_MultLoop_acc_4605_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_22_itm_1  =
      conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_937_nl))) + conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_4605_nl)));
  assign nl_MultLoop_acc_1384_nl = conv_s2u_12_19(data_rsci_idat[89:78]) + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_1384_nl = nl_MultLoop_acc_1384_nl[18:0];
  assign nl_MultLoop_acc_1400_nl = conv_s2u_15_19(data_rsci_idat[827:813]) + conv_s2u_18_19(data_rsci_idat[827:810]);
  assign MultLoop_acc_1400_nl = nl_MultLoop_acc_1400_nl[18:0];
  assign nl_MultLoop_acc_945_nl = conv_s2u_15_18(data_rsci_idat[809:795]) - (data_rsci_idat[809:792]);
  assign MultLoop_acc_945_nl = nl_MultLoop_acc_945_nl[17:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_8_nl = ~((data_rsci_idat[62:54]!=9'b000000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = conv_s2s_11_12(readslicef_18_11_7((MultLoop_acc_945_nl)))
      + conv_s2s_9_12(~ (data_rsci_idat[71:63])) + conv_u2s_1_12(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_8_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl[11:0];
  assign nl_MultLoop_acc_918_nl = conv_s2u_16_18(data_rsci_idat[323:308]) - (data_rsci_idat[323:306]);
  assign MultLoop_acc_918_nl = nl_MultLoop_acc_918_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl = conv_s2s_13_14(readslicef_19_13_6((MultLoop_acc_1400_nl)))
      + conv_s2s_12_14(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_12_nl)
      + conv_s2s_12_14(readslicef_18_12_6((MultLoop_acc_918_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl[13:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl = (readslicef_19_15_4((MultLoop_acc_1384_nl)))
      + conv_s2s_14_15(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_15_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl[14:0];
  assign nl_MultLoop_acc_1945_nl = (~ (data_rsci_idat[773:756])) + conv_s2s_14_18(data_rsci_idat[773:760]);
  assign MultLoop_acc_1945_nl = nl_MultLoop_acc_1945_nl[17:0];
  assign nl_MultLoop_acc_1398_nl = conv_s2u_18_20(MultLoop_acc_1945_nl) + ({(data_rsci_idat[773:756])
      , 2'b01});
  assign MultLoop_acc_1398_nl = nl_MultLoop_acc_1398_nl[19:0];
  assign nl_MultLoop_acc_1947_nl = conv_s2s_20_21({(~ (data_rsci_idat[791:774]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1946_cse_1);
  assign MultLoop_acc_1947_nl = nl_MultLoop_acc_1947_nl[20:0];
  assign nl_MultLoop_acc_1399_nl = conv_s2u_21_22(MultLoop_acc_1947_nl) + ({(data_rsci_idat[791:774])
      , 4'b0100});
  assign MultLoop_acc_1399_nl = nl_MultLoop_acc_1399_nl[21:0];
  assign nl_MultLoop_acc_1944_nl = conv_s2s_18_19(data_rsci_idat[215:198]) + conv_s2s_15_19(data_rsci_idat[215:201]);
  assign MultLoop_acc_1944_nl = nl_MultLoop_acc_1944_nl[18:0];
  assign nl_MultLoop_acc_1387_nl = conv_s2u_19_22(MultLoop_acc_1944_nl) + conv_s2u_21_22({(data_rsci_idat[215:198])
      , 3'b000});
  assign MultLoop_acc_1387_nl = nl_MultLoop_acc_1387_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_47_itm_1  =
      conv_s2s_15_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_20_nl)
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1398_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1399_nl)))
      + conv_s2s_15_18(MultLoop_acc_1275_itm_20_5[15:1]) + conv_s2s_15_18(readslicef_22_15_7((MultLoop_acc_1387_nl)));
  assign nl_MultLoop_acc_1951_nl = ({(data_rsci_idat[737:720]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[737:720])) , 4'b0100}) + conv_s2s_21_24(MultLoop_acc_1949_cse_1);
  assign MultLoop_acc_1951_nl = nl_MultLoop_acc_1951_nl[23:0];
  assign nl_MultLoop_acc_4024_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_1951_nl)))
      + (~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_4024_nl = nl_MultLoop_acc_4024_nl[17:0];
  assign nl_MultLoop_acc_1952_nl = ({(data_rsci_idat[755:738]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[755:738]));
  assign MultLoop_acc_1952_nl = nl_MultLoop_acc_1952_nl[19:0];
  assign nl_MultLoop_acc_942_nl = conv_s2s_24_25({(data_rsci_idat[755:738]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[755:738]) , 4'b0000}) + conv_s2s_20_25(MultLoop_acc_1952_nl);
  assign MultLoop_acc_942_nl = nl_MultLoop_acc_942_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_34_itm_1  =
      conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4024_nl))) + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_942_nl)));
  assign nl_MultLoop_acc_1954_nl = (~ (data_rsci_idat[719:702])) + conv_s2s_16_18(data_rsci_idat[719:704]);
  assign MultLoop_acc_1954_nl = nl_MultLoop_acc_1954_nl[17:0];
  assign nl_MultLoop_acc_1955_nl = conv_s2s_20_21({(~ (data_rsci_idat[719:702]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1954_nl);
  assign MultLoop_acc_1955_nl = nl_MultLoop_acc_1955_nl[20:0];
  assign nl_MultLoop_acc_1397_nl = conv_s2u_21_23(MultLoop_acc_1955_nl) + ({(data_rsci_idat[719:702])
      , 5'b00100});
  assign MultLoop_acc_1397_nl = nl_MultLoop_acc_1397_nl[22:0];
  assign nl_MultLoop_acc_936_nl = conv_s2s_24_25({(~ (data_rsci_idat[647:630])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[647:630])) , 4'b0100}) + conv_s2s_21_25(MultLoop_acc_1957_cse_1);
  assign MultLoop_acc_936_nl = nl_MultLoop_acc_936_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_33_itm_1  =
      conv_s2s_16_17(readslicef_23_16_7((MultLoop_acc_1397_nl))) + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_936_nl)));
  assign nl_MultLoop_acc_931_nl = conv_s2s_19_26({MultLoop_MultLoop_conc_700_18_7
      , (~ (data_rsci_idat[546:540]))}) + conv_s2s_25_26({(~ (data_rsci_idat[557:540]))
      , 7'b0000001});
  assign MultLoop_acc_931_nl = nl_MultLoop_acc_931_nl[25:0];
  assign nl_MultLoop_acc_1961_nl = ({(data_rsci_idat[521:504]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_726_18_7
      , (~ (data_rsci_idat[510:504]))});
  assign MultLoop_acc_1961_nl = nl_MultLoop_acc_1961_nl[19:0];
  assign nl_MultLoop_acc_4028_nl = conv_s2u_13_18(readslicef_20_13_7((MultLoop_acc_1961_nl)))
      + (~ (data_rsci_idat[521:504]));
  assign MultLoop_acc_4028_nl = nl_MultLoop_acc_4028_nl[17:0];
  assign nl_MultLoop_acc_4606_nl = conv_s2u_16_19(MultLoop_acc_1962_cse_1[18:3])
      + conv_s2u_18_19(data_rsci_idat[539:522]);
  assign MultLoop_acc_4606_nl = nl_MultLoop_acc_4606_nl[18:0];
  assign nl_MultLoop_acc_4029_nl = conv_s2s_11_12(data_rsci_idat[503:493]) + 12'b000000000001;
  assign MultLoop_acc_4029_nl = nl_MultLoop_acc_4029_nl[11:0];
  assign nl_MultLoop_acc_1964_nl = (~ (data_rsci_idat[503:486])) + conv_s2s_17_18({(MultLoop_acc_4029_nl)
      , (data_rsci_idat[492:488])});
  assign MultLoop_acc_1964_nl = nl_MultLoop_acc_1964_nl[17:0];
  assign nl_MultLoop_acc_1965_nl = ({(data_rsci_idat[503:486]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1964_nl);
  assign MultLoop_acc_1965_nl = nl_MultLoop_acc_1965_nl[19:0];
  assign nl_MultLoop_acc_928_nl = conv_s2u_20_23(MultLoop_acc_1965_nl) + ({(~ (data_rsci_idat[503:486]))
      , 5'b00000});
  assign MultLoop_acc_928_nl = nl_MultLoop_acc_928_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_45_itm_1  =
      conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_931_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4028_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4606_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_928_nl)));
  assign nl_MultLoop_acc_1977_nl = (~ (data_rsci_idat[341:324])) + conv_s2s_12_18(data_rsci_idat[341:330]);
  assign MultLoop_acc_1977_nl = nl_MultLoop_acc_1977_nl[17:0];
  assign nl_MultLoop_acc_1391_nl = conv_s2u_18_20(MultLoop_acc_1977_nl) + ({(data_rsci_idat[341:324])
      , 2'b01});
  assign MultLoop_acc_1391_nl = nl_MultLoop_acc_1391_nl[19:0];
  assign nl_MultLoop_acc_1979_nl = conv_s2s_20_21({(~ (data_rsci_idat[287:270]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_1626_cse_1);
  assign MultLoop_acc_1979_nl = nl_MultLoop_acc_1979_nl[20:0];
  assign nl_MultLoop_acc_1390_nl = conv_s2u_21_22(MultLoop_acc_1979_nl) + ({(data_rsci_idat[287:270])
      , 4'b0100});
  assign MultLoop_acc_1390_nl = nl_MultLoop_acc_1390_nl[21:0];
  assign nl_MultLoop_acc_1967_nl = (~ (data_rsci_idat[467:450])) + conv_s2s_17_18({MultLoop_acc_4030_cse_1
      , (data_rsci_idat[457:452])});
  assign MultLoop_acc_1967_nl = nl_MultLoop_acc_1967_nl[17:0];
  assign nl_MultLoop_acc_1968_nl = ({(data_rsci_idat[467:450]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_1967_nl);
  assign MultLoop_acc_1968_nl = nl_MultLoop_acc_1968_nl[19:0];
  assign nl_MultLoop_acc_1969_nl = conv_s2s_22_23({(data_rsci_idat[467:450]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_1968_nl);
  assign MultLoop_acc_1969_nl = nl_MultLoop_acc_1969_nl[22:0];
  assign nl_MultLoop_acc_4031_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_1969_nl)))
      + (~ (data_rsci_idat[467:450]));
  assign MultLoop_acc_4031_nl = nl_MultLoop_acc_4031_nl[17:0];
  assign nl_MultLoop_acc_1971_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_16_19({MultLoop_acc_4032_cse_1
      , (data_rsci_idat[400:399])});
  assign MultLoop_acc_1971_nl = nl_MultLoop_acc_1971_nl[18:0];
  assign nl_MultLoop_acc_923_nl = conv_s2u_19_20(MultLoop_acc_1971_nl) + ({(~ (data_rsci_idat[413:396]))
      , 2'b00});
  assign MultLoop_acc_923_nl = nl_MultLoop_acc_923_nl[19:0];
  assign nl_MultLoop_acc_1973_nl = ({(data_rsci_idat[431:414]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_844_18_7
      , (~ (data_rsci_idat[420:414]))});
  assign MultLoop_acc_1973_nl = nl_MultLoop_acc_1973_nl[20:0];
  assign nl_MultLoop_acc_1974_nl = conv_s2s_23_24({(data_rsci_idat[431:414]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_1973_nl);
  assign MultLoop_acc_1974_nl = nl_MultLoop_acc_1974_nl[23:0];
  assign nl_MultLoop_acc_4034_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_1974_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_4034_nl = nl_MultLoop_acc_4034_nl[17:0];
  assign nl_MultLoop_acc_922_nl = conv_s2s_25_26({(~ (data_rsci_idat[395:378])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[395:378])) , 5'b00001}) +
      conv_s2s_19_26({MultLoop_MultLoop_conc_818_18_7 , (~ (data_rsci_idat[384:378]))});
  assign MultLoop_acc_922_nl = nl_MultLoop_acc_922_nl[25:0];
  assign nl_MultLoop_acc_1980_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_13_18(data_rsci_idat[251:239]);
  assign MultLoop_acc_1980_nl = nl_MultLoop_acc_1980_nl[17:0];
  assign nl_MultLoop_acc_1388_nl = conv_s2u_18_21(MultLoop_acc_1980_nl) + ({(data_rsci_idat[251:234])
      , 3'b001});
  assign MultLoop_acc_1388_nl = nl_MultLoop_acc_1388_nl[20:0];
  assign nl_MultLoop_acc_1982_nl = conv_s2s_18_19(data_rsci_idat[197:180]) + conv_s2s_17_19({MultLoop_acc_4036_cse_1
      , (data_rsci_idat[186:182])});
  assign MultLoop_acc_1982_nl = nl_MultLoop_acc_1982_nl[18:0];
  assign nl_MultLoop_acc_911_nl = conv_s2u_19_23(MultLoop_acc_1982_nl) + ({(~ (data_rsci_idat[197:180]))
      , 5'b00000});
  assign MultLoop_acc_911_nl = nl_MultLoop_acc_911_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_51_itm_1  =
      conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1391_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1390_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4031_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_923_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4034_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_922_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1388_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_911_nl)));
  assign nl_MultLoop_acc_4442_nl = conv_s2s_14_15(data_rsci_idat[35:22]) + 15'b000000000000001;
  assign MultLoop_acc_4442_nl = nl_MultLoop_acc_4442_nl[14:0];
  assign nl_MultLoop_acc_3386_nl = (~ (data_rsci_idat[35:18])) + conv_s2s_17_18({(MultLoop_acc_4442_nl)
      , (data_rsci_idat[21:20])});
  assign MultLoop_acc_3386_nl = nl_MultLoop_acc_3386_nl[17:0];
  assign nl_MultLoop_acc_1142_nl = conv_s2u_18_21(MultLoop_acc_3386_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[35:18])) , 2'b01});
  assign MultLoop_acc_1142_nl = nl_MultLoop_acc_1142_nl[20:0];
  assign nl_MultLoop_acc_3456_nl = (readslicef_21_13_8((MultLoop_acc_1142_nl))) +
      conv_s2s_12_13(MultLoop_acc_1152_itm_18_3[15:4]);
  assign MultLoop_acc_3456_nl = nl_MultLoop_acc_3456_nl[12:0];
  assign nl_MultLoop_acc_3470_nl = (MultLoop_acc_2807_itm_18_2[16:1]) + conv_s2s_13_16(MultLoop_acc_3456_nl)
      + conv_s2s_13_16(MultLoop_acc_1543_itm_21_6[15:3]) + conv_s2s_13_16(MultLoop_acc_181_itm_22_8[14:2]);
  assign MultLoop_acc_3470_nl = nl_MultLoop_acc_3470_nl[15:0];
  assign nl_MultLoop_acc_4443_nl = conv_s2s_10_11(data_rsci_idat[809:800]) + 11'b00000000001;
  assign MultLoop_acc_4443_nl = nl_MultLoop_acc_4443_nl[10:0];
  assign nl_MultLoop_acc_3444_nl = ({(~ (data_rsci_idat[809:792])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[809:792])
      + conv_s2s_17_20({(MultLoop_acc_4443_nl) , (data_rsci_idat[799:794])});
  assign MultLoop_acc_3444_nl = nl_MultLoop_acc_3444_nl[19:0];
  assign nl_MultLoop_acc_1158_nl = conv_s2u_20_25(MultLoop_acc_3444_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[809:792])) , 6'b000100});
  assign MultLoop_acc_1158_nl = nl_MultLoop_acc_1158_nl[24:0];
  assign nl_MultLoop_acc_3446_nl = ({(data_rsci_idat[647:630]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2568_cse_1);
  assign MultLoop_acc_3446_nl = nl_MultLoop_acc_3446_nl[19:0];
  assign nl_MultLoop_acc_1155_nl = conv_s2u_20_25(MultLoop_acc_3446_nl) + conv_s2u_24_25({(data_rsci_idat[647:630])
      , 6'b000000});
  assign MultLoop_acc_1155_nl = nl_MultLoop_acc_1155_nl[24:0];
  assign nl_MultLoop_acc_3439_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[89:72]));
  assign MultLoop_acc_3439_nl = nl_MultLoop_acc_3439_nl[19:0];
  assign nl_MultLoop_acc_197_nl = conv_s2s_20_23(MultLoop_acc_3439_nl) + conv_s2s_22_23({(data_rsci_idat[89:72])
      , 4'b0000});
  assign MultLoop_acc_197_nl = nl_MultLoop_acc_197_nl[22:0];
  assign nl_MultLoop_acc_4441_nl = conv_s2u_16_19(MultLoop_acc_434_itm_22_7) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_4441_nl = nl_MultLoop_acc_4441_nl[18:0];
  assign nl_MultLoop_acc_3495_itm_1  = conv_s2s_16_18(MultLoop_acc_3470_nl) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1158_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1155_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_197_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4441_nl)));
  assign nl_MultLoop_acc_3448_nl = (~ (data_rsci_idat[341:324])) + conv_s2s_16_18({MultLoop_acc_4122_cse_1
      , (data_rsci_idat[331:327])});
  assign MultLoop_acc_3448_nl = nl_MultLoop_acc_3448_nl[17:0];
  assign nl_MultLoop_acc_3449_nl = conv_s2s_21_22({(~ (data_rsci_idat[341:324]))
      , 3'b001}) + conv_s2s_18_22(MultLoop_acc_3448_nl);
  assign MultLoop_acc_3449_nl = nl_MultLoop_acc_3449_nl[21:0];
  assign nl_MultLoop_acc_1148_nl = conv_s2u_22_24(MultLoop_acc_3449_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[341:324])) , 5'b01000});
  assign MultLoop_acc_1148_nl = nl_MultLoop_acc_1148_nl[23:0];
  assign nl_MultLoop_acc_4445_nl =  -conv_s2s_10_11(data_rsci_idat[359:350]);
  assign MultLoop_acc_4445_nl = nl_MultLoop_acc_4445_nl[10:0];
  assign nl_MultLoop_acc_212_nl = conv_s2s_26_27({(~ (data_rsci_idat[359:342])) ,
      8'b00001000}) + conv_s2s_21_27({(~ (data_rsci_idat[359:342])) , 3'b001}) +
      conv_s2s_19_27({(MultLoop_acc_4445_nl) , (~ (data_rsci_idat[349:342]))});
  assign MultLoop_acc_212_nl = nl_MultLoop_acc_212_nl[26:0];
  assign nl_MultLoop_acc_204_nl = conv_s2s_26_27({(~ (data_rsci_idat[215:198])) ,
      8'b00100000}) + conv_s2s_23_27({(~ (data_rsci_idat[215:198])) , 5'b00100})
      + conv_s2s_20_27({(~ (data_rsci_idat[215:198])) , 2'b01}) + conv_s2s_19_27({MultLoop_MultLoop_conc_746_18_8
      , (~ (data_rsci_idat[205:198]))});
  assign MultLoop_acc_204_nl = nl_MultLoop_acc_204_nl[26:0];
  assign nl_MultLoop_acc_200_nl = conv_s2s_19_25({MultLoop_MultLoop_conc_824_18_6
      , (~ (data_rsci_idat[131:126]))}) + conv_s2s_24_25({(~ (data_rsci_idat[143:126]))
      , 6'b000001});
  assign MultLoop_acc_200_nl = nl_MultLoop_acc_200_nl[24:0];
  assign nl_MultLoop_acc_3494_itm_1  = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1148_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_212_nl))) + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_204_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_200_nl)));
  assign nl_MultLoop_acc_4684_nl = conv_s2u_15_18(MultLoop_acc_1822_cse_1[18:4])
      + (~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_4684_nl = nl_MultLoop_acc_4684_nl[17:0];
  assign nl_MultLoop_acc_1146_nl = conv_s2u_18_21(MultLoop_acc_3063_cse_1) + ({(data_rsci_idat[269:252])
      , 3'b001});
  assign MultLoop_acc_1146_nl = nl_MultLoop_acc_1146_nl[20:0];
  assign nl_MultLoop_acc_4448_nl = conv_s2s_12_13(data_rsci_idat[17:6]) + 13'b0000000000001;
  assign MultLoop_acc_4448_nl = nl_MultLoop_acc_4448_nl[12:0];
  assign nl_MultLoop_acc_3389_nl = conv_s2s_18_19(data_rsci_idat[17:0]) + conv_s2s_17_19({(MultLoop_acc_4448_nl)
      , (data_rsci_idat[5:2])});
  assign MultLoop_acc_3389_nl = nl_MultLoop_acc_3389_nl[18:0];
  assign nl_MultLoop_acc_193_nl = conv_s2u_19_22(MultLoop_acc_3389_nl) + ({(~ (data_rsci_idat[17:0]))
      , 4'b0000});
  assign MultLoop_acc_193_nl = nl_MultLoop_acc_193_nl[21:0];
  assign nl_MultLoop_193_MultLoop_acc_3_nl = (readslicef_22_14_8((MultLoop_acc_193_nl)))
      + 14'b00001000111001;
  assign MultLoop_193_MultLoop_acc_3_nl = nl_MultLoop_193_MultLoop_acc_3_nl[13:0];
  assign nl_MultLoop_acc_3469_itm_1  = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4684_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1146_nl))) + conv_s2s_14_16(MultLoop_193_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_3393_nl = ({(data_rsci_idat[827:810]) , 4'b0001}) + conv_s2s_19_22({MultLoop_acc_4133_itm
      , (~ (data_rsci_idat[816:810]))});
  assign MultLoop_acc_3393_nl = nl_MultLoop_acc_3393_nl[21:0];
  assign nl_MultLoop_acc_4451_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_3393_nl)))
      + (~ (data_rsci_idat[827:810]));
  assign MultLoop_acc_4451_nl = nl_MultLoop_acc_4451_nl[17:0];
  assign nl_MultLoop_acc_3394_nl = conv_s2s_20_21({(~ (data_rsci_idat[737:720]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_3394_nl = nl_MultLoop_acc_3394_nl[20:0];
  assign nl_MultLoop_acc_232_nl = conv_s2s_21_22(MultLoop_acc_3394_nl) + ({(data_rsci_idat[737:720])
      , 4'b0100});
  assign MultLoop_acc_232_nl = nl_MultLoop_acc_232_nl[21:0];
  assign nl_MultLoop_acc_3468_itm_1  = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4451_nl)))
      + conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_232_nl)));
  assign nl_MultLoop_acc_4648_nl = conv_s2u_16_19(MultLoop_acc_2040_itm_18_3) + conv_s2u_18_19(data_rsci_idat[755:738]);
  assign MultLoop_acc_4648_nl = nl_MultLoop_acc_4648_nl[18:0];
  assign nl_MultLoop_acc_4452_nl =  -conv_s2s_13_14(data_rsci_idat[701:689]);
  assign MultLoop_acc_4452_nl = nl_MultLoop_acc_4452_nl[13:0];
  assign nl_MultLoop_acc_230_nl = conv_s2s_23_24({(~ (data_rsci_idat[701:684])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[701:684])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4452_nl)
      , (~ (data_rsci_idat[688:684]))});
  assign MultLoop_acc_230_nl = nl_MultLoop_acc_230_nl[23:0];
  assign nl_MultLoop_acc_3399_nl = ({(data_rsci_idat[683:666]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_838_18_4
      , (~ (data_rsci_idat[669:666]))});
  assign MultLoop_acc_3399_nl = nl_MultLoop_acc_3399_nl[19:0];
  assign nl_MultLoop_acc_229_nl = conv_s2s_20_22(MultLoop_acc_3399_nl) + ({(~ (data_rsci_idat[683:666]))
      , 4'b0000});
  assign MultLoop_acc_229_nl = nl_MultLoop_acc_229_nl[21:0];
  assign nl_MultLoop_acc_226_nl = conv_s2u_15_18(data_rsci_idat[629:615]) - (data_rsci_idat[629:612]);
  assign MultLoop_acc_226_nl = nl_MultLoop_acc_226_nl[17:0];
  assign nl_MultLoop_acc_3482_itm_1  = conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4648_nl)))
      + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_230_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_229_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_226_nl)));
  assign nl_MultLoop_acc_3401_nl = (~ (data_rsci_idat[503:486])) + conv_s2s_16_18({Result_acc_190_cse_1
      , (data_rsci_idat[491:489])});
  assign MultLoop_acc_3401_nl = nl_MultLoop_acc_3401_nl[17:0];
  assign nl_MultLoop_acc_1151_nl = conv_s2u_18_22(MultLoop_acc_3401_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[503:486])) , 3'b001});
  assign MultLoop_acc_1151_nl = nl_MultLoop_acc_1151_nl[21:0];
  assign nl_MultLoop_acc_4455_nl = conv_s2s_11_12(data_rsci_idat[449:439]) + 12'b000000000001;
  assign MultLoop_acc_4455_nl = nl_MultLoop_acc_4455_nl[11:0];
  assign nl_MultLoop_acc_3403_nl = conv_s2s_18_19(data_rsci_idat[449:432]) + conv_s2s_15_19({(MultLoop_acc_4455_nl)
      , (data_rsci_idat[438:436])});
  assign MultLoop_acc_3403_nl = nl_MultLoop_acc_3403_nl[18:0];
  assign nl_MultLoop_acc_217_nl = conv_s2u_19_21(MultLoop_acc_3403_nl) + ({(~ (data_rsci_idat[449:432]))
      , 3'b000});
  assign MultLoop_acc_217_nl = nl_MultLoop_acc_217_nl[20:0];
  assign nl_MultLoop_acc_3481_itm_1  = conv_s2s_15_17(MultLoop_acc_1154_itm_21_6[15:1])
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1151_nl))) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_217_nl)))
      + conv_s2s_15_17(data_rsci_idat[467:453]);
  assign nl_MultLoop_acc_3404_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_15_19(data_rsci_idat[413:399]);
  assign MultLoop_acc_3404_nl = nl_MultLoop_acc_3404_nl[18:0];
  assign nl_MultLoop_acc_1150_nl = conv_s2u_19_22(MultLoop_acc_3404_nl) + conv_s2u_21_22({(data_rsci_idat[413:396])
      , 3'b000});
  assign MultLoop_acc_1150_nl = nl_MultLoop_acc_1150_nl[21:0];
  assign nl_MultLoop_acc_4456_nl = conv_s2s_13_14(data_rsci_idat[431:419]) + 14'b00000000000001;
  assign MultLoop_acc_4456_nl = nl_MultLoop_acc_4456_nl[13:0];
  assign nl_MultLoop_acc_3406_nl = conv_s2s_18_19(data_rsci_idat[431:414]) + conv_s2s_17_19({(MultLoop_acc_4456_nl)
      , (data_rsci_idat[418:416])});
  assign MultLoop_acc_3406_nl = nl_MultLoop_acc_3406_nl[18:0];
  assign nl_MultLoop_acc_216_nl = conv_s2u_19_21(MultLoop_acc_3406_nl) + ({(~ (data_rsci_idat[431:414]))
      , 3'b000});
  assign MultLoop_acc_216_nl = nl_MultLoop_acc_216_nl[20:0];
  assign nl_MultLoop_acc_3408_nl = ({(data_rsci_idat[377:360]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_800_18_7
      , (~ (data_rsci_idat[366:360]))});
  assign MultLoop_acc_3408_nl = nl_MultLoop_acc_3408_nl[22:0];
  assign nl_MultLoop_acc_4458_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3408_nl)))
      + (~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_4458_nl = nl_MultLoop_acc_4458_nl[17:0];
  assign nl_MultLoop_acc_4459_nl =  -conv_s2s_13_14(data_rsci_idat[287:275]);
  assign MultLoop_acc_4459_nl = nl_MultLoop_acc_4459_nl[13:0];
  assign nl_MultLoop_acc_208_nl = conv_s2s_19_24({(MultLoop_acc_4459_nl) , (~ (data_rsci_idat[274:270]))})
      + conv_s2s_23_24({(~ (data_rsci_idat[287:270])) , 5'b00001});
  assign MultLoop_acc_208_nl = nl_MultLoop_acc_208_nl[23:0];
  assign nl_MultLoop_acc_3480_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1150_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_216_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4458_nl)))
      + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_208_nl)));
  assign nl_MultLoop_acc_4460_nl =  -conv_s2s_12_13(data_rsci_idat[161:150]);
  assign MultLoop_acc_4460_nl = nl_MultLoop_acc_4460_nl[12:0];
  assign nl_MultLoop_acc_201_nl = conv_s2s_24_25({(~ (data_rsci_idat[161:144])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[161:144])) , 2'b01}) + conv_s2s_19_25({(MultLoop_acc_4460_nl)
      , (~ (data_rsci_idat[149:144]))});
  assign MultLoop_acc_201_nl = nl_MultLoop_acc_201_nl[24:0];
  assign nl_MultLoop_acc_4649_nl = conv_s2u_16_19(MultLoop_acc_2252_itm_20_5) + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_4649_nl = nl_MultLoop_acc_4649_nl[18:0];
  assign nl_MultLoop_acc_3413_nl = conv_s2s_18_19(data_rsci_idat[53:36]) + conv_s2s_16_19(data_rsci_idat[53:38]);
  assign MultLoop_acc_3413_nl = nl_MultLoop_acc_3413_nl[18:0];
  assign nl_MultLoop_acc_1143_nl = conv_s2u_19_22(MultLoop_acc_3413_nl) + conv_s2u_21_22({(data_rsci_idat[53:36])
      , 3'b000});
  assign MultLoop_acc_1143_nl = nl_MultLoop_acc_1143_nl[21:0];
  assign nl_MultLoop_acc_3479_itm_1  = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_201_nl)))
      + conv_s2s_15_17(MultLoop_acc_1145_itm_22_7[15:1]) + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4649_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1143_nl)));
  assign nl_MultLoop_acc_238_nl = conv_s2s_25_26({(~ (data_rsci_idat[845:828])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[845:828])) , 5'b00100}) +
      conv_s2s_20_26({(~ (data_rsci_idat[845:828])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_696_18_7
      , (~ (data_rsci_idat[834:828]))});
  assign MultLoop_acc_238_nl = nl_MultLoop_acc_238_nl[25:0];
  assign nl_MultLoop_acc_3419_nl = ({(data_rsci_idat[773:756]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[773:756])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_688_18_7
      , (~ (data_rsci_idat[762:756]))});
  assign MultLoop_acc_3419_nl = nl_MultLoop_acc_3419_nl[22:0];
  assign nl_MultLoop_acc_4463_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_3419_nl)))
      + (~ (data_rsci_idat[773:756]));
  assign MultLoop_acc_4463_nl = nl_MultLoop_acc_4463_nl[17:0];
  assign nl_MultLoop_acc_3478_itm_1  = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_238_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4463_nl)));
  assign nl_MultLoop_acc_3421_nl = conv_s2s_20_21({(data_rsci_idat[791:774]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[791:774]) + conv_s2s_16_21(data_rsci_idat[791:776]);
  assign MultLoop_acc_3421_nl = nl_MultLoop_acc_3421_nl[20:0];
  assign nl_MultLoop_acc_1157_nl = conv_s2u_21_24(MultLoop_acc_3421_nl) + conv_s2u_23_24({(data_rsci_idat[791:774])
      , 5'b00000});
  assign MultLoop_acc_1157_nl = nl_MultLoop_acc_1157_nl[23:0];
  assign nl_MultLoop_acc_1153_nl = conv_s2u_15_19(data_rsci_idat[593:579]) + conv_s2u_18_19(data_rsci_idat[593:576]);
  assign MultLoop_acc_1153_nl = nl_MultLoop_acc_1153_nl[18:0];
  assign nl_MultLoop_acc_4464_nl = conv_s2s_11_12(data_rsci_idat[521:511]) + 12'b000000000001;
  assign MultLoop_acc_4464_nl = nl_MultLoop_acc_4464_nl[11:0];
  assign nl_MultLoop_acc_3423_nl = conv_s2s_18_19(data_rsci_idat[521:504]) + conv_s2s_15_19({(MultLoop_acc_4464_nl)
      , (data_rsci_idat[510:508])});
  assign MultLoop_acc_3423_nl = nl_MultLoop_acc_3423_nl[18:0];
  assign nl_MultLoop_acc_220_nl = conv_s2u_19_21(MultLoop_acc_3423_nl) + ({(~ (data_rsci_idat[521:504]))
      , 3'b000});
  assign MultLoop_acc_220_nl = nl_MultLoop_acc_220_nl[20:0];
  assign nl_MultLoop_acc_3490_itm_1  = conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1157_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1153_nl))) + conv_s2s_16_18(MultLoop_acc_2390_cse_1[20:5])
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_220_nl)));
  assign nl_MultLoop_acc_4469_nl = conv_s2s_13_14(data_rsci_idat[323:311]) + 14'b00000000000001;
  assign MultLoop_acc_4469_nl = nl_MultLoop_acc_4469_nl[13:0];
  assign nl_MultLoop_acc_3432_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_17_18({(MultLoop_acc_4469_nl)
      , (data_rsci_idat[310:308])});
  assign MultLoop_acc_3432_nl = nl_MultLoop_acc_3432_nl[17:0];
  assign nl_MultLoop_acc_1147_nl = conv_s2u_18_22(MultLoop_acc_3432_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[323:306])) , 3'b001});
  assign MultLoop_acc_1147_nl = nl_MultLoop_acc_1147_nl[21:0];
  assign nl_MultLoop_acc_3434_nl = (~ (data_rsci_idat[233:216])) + conv_s2s_17_18({MultLoop_acc_3974_cse_1
      , (data_rsci_idat[223:218])});
  assign MultLoop_acc_3434_nl = nl_MultLoop_acc_3434_nl[17:0];
  assign nl_MultLoop_acc_3435_nl = ({(data_rsci_idat[233:216]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3434_nl);
  assign MultLoop_acc_3435_nl = nl_MultLoop_acc_3435_nl[19:0];
  assign nl_MultLoop_acc_3436_nl = conv_s2s_22_23({(data_rsci_idat[233:216]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_3435_nl);
  assign MultLoop_acc_3436_nl = nl_MultLoop_acc_3436_nl[22:0];
  assign nl_MultLoop_acc_4471_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3436_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_4471_nl = nl_MultLoop_acc_4471_nl[17:0];
  assign nl_MultLoop_acc_221_nl = conv_s2s_19_25({MultLoop_MultLoop_conc_852_18_6
      , (~ (data_rsci_idat[527:522]))}) + conv_s2s_24_25({(~ (data_rsci_idat[539:522]))
      , 6'b000001});
  assign MultLoop_acc_221_nl = nl_MultLoop_acc_221_nl[24:0];
  assign nl_MultLoop_acc_4466_nl = conv_s2s_11_12(data_rsci_idat[485:475]) + 12'b000000000001;
  assign MultLoop_acc_4466_nl = nl_MultLoop_acc_4466_nl[11:0];
  assign nl_MultLoop_acc_3426_nl = (~ (data_rsci_idat[485:468])) + conv_s2s_16_18({(MultLoop_acc_4466_nl)
      , (data_rsci_idat[474:471])});
  assign MultLoop_acc_3426_nl = nl_MultLoop_acc_3426_nl[17:0];
  assign nl_MultLoop_acc_3427_nl = ({(data_rsci_idat[485:468]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3426_nl);
  assign MultLoop_acc_3427_nl = nl_MultLoop_acc_3427_nl[19:0];
  assign nl_MultLoop_acc_218_nl = conv_s2u_20_22(MultLoop_acc_3427_nl) + ({(~ (data_rsci_idat[485:468]))
      , 4'b0000});
  assign MultLoop_acc_218_nl = nl_MultLoop_acc_218_nl[21:0];
  assign nl_MultLoop_acc_1149_nl = conv_s2u_12_19(data_rsci_idat[395:384]) + conv_s2u_18_19(data_rsci_idat[395:378]);
  assign MultLoop_acc_1149_nl = nl_MultLoop_acc_1149_nl[18:0];
  assign nl_MultLoop_acc_4467_nl =  -conv_s2s_10_11(data_rsci_idat[305:296]);
  assign MultLoop_acc_4467_nl = nl_MultLoop_acc_4467_nl[10:0];
  assign nl_MultLoop_acc_3429_nl = ({(data_rsci_idat[305:288]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4467_nl)
      , (~ (data_rsci_idat[295:288]))});
  assign MultLoop_acc_3429_nl = nl_MultLoop_acc_3429_nl[20:0];
  assign nl_MultLoop_acc_3430_nl = conv_s2s_23_24({(data_rsci_idat[305:288]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_3429_nl);
  assign MultLoop_acc_3430_nl = nl_MultLoop_acc_3430_nl[23:0];
  assign nl_MultLoop_acc_4468_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3430_nl)))
      + (~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_4468_nl = nl_MultLoop_acc_4468_nl[17:0];
  assign nl_MultLoop_acc_4650_nl = conv_s2u_19_20(MultLoop_acc_3213_itm_21_3_1) +
      ({(data_rsci_idat[251:234]) , 2'b01});
  assign MultLoop_acc_4650_nl = nl_MultLoop_acc_4650_nl[19:0];
  assign nl_MultLoop_acc_3438_nl = conv_s2s_21_22({(~ (data_rsci_idat[197:180]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_3438_nl = nl_MultLoop_acc_3438_nl[21:0];
  assign nl_MultLoop_acc_203_nl = conv_s2s_22_23(MultLoop_acc_3438_nl) + ({(data_rsci_idat[197:180])
      , 5'b01000});
  assign MultLoop_acc_203_nl = nl_MultLoop_acc_203_nl[22:0];
  assign nl_MultLoop_acc_3496_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1147_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4471_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_221_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_218_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1149_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4468_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_4650_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_203_nl)));
  assign nl_MultLoop_acc_2063_nl = (~ (data_rsci_idat[215:198])) + conv_s2s_13_18(data_rsci_idat[215:203]);
  assign MultLoop_acc_2063_nl = nl_MultLoop_acc_2063_nl[17:0];
  assign nl_MultLoop_acc_1368_nl = conv_s2u_18_20(MultLoop_acc_2063_nl) + ({(data_rsci_idat[215:198])
      , 2'b01});
  assign MultLoop_acc_1368_nl = nl_MultLoop_acc_1368_nl[19:0];
  assign nl_MultLoop_acc_4040_nl = conv_s2s_11_12(data_rsci_idat[179:169]) + 12'b000000000001;
  assign MultLoop_acc_4040_nl = nl_MultLoop_acc_4040_nl[11:0];
  assign nl_MultLoop_acc_2066_nl = ({(~ (data_rsci_idat[179:162])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[179:162])
      + conv_s2s_17_21({(MultLoop_acc_4040_nl) , (data_rsci_idat[168:164])});
  assign MultLoop_acc_2066_nl = nl_MultLoop_acc_2066_nl[20:0];
  assign nl_MultLoop_acc_1366_nl = conv_s2u_21_24(MultLoop_acc_2066_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[179:162])) , 5'b01000});
  assign MultLoop_acc_1366_nl = nl_MultLoop_acc_1366_nl[23:0];
  assign nl_MultLoop_acc_2056_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_12_18(data_rsci_idat[269:258]);
  assign MultLoop_acc_2056_nl = nl_MultLoop_acc_2056_nl[17:0];
  assign nl_MultLoop_acc_1369_nl = conv_s2u_18_20(MultLoop_acc_2056_nl) + ({(data_rsci_idat[269:252])
      , 2'b01});
  assign MultLoop_acc_1369_nl = nl_MultLoop_acc_1369_nl[19:0];
  assign nl_MultLoop_acc_2058_nl = conv_s2s_21_22({(data_rsci_idat[287:270]) , 3'b000})
      + conv_s2s_19_22(MultLoop_acc_2057_cse_1);
  assign MultLoop_acc_2058_nl = nl_MultLoop_acc_2058_nl[21:0];
  assign nl_MultLoop_acc_1370_nl = conv_s2u_22_24(MultLoop_acc_2058_nl) + conv_s2u_23_24({(data_rsci_idat[287:270])
      , 5'b00000});
  assign MultLoop_acc_1370_nl = nl_MultLoop_acc_1370_nl[23:0];
  assign nl_MultLoop_acc_2060_nl = ({(data_rsci_idat[251:234]) , 6'b000001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_770_18_8
      , (~ (data_rsci_idat[241:234]))});
  assign MultLoop_acc_2060_nl = nl_MultLoop_acc_2060_nl[23:0];
  assign nl_MultLoop_acc_4038_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_2060_nl)))
      + (~ (data_rsci_idat[251:234]));
  assign MultLoop_acc_4038_nl = nl_MultLoop_acc_4038_nl[17:0];
  assign nl_MultLoop_acc_2062_nl = (~ (data_rsci_idat[197:180])) + conv_s2s_16_18({MultLoop_acc_4036_cse_1
      , (data_rsci_idat[186:183])});
  assign MultLoop_acc_2062_nl = nl_MultLoop_acc_2062_nl[17:0];
  assign nl_MultLoop_acc_1367_nl = conv_s2u_18_23(MultLoop_acc_2062_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[197:180])) , 4'b0001});
  assign MultLoop_acc_1367_nl = nl_MultLoop_acc_1367_nl[22:0];
  assign nl_MultLoop_acc_2067_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_15_18(data_rsci_idat[89:75]);
  assign MultLoop_acc_2067_nl = nl_MultLoop_acc_2067_nl[17:0];
  assign nl_MultLoop_acc_1363_nl = conv_s2u_18_21(MultLoop_acc_2067_nl) + ({(data_rsci_idat[89:72])
      , 3'b001});
  assign MultLoop_acc_1363_nl = nl_MultLoop_acc_1363_nl[20:0];
  assign nl_MultLoop_acc_2068_nl = (MultLoop_acc_856_itm_22_7[15:1]) + 15'b111111111110101;
  assign MultLoop_acc_2068_nl = nl_MultLoop_acc_2068_nl[14:0];
  assign nl_MultLoop_acc_855_nl = conv_s2u_14_19(data_rsci_idat[17:4]) + conv_s2u_18_19(data_rsci_idat[17:0]);
  assign MultLoop_acc_855_nl = nl_MultLoop_acc_855_nl[18:0];
  assign nl_MultLoop_866_MultLoop_acc_3_nl = conv_s2s_15_16(MultLoop_acc_2068_nl)
      + (readslicef_19_16_3((MultLoop_acc_855_nl)));
  assign MultLoop_866_MultLoop_acc_3_nl = nl_MultLoop_866_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_2120_itm_1  = conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1368_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1366_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1369_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1370_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4038_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1367_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1363_nl)))
      + conv_s2s_16_18(MultLoop_866_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_4607_nl = conv_s2u_13_19(MultLoop_acc_2073_cse_1[18:6])
      + conv_s2u_18_19(data_rsci_idat[665:648]);
  assign MultLoop_acc_4607_nl = nl_MultLoop_acc_4607_nl[18:0];
  assign nl_MultLoop_acc_2074_nl = ({(data_rsci_idat[593:576]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[593:576]));
  assign MultLoop_acc_2074_nl = nl_MultLoop_acc_2074_nl[20:0];
  assign nl_MultLoop_acc_2075_nl = conv_s2s_24_25({(data_rsci_idat[593:576]) , 6'b000000})
      + conv_s2s_21_25(MultLoop_acc_2074_nl);
  assign MultLoop_acc_2075_nl = nl_MultLoop_acc_2075_nl[24:0];
  assign nl_MultLoop_acc_4044_nl = conv_s2u_17_19(readslicef_25_17_8((MultLoop_acc_2075_nl)))
      + conv_s2u_18_19(data_rsci_idat[593:576]);
  assign MultLoop_acc_4044_nl = nl_MultLoop_acc_4044_nl[18:0];
  assign nl_MultLoop_acc_2070_nl = ({(data_rsci_idat[53:36]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_802_18_8
      , (~ (data_rsci_idat[43:36]))});
  assign MultLoop_acc_2070_nl = nl_MultLoop_acc_2070_nl[20:0];
  assign nl_MultLoop_acc_4042_nl = conv_s2u_13_18(readslicef_21_13_8((MultLoop_acc_2070_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_4042_nl = nl_MultLoop_acc_4042_nl[17:0];
  assign nl_MultLoop_acc_1362_nl = conv_s2u_18_24(MultLoop_acc_1636_cse_1) + conv_s2u_23_24({(~
      (data_rsci_idat[71:54])) , 5'b00001});
  assign MultLoop_acc_1362_nl = nl_MultLoop_acc_1362_nl[23:0];
  assign nl_MultLoop_acc_2119_itm_1  = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4607_nl)))
      + conv_s2s_17_18(MultLoop_acc_1993_itm_18_2) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4044_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4042_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1362_nl)));
  assign nl_MultLoop_acc_2076_nl = ({(data_rsci_idat[611:594]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[611:594]));
  assign MultLoop_acc_2076_nl = nl_MultLoop_acc_2076_nl[19:0];
  assign nl_MultLoop_acc_2077_nl = conv_s2s_24_25({(data_rsci_idat[611:594]) , 6'b000000})
      + conv_s2s_20_25(MultLoop_acc_2076_nl);
  assign MultLoop_acc_2077_nl = nl_MultLoop_acc_2077_nl[24:0];
  assign nl_MultLoop_acc_4045_nl = conv_s2u_17_19(readslicef_25_17_8((MultLoop_acc_2077_nl)))
      + conv_s2u_18_19(data_rsci_idat[611:594]);
  assign MultLoop_acc_4045_nl = nl_MultLoop_acc_4045_nl[18:0];
  assign nl_MultLoop_acc_2078_nl = ({(data_rsci_idat[395:378]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[395:378]));
  assign MultLoop_acc_2078_nl = nl_MultLoop_acc_2078_nl[21:0];
  assign nl_MultLoop_acc_874_nl = conv_s2s_22_25(MultLoop_acc_2078_nl) + conv_s2s_24_25({(data_rsci_idat[395:378])
      , 6'b000000});
  assign MultLoop_acc_874_nl = nl_MultLoop_acc_874_nl[24:0];
  assign nl_MultLoop_acc_2080_nl = ({(data_rsci_idat[125:108]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2079_cse_1);
  assign MultLoop_acc_2080_nl = nl_MultLoop_acc_2080_nl[19:0];
  assign nl_MultLoop_acc_1365_nl = conv_s2u_20_23(MultLoop_acc_2080_nl) + conv_s2u_22_23({(data_rsci_idat[125:108])
      , 4'b0000});
  assign MultLoop_acc_1365_nl = nl_MultLoop_acc_1365_nl[22:0];
  assign nl_MultLoop_acc_4608_nl = conv_s2u_14_19(Result_acc_111_cse_1[18:5]) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_4608_nl = nl_MultLoop_acc_4608_nl[18:0];
  assign nl_MultLoop_acc_2118_itm_1  = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4045_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_874_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1365_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4608_nl)));
  assign nl_MultLoop_acc_4046_nl =  -conv_s2s_15_16(data_rsci_idat[719:705]);
  assign MultLoop_acc_4046_nl = nl_MultLoop_acc_4046_nl[15:0];
  assign nl_MultLoop_acc_892_nl = conv_s2s_19_22({(MultLoop_acc_4046_nl) , (~ (data_rsci_idat[704:702]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[719:702])) , 3'b001});
  assign MultLoop_acc_892_nl = nl_MultLoop_acc_892_nl[21:0];
  assign nl_MultLoop_acc_4667_nl = conv_s2u_19_20(Result_acc_102_itm_20_2_1) + ({(data_rsci_idat[521:504])
      , 2'b01});
  assign MultLoop_acc_4667_nl = nl_MultLoop_acc_4667_nl[19:0];
  assign nl_MultLoop_acc_2012_nl = ({(data_rsci_idat[539:522]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_852_18_6
      , (~ (data_rsci_idat[527:522]))});
  assign MultLoop_acc_2012_nl = nl_MultLoop_acc_2012_nl[21:0];
  assign nl_MultLoop_acc_4048_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2012_nl)))
      + (~ (data_rsci_idat[539:522]));
  assign MultLoop_acc_4048_nl = nl_MultLoop_acc_4048_nl[17:0];
  assign nl_MultLoop_acc_2014_nl = conv_s2s_18_19(data_rsci_idat[449:432]) + conv_s2s_16_19({MultLoop_MultLoop_conc_768_15_2
      , (data_rsci_idat[436:435])});
  assign MultLoop_acc_2014_nl = nl_MultLoop_acc_2014_nl[18:0];
  assign nl_MultLoop_acc_877_nl = conv_s2u_19_20(MultLoop_acc_2014_nl) + ({(~ (data_rsci_idat[449:432]))
      , 2'b00});
  assign MultLoop_acc_877_nl = nl_MultLoop_acc_877_nl[19:0];
  assign nl_MultLoop_acc_2091_itm_1  = conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_892_nl)))
      + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_4667_nl))) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4048_nl)))
      + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_877_nl)));
  assign nl_MultLoop_acc_4609_nl = conv_s2u_19_20(MultLoop_acc_1512_itm_20_2_1) +
      ({(data_rsci_idat[845:828]) , 2'b01});
  assign MultLoop_acc_4609_nl = nl_MultLoop_acc_4609_nl[19:0];
  assign nl_MultLoop_acc_4050_nl =  -conv_s2s_14_15(data_rsci_idat[647:634]);
  assign MultLoop_acc_4050_nl = nl_MultLoop_acc_4050_nl[14:0];
  assign nl_MultLoop_acc_888_nl = conv_s2s_19_23({(MultLoop_acc_4050_nl) , (~ (data_rsci_idat[633:630]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[647:630])) , 4'b0001});
  assign MultLoop_acc_888_nl = nl_MultLoop_acc_888_nl[22:0];
  assign nl_MultLoop_acc_2082_nl = (readslicef_23_13_10((MultLoop_acc_888_nl))) +
      conv_s2s_9_13(data_rsci_idat[143:135]);
  assign MultLoop_acc_2082_nl = nl_MultLoop_acc_2082_nl[12:0];
  assign nl_MultLoop_acc_2090_itm_1  = conv_s2s_15_16(readslicef_20_15_5((MultLoop_acc_4609_nl)))
      + conv_s2s_14_16(MultLoop_acc_119_itm_23_9[14:1]) + conv_s2s_13_16(MultLoop_acc_2082_nl);
  assign nl_MultLoop_acc_2016_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_13_18(data_rsci_idat[557:545]);
  assign MultLoop_acc_2016_nl = nl_MultLoop_acc_2016_nl[17:0];
  assign nl_MultLoop_acc_1374_nl = conv_s2u_18_20(MultLoop_acc_2016_nl) + ({(data_rsci_idat[557:540])
      , 2'b01});
  assign MultLoop_acc_1374_nl = nl_MultLoop_acc_1374_nl[19:0];
  assign nl_MultLoop_acc_4610_nl = conv_s2u_16_19(MultLoop_acc_1727_cse_1[18:3])
      + conv_s2u_18_19(data_rsci_idat[575:558]);
  assign MultLoop_acc_4610_nl = nl_MultLoop_acc_4610_nl[18:0];
  assign nl_MultLoop_acc_2018_nl = (~ (data_rsci_idat[485:468])) + conv_s2s_15_18(data_rsci_idat[485:471]);
  assign MultLoop_acc_2018_nl = nl_MultLoop_acc_2018_nl[17:0];
  assign nl_MultLoop_acc_2019_nl = conv_s2s_20_21({(~ (data_rsci_idat[485:468]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2018_nl);
  assign MultLoop_acc_2019_nl = nl_MultLoop_acc_2019_nl[20:0];
  assign nl_MultLoop_acc_1373_nl = conv_s2u_21_22(MultLoop_acc_2019_nl) + ({(data_rsci_idat[485:468])
      , 4'b0100});
  assign MultLoop_acc_1373_nl = nl_MultLoop_acc_1373_nl[21:0];
  assign nl_MultLoop_acc_2105_itm_1  = conv_s2s_15_17(MultLoop_acc_4592_itm_18_3[15:1])
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1374_nl))) + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4610_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1373_nl)));
  assign nl_MultLoop_acc_4051_nl = conv_s2s_12_13(data_rsci_idat[359:348]) + 13'b0000000000001;
  assign MultLoop_acc_4051_nl = nl_MultLoop_acc_4051_nl[12:0];
  assign nl_MultLoop_acc_2021_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_17_18({(MultLoop_acc_4051_nl)
      , (data_rsci_idat[347:344])});
  assign MultLoop_acc_2021_nl = nl_MultLoop_acc_2021_nl[17:0];
  assign nl_MultLoop_acc_1371_nl = conv_s2u_18_23(MultLoop_acc_2021_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[359:342])) , 4'b0001});
  assign MultLoop_acc_1371_nl = nl_MultLoop_acc_1371_nl[22:0];
  assign nl_MultLoop_acc_2023_nl = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_734_18_7
      , (~ (data_rsci_idat[294:288]))});
  assign MultLoop_acc_2023_nl = nl_MultLoop_acc_2023_nl[19:0];
  assign nl_MultLoop_acc_2024_nl = conv_s2s_23_24({(data_rsci_idat[305:288]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_2023_nl);
  assign MultLoop_acc_2024_nl = nl_MultLoop_acc_2024_nl[23:0];
  assign nl_MultLoop_acc_4053_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_2024_nl)))
      + (~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_4053_nl = nl_MultLoop_acc_4053_nl[17:0];
  assign nl_MultLoop_acc_4611_nl = conv_s2u_16_19(MultLoop_acc_2026_itm_21_6) + conv_s2u_18_19(data_rsci_idat[233:216]);
  assign MultLoop_acc_4611_nl = nl_MultLoop_acc_4611_nl[18:0];
  assign nl_MultLoop_acc_2104_itm_1  = conv_s2s_15_17(MultLoop_acc_408_itm_23_9)
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1371_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4053_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4611_nl)));
  assign nl_MultLoop_acc_2028_nl = ({(data_rsci_idat[863:846]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_720_18_7
      , (~ (data_rsci_idat[852:846]))});
  assign MultLoop_acc_2028_nl = nl_MultLoop_acc_2028_nl[22:0];
  assign nl_MultLoop_acc_4055_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_2028_nl)))
      + (~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_4055_nl = nl_MultLoop_acc_4055_nl[17:0];
  assign nl_MultLoop_acc_897_nl = conv_s2s_24_25({(~ (data_rsci_idat[809:792])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[809:792])) , 4'b0100}) + conv_s2s_21_25(MultLoop_acc_2030_cse_1);
  assign MultLoop_acc_897_nl = nl_MultLoop_acc_897_nl[24:0];
  assign nl_MultLoop_acc_2103_itm_1  = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4055_nl)))
      + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_897_nl)));
  assign nl_MultLoop_acc_2032_nl = (~ (data_rsci_idat[827:810])) + conv_s2s_13_18(data_rsci_idat[827:815]);
  assign MultLoop_acc_2032_nl = nl_MultLoop_acc_2032_nl[17:0];
  assign nl_MultLoop_acc_1383_nl = conv_s2u_18_21(MultLoop_acc_2032_nl) + ({(data_rsci_idat[827:810])
      , 3'b001});
  assign MultLoop_acc_1383_nl = nl_MultLoop_acc_1383_nl[20:0];
  assign nl_MultLoop_acc_4612_nl = conv_s2u_18_19(data_rsci_idat[773:756]) + conv_s2u_16_19(MultLoop_acc_1723_cse_1[19:4]);
  assign MultLoop_acc_4612_nl = nl_MultLoop_acc_4612_nl[18:0];
  assign nl_MultLoop_acc_4057_nl = conv_s2u_16_19(readslicef_19_16_3((MultLoop_acc_4612_nl)))
      + conv_s2u_18_19(data_rsci_idat[773:756]);
  assign MultLoop_acc_4057_nl = nl_MultLoop_acc_4057_nl[18:0];
  assign nl_MultLoop_acc_2036_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2035_cse_1);
  assign MultLoop_acc_2036_nl = nl_MultLoop_acc_2036_nl[19:0];
  assign nl_MultLoop_acc_2037_nl = ({(~ (data_rsci_idat[791:774])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2036_nl);
  assign MultLoop_acc_2037_nl = nl_MultLoop_acc_2037_nl[21:0];
  assign nl_MultLoop_acc_1382_nl = conv_s2u_22_24(MultLoop_acc_2037_nl) + ({(data_rsci_idat[791:774])
      , 6'b010000});
  assign MultLoop_acc_1382_nl = nl_MultLoop_acc_1382_nl[23:0];
  assign nl_MultLoop_acc_2039_nl = (~ (data_rsci_idat[737:720])) + conv_s2s_16_18({MultLoop_MultLoop_conc_714_15_2
      , (data_rsci_idat[724:723])});
  assign MultLoop_acc_2039_nl = nl_MultLoop_acc_2039_nl[17:0];
  assign nl_MultLoop_acc_1380_nl = conv_s2u_18_21(MultLoop_acc_2039_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[737:720])) , 2'b01});
  assign MultLoop_acc_1380_nl = nl_MultLoop_acc_1380_nl[20:0];
  assign nl_MultLoop_acc_2115_itm_1  = conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1383_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4057_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1382_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1380_nl)));
  assign nl_MultLoop_acc_2046_nl = ({(~ (data_rsci_idat[413:396])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[413:396])
      + conv_s2s_16_20(data_rsci_idat[413:398]);
  assign MultLoop_acc_2046_nl = nl_MultLoop_acc_2046_nl[19:0];
  assign nl_MultLoop_acc_2047_nl = conv_s2s_22_23({(~ (data_rsci_idat[413:396]))
      , 4'b0100}) + conv_s2s_20_23(MultLoop_acc_2046_nl);
  assign MultLoop_acc_2047_nl = nl_MultLoop_acc_2047_nl[22:0];
  assign nl_MultLoop_acc_1372_nl = conv_s2u_23_24(MultLoop_acc_2047_nl) + ({(data_rsci_idat[413:396])
      , 6'b010000});
  assign MultLoop_acc_1372_nl = nl_MultLoop_acc_1372_nl[23:0];
  assign nl_MultLoop_acc_2050_nl = ({(data_rsci_idat[377:360]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[377:360])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_800_18_7
      , (~ (data_rsci_idat[366:360]))});
  assign MultLoop_acc_2050_nl = nl_MultLoop_acc_2050_nl[22:0];
  assign nl_MultLoop_acc_4062_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_2050_nl)))
      + (~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_4062_nl = nl_MultLoop_acc_4062_nl[17:0];
  assign nl_MultLoop_acc_4613_nl = conv_s2u_15_19(MultLoop_acc_2040_itm_18_3[15:1])
      + conv_s2u_18_19(data_rsci_idat[755:738]);
  assign MultLoop_acc_4613_nl = nl_MultLoop_acc_4613_nl[18:0];
  assign nl_MultLoop_acc_4059_nl = conv_s2s_12_13(data_rsci_idat[629:618]) + 13'b0000000000001;
  assign MultLoop_acc_4059_nl = nl_MultLoop_acc_4059_nl[12:0];
  assign nl_MultLoop_acc_2042_nl = (~ (data_rsci_idat[629:612])) + conv_s2s_17_18({(MultLoop_acc_4059_nl)
      , (data_rsci_idat[617:614])});
  assign MultLoop_acc_2042_nl = nl_MultLoop_acc_2042_nl[17:0];
  assign nl_MultLoop_acc_1376_nl = conv_s2u_18_23(MultLoop_acc_2042_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[629:612])) , 4'b0001});
  assign MultLoop_acc_1376_nl = nl_MultLoop_acc_1376_nl[22:0];
  assign nl_MultLoop_acc_2044_nl = conv_s2s_18_19(data_rsci_idat[467:450]) + conv_s2s_14_19({MultLoop_acc_4030_cse_1
      , (data_rsci_idat[457:455])});
  assign MultLoop_acc_2044_nl = nl_MultLoop_acc_2044_nl[18:0];
  assign nl_MultLoop_acc_878_nl = conv_s2u_19_21(MultLoop_acc_2044_nl) + ({(~ (data_rsci_idat[467:450]))
      , 3'b000});
  assign MultLoop_acc_878_nl = nl_MultLoop_acc_878_nl[20:0];
  assign nl_MultLoop_acc_4063_nl =  -conv_s2s_11_12(data_rsci_idat[341:331]);
  assign MultLoop_acc_4063_nl = nl_MultLoop_acc_4063_nl[11:0];
  assign nl_MultLoop_acc_2052_nl = ({(data_rsci_idat[341:324]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4063_nl)
      , (~ (data_rsci_idat[330:324]))});
  assign MultLoop_acc_2052_nl = nl_MultLoop_acc_2052_nl[20:0];
  assign nl_MultLoop_acc_2053_nl = ({(~ (data_rsci_idat[341:324])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_2052_nl);
  assign MultLoop_acc_2053_nl = nl_MultLoop_acc_2053_nl[22:0];
  assign nl_MultLoop_acc_871_nl = conv_s2s_23_26(MultLoop_acc_2053_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[341:324])) , 7'b0100000});
  assign MultLoop_acc_871_nl = nl_MultLoop_acc_871_nl[25:0];
  assign nl_MultLoop_acc_2055_nl = conv_s2s_24_25({(~ (data_rsci_idat[323:306]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[323:306])) , 4'b0001}) +
      conv_s2s_18_25(~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_2055_nl = nl_MultLoop_acc_2055_nl[24:0];
  assign nl_MultLoop_acc_870_nl = conv_s2s_25_26(MultLoop_acc_2055_nl) + ({(data_rsci_idat[323:306])
      , 8'b01000000});
  assign MultLoop_acc_870_nl = nl_MultLoop_acc_870_nl[25:0];
  assign nl_MultLoop_acc_2121_itm_1  = conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1372_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4062_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4613_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1376_nl))) + conv_s2s_16_18(data_rsci_idat[161:146])
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_878_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_871_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_870_nl)));
  assign nl_MultLoop_acc_4415_nl = conv_s2s_13_14(data_rsci_idat[467:455]) + 14'b00000000000001;
  assign MultLoop_acc_4415_nl = nl_MultLoop_acc_4415_nl[13:0];
  assign nl_MultLoop_acc_3328_nl = (~ (data_rsci_idat[467:450])) + conv_s2s_17_18({(MultLoop_acc_4415_nl)
      , (data_rsci_idat[454:452])});
  assign MultLoop_acc_3328_nl = nl_MultLoop_acc_3328_nl[17:0];
  assign nl_MultLoop_acc_1167_nl = conv_s2u_18_22(MultLoop_acc_3328_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[467:450])) , 3'b001});
  assign MultLoop_acc_1167_nl = nl_MultLoop_acc_1167_nl[21:0];
  assign nl_MultLoop_acc_3329_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_14_19(data_rsci_idat[413:400]);
  assign MultLoop_acc_3329_nl = nl_MultLoop_acc_3329_nl[18:0];
  assign nl_MultLoop_acc_1166_nl = conv_s2u_19_21(MultLoop_acc_3329_nl) + conv_s2u_20_21({(data_rsci_idat[413:396])
      , 2'b00});
  assign MultLoop_acc_1166_nl = nl_MultLoop_acc_1166_nl[20:0];
  assign nl_MultLoop_acc_256_nl = conv_s2s_25_26({(~ (data_rsci_idat[305:288])) ,
      7'b0000100}) + conv_s2s_20_26({(~ (data_rsci_idat[305:288])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_734_18_7
      , (~ (data_rsci_idat[294:288]))});
  assign MultLoop_acc_256_nl = nl_MultLoop_acc_256_nl[25:0];
  assign nl_MultLoop_acc_4417_nl =  -conv_s2s_10_11(data_rsci_idat[269:260]);
  assign MultLoop_acc_4417_nl = nl_MultLoop_acc_4417_nl[10:0];
  assign nl_MultLoop_acc_254_nl = conv_s2s_26_27({(~ (data_rsci_idat[269:252])) ,
      8'b00010000}) + conv_s2s_22_27({(~ (data_rsci_idat[269:252])) , 4'b0100}) +
      conv_s2s_20_27({(~ (data_rsci_idat[269:252])) , 2'b01}) + conv_s2s_19_27({(MultLoop_acc_4417_nl)
      , (~ (data_rsci_idat[259:252]))});
  assign MultLoop_acc_254_nl = nl_MultLoop_acc_254_nl[26:0];
  assign nl_MultLoop_acc_3378_itm_1  = conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1167_nl)))
      + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1166_nl))) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_256_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_254_nl)));
  assign nl_MultLoop_acc_243_nl = conv_s2u_13_18(data_rsci_idat[71:59]) - (data_rsci_idat[71:54]);
  assign MultLoop_acc_243_nl = nl_MultLoop_acc_243_nl[17:0];
  assign nl_MultLoop_acc_240_nl = conv_s2u_15_18(data_rsci_idat[17:3]) - (data_rsci_idat[17:0]);
  assign MultLoop_acc_240_nl = nl_MultLoop_acc_240_nl[17:0];
  assign nl_MultLoop_241_MultLoop_acc_3_nl = (readslicef_18_13_5((MultLoop_acc_240_nl)))
      + 13'b0000010101001;
  assign MultLoop_241_MultLoop_acc_3_nl = nl_MultLoop_241_MultLoop_acc_3_nl[12:0];
  assign nl_MultLoop_acc_242_nl = conv_s2u_15_18(data_rsci_idat[53:39]) - (data_rsci_idat[53:36]);
  assign MultLoop_acc_242_nl = nl_MultLoop_acc_242_nl[17:0];
  assign nl_MultLoop_acc_3341_nl = conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_243_nl)))
      + conv_s2s_13_15(MultLoop_241_MultLoop_acc_3_nl) + conv_s2s_11_15(readslicef_18_11_7((MultLoop_acc_242_nl)));
  assign MultLoop_acc_3341_nl = nl_MultLoop_acc_3341_nl[14:0];
  assign nl_MultLoop_acc_4645_nl = ({(data_rsci_idat[35:18]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_3338_itm_20_2_1);
  assign MultLoop_acc_4645_nl = nl_MultLoop_acc_4645_nl[19:0];
  assign nl_MultLoop_acc_4419_nl = conv_s2u_15_19(readslicef_20_15_5((MultLoop_acc_4645_nl)))
      + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_4419_nl = nl_MultLoop_acc_4419_nl[18:0];
  assign nl_MultLoop_244_MultLoop_acc_3_nl = conv_s2s_15_16(MultLoop_acc_3341_nl)
      + (readslicef_19_16_3((MultLoop_acc_4419_nl)));
  assign MultLoop_244_MultLoop_acc_3_nl = nl_MultLoop_244_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_3342_nl = conv_s2s_18_19(data_rsci_idat[89:72]) + conv_s2s_16_19(data_rsci_idat[89:74]);
  assign MultLoop_acc_3342_nl = nl_MultLoop_acc_3342_nl[18:0];
  assign nl_MultLoop_acc_1159_nl = conv_s2u_19_22(MultLoop_acc_3342_nl) + conv_s2u_21_22({(data_rsci_idat[89:72])
      , 3'b000});
  assign MultLoop_acc_1159_nl = nl_MultLoop_acc_1159_nl[21:0];
  assign nl_MultLoop_acc_247_nl = conv_s2s_24_25({(~ (data_rsci_idat[143:126])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[143:126])) , 4'b0001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_824_18_6
      , (~ (data_rsci_idat[131:126]))});
  assign MultLoop_acc_247_nl = nl_MultLoop_acc_247_nl[24:0];
  assign nl_MultLoop_acc_3343_nl = (MultLoop_acc_1848_itm_21_6[15:3]) + conv_s2s_12_13(Result_acc_111_cse_1[18:7]);
  assign MultLoop_acc_3343_nl = nl_MultLoop_acc_3343_nl[12:0];
  assign nl_MultLoop_acc_3344_nl = (readslicef_25_15_10((MultLoop_acc_247_nl))) +
      conv_s2s_13_15(MultLoop_acc_3343_nl);
  assign MultLoop_acc_3344_nl = nl_MultLoop_acc_3344_nl[14:0];
  assign nl_MultLoop_248_MultLoop_acc_3_nl = conv_s2s_16_17(MultLoop_244_MultLoop_acc_3_nl)
      + conv_s2s_16_17(readslicef_22_16_6((MultLoop_acc_1159_nl))) + conv_s2s_15_17(MultLoop_acc_3344_nl);
  assign MultLoop_248_MultLoop_acc_3_nl = nl_MultLoop_248_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_4420_nl =  -conv_s2s_16_17(data_rsci_idat[557:542]);
  assign MultLoop_acc_4420_nl = nl_MultLoop_acc_4420_nl[16:0];
  assign nl_MultLoop_acc_269_nl = conv_s2s_19_21({(MultLoop_acc_4420_nl) , (~ (data_rsci_idat[541:540]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[557:540])) , 2'b01});
  assign MultLoop_acc_269_nl = nl_MultLoop_acc_269_nl[20:0];
  assign nl_MultLoop_acc_4421_nl =  -conv_s2s_15_16(data_rsci_idat[197:183]);
  assign MultLoop_acc_4421_nl = nl_MultLoop_acc_4421_nl[15:0];
  assign nl_MultLoop_acc_250_nl = conv_s2s_19_22({(MultLoop_acc_4421_nl) , (~ (data_rsci_idat[182:180]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[197:180])) , 3'b001});
  assign MultLoop_acc_250_nl = nl_MultLoop_acc_250_nl[21:0];
  assign nl_MultLoop_acc_3346_nl = (readslicef_22_13_9((MultLoop_acc_250_nl))) +
      conv_s2s_9_13(data_rsci_idat[449:441]);
  assign MultLoop_acc_3346_nl = nl_MultLoop_acc_3346_nl[12:0];
  assign nl_MultLoop_acc_3348_nl = (readslicef_21_14_7((MultLoop_acc_269_nl))) +
      conv_s2s_13_14(MultLoop_acc_3346_nl);
  assign MultLoop_acc_3348_nl = nl_MultLoop_acc_3348_nl[13:0];
  assign nl_MultLoop_acc_3267_nl = conv_s2s_20_21({(~ (data_rsci_idat[791:774]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[791:774]));
  assign MultLoop_acc_3267_nl = nl_MultLoop_acc_3267_nl[20:0];
  assign nl_MultLoop_acc_282_nl = conv_s2s_21_22(MultLoop_acc_3267_nl) + ({(data_rsci_idat[791:774])
      , 4'b0100});
  assign MultLoop_acc_282_nl = nl_MultLoop_acc_282_nl[21:0];
  assign nl_MultLoop_acc_1163_nl = conv_s2u_18_21(MultLoop_acc_2574_cse_1) + ({(data_rsci_idat[341:324])
      , 3'b001});
  assign MultLoop_acc_1163_nl = nl_MultLoop_acc_1163_nl[20:0];
  assign nl_MultLoop_acc_3271_nl = conv_s2s_18_19(data_rsci_idat[593:576]) + conv_s2s_17_19({MultLoop_MultLoop_conc_772_16_2
      , (data_rsci_idat[579:578])});
  assign MultLoop_acc_3271_nl = nl_MultLoop_acc_3271_nl[18:0];
  assign nl_MultLoop_acc_271_nl = conv_s2u_19_20(MultLoop_acc_3271_nl) + ({(~ (data_rsci_idat[593:576]))
      , 2'b00});
  assign MultLoop_acc_271_nl = nl_MultLoop_acc_271_nl[19:0];
  assign nl_MultLoop_acc_3368_itm_1  = conv_s2s_17_18(MultLoop_248_MultLoop_acc_3_nl)
      + conv_s2s_14_18(MultLoop_acc_3348_nl) + conv_s2s_13_18(readslicef_22_13_9((MultLoop_acc_282_nl)))
      + conv_s2s_13_18(readslicef_21_13_8((MultLoop_acc_1163_nl))) + conv_s2s_14_18(MultLoop_acc_1541_itm_18_2[16:3])
      + conv_s2s_14_18(readslicef_20_14_6((MultLoop_acc_271_nl)));
  assign nl_MultLoop_acc_3274_nl = conv_s2s_20_21({(~ (data_rsci_idat[845:828]))
      , 2'b01}) + conv_s2s_18_21(Result_acc_143_cse_1);
  assign MultLoop_acc_3274_nl = nl_MultLoop_acc_3274_nl[20:0];
  assign nl_MultLoop_acc_1174_nl = conv_s2u_21_22(MultLoop_acc_3274_nl) + ({(data_rsci_idat[845:828])
      , 4'b0100});
  assign MultLoop_acc_1174_nl = nl_MultLoop_acc_1174_nl[21:0];
  assign nl_MultLoop_acc_3275_nl = (~ (data_rsci_idat[809:792])) + conv_s2s_14_18(data_rsci_idat[809:796]);
  assign MultLoop_acc_3275_nl = nl_MultLoop_acc_3275_nl[17:0];
  assign nl_MultLoop_acc_1173_nl = conv_s2u_18_20(MultLoop_acc_3275_nl) + ({(data_rsci_idat[809:792])
      , 2'b01});
  assign MultLoop_acc_1173_nl = nl_MultLoop_acc_1173_nl[19:0];
  assign nl_MultLoop_acc_3277_nl = conv_s2s_20_21({(data_rsci_idat[719:702]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_2566_cse_1);
  assign MultLoop_acc_3277_nl = nl_MultLoop_acc_3277_nl[20:0];
  assign nl_MultLoop_acc_1172_nl = conv_s2u_21_23(MultLoop_acc_3277_nl) + conv_s2u_22_23({(data_rsci_idat[719:702])
      , 4'b0000});
  assign MultLoop_acc_1172_nl = nl_MultLoop_acc_1172_nl[22:0];
  assign nl_MultLoop_acc_3279_nl = ({(~ (data_rsci_idat[665:648])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_1743_cse_1);
  assign MultLoop_acc_3279_nl = nl_MultLoop_acc_3279_nl[22:0];
  assign nl_MultLoop_acc_275_nl = conv_s2s_23_25(MultLoop_acc_3279_nl) + ({(data_rsci_idat[665:648])
      , 7'b0100000});
  assign MultLoop_acc_275_nl = nl_MultLoop_acc_275_nl[24:0];
  assign nl_MultLoop_acc_3367_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1174_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1173_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1172_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_275_nl)));
  assign nl_MultLoop_acc_4646_nl = conv_s2u_19_21(MultLoop_acc_2385_cse_1[20:2])
      + ({(data_rsci_idat[683:666]) , 3'b001});
  assign MultLoop_acc_4646_nl = nl_MultLoop_acc_4646_nl[20:0];
  assign nl_MultLoop_acc_4647_nl = conv_s2u_15_19(MultLoop_acc_3281_itm_20_6) + conv_s2u_18_19(data_rsci_idat[647:630]);
  assign MultLoop_acc_4647_nl = nl_MultLoop_acc_4647_nl[18:0];
  assign nl_MultLoop_acc_3282_nl = conv_s2s_20_21({(~ (data_rsci_idat[575:558]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[575:558]));
  assign MultLoop_acc_3282_nl = nl_MultLoop_acc_3282_nl[20:0];
  assign nl_MultLoop_acc_270_nl = conv_s2s_21_22(MultLoop_acc_3282_nl) + ({(data_rsci_idat[575:558])
      , 4'b0100});
  assign MultLoop_acc_270_nl = nl_MultLoop_acc_270_nl[21:0];
  assign nl_MultLoop_acc_3284_nl = conv_s2s_20_21({(data_rsci_idat[503:486]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_3283_cse);
  assign MultLoop_acc_3284_nl = nl_MultLoop_acc_3284_nl[20:0];
  assign nl_MultLoop_acc_1169_nl = conv_s2u_21_23(MultLoop_acc_3284_nl) + conv_s2u_22_23({(data_rsci_idat[503:486])
      , 4'b0000});
  assign MultLoop_acc_1169_nl = nl_MultLoop_acc_1169_nl[22:0];
  assign nl_MultLoop_acc_3366_itm_1  = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_4646_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4647_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_270_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1169_nl)));
  assign nl_MultLoop_acc_3289_nl = ({(~ (data_rsci_idat[863:846])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[863:846])
      + conv_s2s_17_20({MultLoop_acc_4011_cse_1 , (data_rsci_idat[853:848])});
  assign MultLoop_acc_3289_nl = nl_MultLoop_acc_3289_nl[19:0];
  assign nl_MultLoop_acc_3290_nl = ({(data_rsci_idat[863:846]) , 4'b0100}) + conv_s2s_20_22(MultLoop_acc_3289_nl);
  assign MultLoop_acc_3290_nl = nl_MultLoop_acc_3290_nl[21:0];
  assign nl_MultLoop_acc_4424_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3290_nl)))
      + (~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_4424_nl = nl_MultLoop_acc_4424_nl[17:0];
  assign nl_MultLoop_acc_1164_nl = conv_s2u_15_19(data_rsci_idat[377:363]) + conv_s2u_18_19(data_rsci_idat[377:360]);
  assign MultLoop_acc_1164_nl = nl_MultLoop_acc_1164_nl[18:0];
  assign nl_MultLoop_acc_3286_nl = conv_s2s_22_23({(~ (data_rsci_idat[179:162]))
      , 4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_18_23(~
      (data_rsci_idat[179:162]));
  assign MultLoop_acc_3286_nl = nl_MultLoop_acc_3286_nl[22:0];
  assign nl_MultLoop_acc_249_nl = conv_s2s_23_24(MultLoop_acc_3286_nl) + ({(data_rsci_idat[179:162])
      , 6'b010000});
  assign MultLoop_acc_249_nl = nl_MultLoop_acc_249_nl[23:0];
  assign nl_MultLoop_acc_3365_itm_1  = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4424_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_1164_nl))) + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_249_nl)));
  assign nl_MultLoop_acc_284_nl = conv_s2s_25_26({(~ (data_rsci_idat[827:810])) ,
      7'b0010000}) + conv_s2s_22_26({(~ (data_rsci_idat[827:810])) , 4'b0001}) +
      conv_s2s_19_26({MultLoop_acc_4133_itm , (~ (data_rsci_idat[816:810]))});
  assign MultLoop_acc_284_nl = nl_MultLoop_acc_284_nl[25:0];
  assign nl_MultLoop_acc_3293_nl = conv_s2s_21_22({(~ (data_rsci_idat[773:756]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[773:756]));
  assign MultLoop_acc_3293_nl = nl_MultLoop_acc_3293_nl[21:0];
  assign nl_MultLoop_acc_281_nl = conv_s2s_22_24(MultLoop_acc_3293_nl) + ({(data_rsci_idat[773:756])
      , 6'b001000});
  assign MultLoop_acc_281_nl = nl_MultLoop_acc_281_nl[23:0];
  assign nl_MultLoop_acc_3295_nl = ({(data_rsci_idat[737:720]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_820_18_8
      , (~ (data_rsci_idat[727:720]))});
  assign MultLoop_acc_3295_nl = nl_MultLoop_acc_3295_nl[19:0];
  assign nl_MultLoop_acc_3296_nl = conv_s2s_24_25({(data_rsci_idat[737:720]) , 6'b000000})
      + conv_s2s_20_25(MultLoop_acc_3295_nl);
  assign MultLoop_acc_3296_nl = nl_MultLoop_acc_3296_nl[24:0];
  assign nl_MultLoop_acc_4427_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_3296_nl)))
      + (~ (data_rsci_idat[737:720]));
  assign MultLoop_acc_4427_nl = nl_MultLoop_acc_4427_nl[17:0];
  assign nl_MultLoop_acc_280_nl = conv_s2s_24_25({(~ (data_rsci_idat[755:738])) ,
      6'b001000}) + conv_s2s_21_25({(~ (data_rsci_idat[755:738])) , 3'b001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_842_18_6
      , (~ (data_rsci_idat[743:738]))});
  assign MultLoop_acc_280_nl = nl_MultLoop_acc_280_nl[24:0];
  assign nl_MultLoop_acc_3375_itm_1  = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_284_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_281_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4427_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_280_nl)));
  assign nl_MultLoop_acc_4429_nl = conv_s2s_10_11(data_rsci_idat[611:602]) + 11'b00000000001;
  assign MultLoop_acc_4429_nl = nl_MultLoop_acc_4429_nl[10:0];
  assign nl_MultLoop_acc_3300_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_17_18({(MultLoop_acc_4429_nl)
      , (data_rsci_idat[601:596])});
  assign MultLoop_acc_3300_nl = nl_MultLoop_acc_3300_nl[17:0];
  assign nl_MultLoop_acc_3301_nl = ({(data_rsci_idat[611:594]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_3300_nl);
  assign MultLoop_acc_3301_nl = nl_MultLoop_acc_3301_nl[21:0];
  assign nl_MultLoop_acc_4430_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3301_nl)))
      + (~ (data_rsci_idat[611:594]));
  assign MultLoop_acc_4430_nl = nl_MultLoop_acc_4430_nl[17:0];
  assign nl_MultLoop_acc_4431_nl =  -conv_s2s_10_11(data_rsci_idat[521:512]);
  assign MultLoop_acc_4431_nl = nl_MultLoop_acc_4431_nl[10:0];
  assign nl_MultLoop_acc_3303_nl = ({(data_rsci_idat[521:504]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4431_nl)
      , (~ (data_rsci_idat[511:504]))});
  assign MultLoop_acc_3303_nl = nl_MultLoop_acc_3303_nl[19:0];
  assign nl_MultLoop_acc_3304_nl = conv_s2s_23_24({(data_rsci_idat[521:504]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_3303_nl);
  assign MultLoop_acc_3304_nl = nl_MultLoop_acc_3304_nl[23:0];
  assign nl_MultLoop_acc_4432_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3304_nl)))
      + (~ (data_rsci_idat[521:504]));
  assign MultLoop_acc_4432_nl = nl_MultLoop_acc_4432_nl[17:0];
  assign nl_MultLoop_acc_3362_itm_1  = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4430_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4432_nl)));
  assign nl_MultLoop_acc_268_nl = conv_s2s_18_26(~ (data_rsci_idat[539:522])) + ({(data_rsci_idat[539:522])
      , 8'b00000001});
  assign MultLoop_acc_268_nl = nl_MultLoop_acc_268_nl[25:0];
  assign nl_MultLoop_acc_4433_nl =  -conv_s2s_10_11(data_rsci_idat[431:422]);
  assign MultLoop_acc_4433_nl = nl_MultLoop_acc_4433_nl[10:0];
  assign nl_MultLoop_acc_3308_nl = ({(data_rsci_idat[431:414]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[431:414])) , 4'b0100}) + conv_s2s_20_24({(~ (data_rsci_idat[431:414]))
      , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4433_nl) , (~ (data_rsci_idat[421:414]))});
  assign MultLoop_acc_3308_nl = nl_MultLoop_acc_3308_nl[23:0];
  assign nl_MultLoop_acc_4434_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3308_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_4434_nl = nl_MultLoop_acc_4434_nl[17:0];
  assign nl_MultLoop_acc_3361_itm_1  = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_268_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4434_nl)));
  assign nl_MultLoop_acc_3309_nl = conv_s2s_18_19(data_rsci_idat[395:378]) + conv_s2s_15_19(data_rsci_idat[395:381]);
  assign MultLoop_acc_3309_nl = nl_MultLoop_acc_3309_nl[18:0];
  assign nl_MultLoop_acc_1165_nl = conv_s2u_19_21(MultLoop_acc_3309_nl) + conv_s2u_20_21({(data_rsci_idat[395:378])
      , 2'b00});
  assign MultLoop_acc_1165_nl = nl_MultLoop_acc_1165_nl[20:0];
  assign nl_MultLoop_acc_4435_nl = conv_s2s_11_12(data_rsci_idat[359:349]) + 12'b000000000001;
  assign MultLoop_acc_4435_nl = nl_MultLoop_acc_4435_nl[11:0];
  assign nl_MultLoop_acc_3311_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_17_18({(MultLoop_acc_4435_nl)
      , (data_rsci_idat[348:344])});
  assign MultLoop_acc_3311_nl = nl_MultLoop_acc_3311_nl[17:0];
  assign nl_MultLoop_acc_3312_nl = ({(data_rsci_idat[359:342]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_3311_nl);
  assign MultLoop_acc_3312_nl = nl_MultLoop_acc_3312_nl[20:0];
  assign nl_MultLoop_acc_259_nl = conv_s2u_21_23(MultLoop_acc_3312_nl) + ({(~ (data_rsci_idat[359:342]))
      , 5'b00000});
  assign MultLoop_acc_259_nl = nl_MultLoop_acc_259_nl[22:0];
  assign nl_MultLoop_acc_4436_nl =  -conv_s2s_11_12(data_rsci_idat[323:313]);
  assign MultLoop_acc_4436_nl = nl_MultLoop_acc_4436_nl[11:0];
  assign nl_MultLoop_acc_3314_nl = ({(data_rsci_idat[323:306]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4436_nl)
      , (~ (data_rsci_idat[312:306]))});
  assign MultLoop_acc_3314_nl = nl_MultLoop_acc_3314_nl[19:0];
  assign nl_MultLoop_acc_3315_nl = conv_s2s_23_24({(data_rsci_idat[323:306]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_3314_nl);
  assign MultLoop_acc_3315_nl = nl_MultLoop_acc_3315_nl[23:0];
  assign nl_MultLoop_acc_4437_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_3315_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_4437_nl = nl_MultLoop_acc_4437_nl[17:0];
  assign nl_MultLoop_acc_3316_nl = conv_s2s_22_23({(~ (data_rsci_idat[287:270]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_3316_nl = nl_MultLoop_acc_3316_nl[22:0];
  assign nl_MultLoop_acc_255_nl = conv_s2s_23_26(MultLoop_acc_3316_nl) + ({(data_rsci_idat[287:270])
      , 8'b00010000});
  assign MultLoop_acc_255_nl = nl_MultLoop_acc_255_nl[25:0];
  assign nl_MultLoop_acc_3373_itm_1  = conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1165_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_259_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4437_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_255_nl)));
  assign nl_MultLoop_acc_3323_nl = conv_s2s_18_19(data_rsci_idat[629:612]) + conv_s2s_15_19(data_rsci_idat[629:615]);
  assign MultLoop_acc_3323_nl = nl_MultLoop_acc_3323_nl[18:0];
  assign nl_MultLoop_acc_1170_nl = conv_s2u_19_23(MultLoop_acc_3323_nl) + conv_s2u_22_23({(data_rsci_idat[629:612])
      , 4'b0000});
  assign MultLoop_acc_1170_nl = nl_MultLoop_acc_1170_nl[22:0];
  assign nl_MultLoop_acc_4440_nl = conv_s2s_10_11(data_rsci_idat[485:476]) + 11'b00000000001;
  assign MultLoop_acc_4440_nl = nl_MultLoop_acc_4440_nl[10:0];
  assign nl_MultLoop_acc_3326_nl = ({(~ (data_rsci_idat[485:468])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[485:468])
      + conv_s2s_16_20({(MultLoop_acc_4440_nl) , (data_rsci_idat[475:471])});
  assign MultLoop_acc_3326_nl = nl_MultLoop_acc_3326_nl[19:0];
  assign nl_MultLoop_acc_1168_nl = conv_s2u_20_24(MultLoop_acc_3326_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[485:468])) , 5'b00100});
  assign MultLoop_acc_1168_nl = nl_MultLoop_acc_1168_nl[23:0];
  assign nl_MultLoop_acc_4438_nl =  -conv_s2s_13_14(data_rsci_idat[233:221]);
  assign MultLoop_acc_4438_nl = nl_MultLoop_acc_4438_nl[13:0];
  assign nl_MultLoop_acc_3318_nl = ({(data_rsci_idat[233:216]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4438_nl)
      , (~ (data_rsci_idat[220:216]))});
  assign MultLoop_acc_3318_nl = nl_MultLoop_acc_3318_nl[20:0];
  assign nl_MultLoop_acc_252_nl = conv_s2s_21_23(MultLoop_acc_3318_nl) + ({(~ (data_rsci_idat[233:216]))
      , 5'b00000});
  assign MultLoop_acc_252_nl = nl_MultLoop_acc_252_nl[22:0];
  assign nl_MultLoop_acc_3320_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_17_18({MultLoop_acc_3941_cse_1
      , (data_rsci_idat[240:236])});
  assign MultLoop_acc_3320_nl = nl_MultLoop_acc_3320_nl[17:0];
  assign nl_MultLoop_acc_1162_nl = conv_s2u_18_24(MultLoop_acc_3320_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[251:234])) , 5'b00001});
  assign MultLoop_acc_1162_nl = nl_MultLoop_acc_1162_nl[23:0];
  assign nl_MultLoop_acc_3321_nl = (~ (data_rsci_idat[215:198])) + conv_s2s_14_18(data_rsci_idat[215:202]);
  assign MultLoop_acc_3321_nl = nl_MultLoop_acc_3321_nl[17:0];
  assign nl_MultLoop_acc_1161_nl = conv_s2u_18_20(MultLoop_acc_3321_nl) + ({(data_rsci_idat[215:198])
      , 2'b01});
  assign MultLoop_acc_1161_nl = nl_MultLoop_acc_1161_nl[19:0];
  assign nl_MultLoop_acc_4694_nl = conv_s2u_19_22(MultLoop_acc_4690[22:4]) + ({(data_rsci_idat[161:144])
      , 4'b0001});
  assign MultLoop_acc_4694_nl = nl_MultLoop_acc_4694_nl[21:0];
  assign nl_MultLoop_acc_3379_itm_1  = conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1170_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1168_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_252_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1162_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1161_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_4694_nl)));
  assign nl_MultLoop_acc_4668_nl = conv_s2u_19_23(MultLoop_acc_1957_cse_1[20:2])
      + conv_s2u_22_23({(~ (data_rsci_idat[647:630])) , 4'b0001});
  assign MultLoop_acc_4668_nl = nl_MultLoop_acc_4668_nl[22:0];
  assign nl_MultLoop_acc_4066_nl = conv_s2s_11_12(data_rsci_idat[575:565]) + 12'b000000000001;
  assign MultLoop_acc_4066_nl = nl_MultLoop_acc_4066_nl[11:0];
  assign nl_MultLoop_acc_2177_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_17_18({(MultLoop_acc_4066_nl)
      , (data_rsci_idat[564:560])});
  assign MultLoop_acc_2177_nl = nl_MultLoop_acc_2177_nl[17:0];
  assign nl_MultLoop_acc_2178_nl = conv_s2s_20_21({(~ (data_rsci_idat[575:558]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2177_nl);
  assign MultLoop_acc_2178_nl = nl_MultLoop_acc_2178_nl[20:0];
  assign nl_MultLoop_acc_1356_nl = conv_s2u_21_24(MultLoop_acc_2178_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[575:558])) , 5'b00100});
  assign MultLoop_acc_1356_nl = nl_MultLoop_acc_1356_nl[23:0];
  assign nl_MultLoop_acc_2182_nl = ({(~ (data_rsci_idat[431:414])) , 4'b0000}) +
      conv_s2s_20_22({(data_rsci_idat[431:414]) , 2'b00}) + conv_s2s_18_22(data_rsci_idat[431:414])
      + conv_s2s_17_22({MultLoop_MultLoop_conc_680_16_6 , (data_rsci_idat[421:416])});
  assign MultLoop_acc_2182_nl = nl_MultLoop_acc_2182_nl[21:0];
  assign nl_MultLoop_acc_1352_nl = conv_s2u_22_25(MultLoop_acc_2182_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[431:414])) , 6'b010000});
  assign MultLoop_acc_1352_nl = nl_MultLoop_acc_1352_nl[24:0];
  assign nl_MultLoop_acc_2173_nl = ({(data_rsci_idat[89:72]) , 5'b00001}) + conv_s2s_18_23(~
      (data_rsci_idat[89:72]));
  assign MultLoop_acc_2173_nl = nl_MultLoop_acc_2173_nl[22:0];
  assign nl_MultLoop_acc_4064_nl = conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_2173_nl)))
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_4064_nl = nl_MultLoop_acc_4064_nl[18:0];
  assign nl_MultLoop_acc_806_nl = (MultLoop_acc_807_itm_21_6[15:1]) + 15'b000000010100101;
  assign MultLoop_acc_806_nl = nl_MultLoop_acc_806_nl[14:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_96_itm_1  =
      conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_4668_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1356_nl)))
      + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1352_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4064_nl)))
      + conv_s2s_16_18({(MultLoop_acc_806_nl) , (MultLoop_acc_807_itm_21_6[0])});
  assign nl_MultLoop_acc_828_nl = conv_s2s_25_26({(~ (data_rsci_idat[395:378])) ,
      7'b0010000}) + conv_s2s_22_26({(~ (data_rsci_idat[395:378])) , 4'b0100}) +
      conv_s2s_20_26({(~ (data_rsci_idat[395:378])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_818_18_7
      , (~ (data_rsci_idat[384:378]))});
  assign MultLoop_acc_828_nl = nl_MultLoop_acc_828_nl[25:0];
  assign nl_MultLoop_acc_4069_nl =  -conv_s2s_13_14(data_rsci_idat[269:257]);
  assign MultLoop_acc_4069_nl = nl_MultLoop_acc_4069_nl[13:0];
  assign nl_MultLoop_acc_821_nl = conv_s2s_23_24({(~ (data_rsci_idat[269:252])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[269:252])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4069_nl)
      , (~ (data_rsci_idat[256:252]))});
  assign MultLoop_acc_821_nl = nl_MultLoop_acc_821_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_86_itm_1  =
      conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_828_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_821_nl)));
  assign nl_MultLoop_acc_4070_nl =  -conv_s2s_13_14(data_rsci_idat[161:149]);
  assign MultLoop_acc_4070_nl = nl_MultLoop_acc_4070_nl[13:0];
  assign nl_MultLoop_acc_815_nl = conv_s2s_23_24({(~ (data_rsci_idat[161:144])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[161:144])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4070_nl)
      , (~ (data_rsci_idat[148:144]))});
  assign MultLoop_acc_815_nl = nl_MultLoop_acc_815_nl[23:0];
  assign nl_MultLoop_acc_4071_nl = conv_s2s_14_15(data_rsci_idat[845:832]) + 15'b000000000000001;
  assign MultLoop_acc_4071_nl = nl_MultLoop_acc_4071_nl[14:0];
  assign nl_MultLoop_acc_2129_nl = conv_s2s_18_19(data_rsci_idat[845:828]) + conv_s2s_17_19({(MultLoop_acc_4071_nl)
      , (data_rsci_idat[831:830])});
  assign MultLoop_acc_2129_nl = nl_MultLoop_acc_2129_nl[18:0];
  assign nl_MultLoop_acc_852_nl = conv_s2u_19_20(MultLoop_acc_2129_nl) + ({(~ (data_rsci_idat[845:828]))
      , 2'b00});
  assign MultLoop_acc_852_nl = nl_MultLoop_acc_852_nl[19:0];
  assign nl_MultLoop_acc_2127_nl = conv_s2s_20_21({(~ (data_rsci_idat[71:54])) ,
      2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_2127_nl = nl_MultLoop_acc_2127_nl[20:0];
  assign nl_MultLoop_acc_810_nl = conv_s2s_21_22(MultLoop_acc_2127_nl) + ({(data_rsci_idat[71:54])
      , 4'b0100});
  assign MultLoop_acc_810_nl = nl_MultLoop_acc_810_nl[21:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_7_nl = ~((data_rsci_idat[435:432]!=4'b0000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl = conv_s2s_13_14(readslicef_20_13_7((MultLoop_acc_852_nl)))
      + conv_s2s_12_14(readslicef_22_12_10((MultLoop_acc_810_nl))) + conv_u2s_1_14(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_7_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl[13:0];
  assign nl_MultLoop_acc_1361_nl = conv_s2u_15_19(data_rsci_idat[863:849]) + conv_s2u_18_19(data_rsci_idat[863:846]);
  assign MultLoop_acc_1361_nl = nl_MultLoop_acc_1361_nl[18:0];
  assign nl_MultLoop_acc_848_nl = conv_s2s_23_24({(~ (data_rsci_idat[773:756])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[773:756])) , 3'b001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_760_18_5
      , (~ (data_rsci_idat[760:756]))});
  assign MultLoop_acc_848_nl = nl_MultLoop_acc_848_nl[23:0];
  assign nl_MultLoop_acc_4073_nl =  -conv_s2s_14_15(data_rsci_idat[593:580]);
  assign MultLoop_acc_4073_nl = nl_MultLoop_acc_4073_nl[14:0];
  assign nl_MultLoop_acc_838_nl = conv_s2s_19_23({(MultLoop_acc_4073_nl) , (~ (data_rsci_idat[579:576]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[593:576])) , 4'b0001});
  assign MultLoop_acc_838_nl = nl_MultLoop_acc_838_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_71_itm_1  =
      conv_s2s_14_16(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_57_nl)
      + conv_s2s_14_16(readslicef_19_14_5((MultLoop_acc_1361_nl))) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_848_nl)))
      + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_838_nl)));
  assign nl_MultLoop_acc_1355_nl = conv_s2u_18_20(MultLoop_acc_2133_cse_1) + ({(data_rsci_idat[521:504])
      , 2'b01});
  assign MultLoop_acc_1355_nl = nl_MultLoop_acc_1355_nl[19:0];
  assign nl_MultLoop_acc_1353_nl = conv_s2u_16_19(data_rsci_idat[467:452]) + conv_s2u_18_19(data_rsci_idat[467:450]);
  assign MultLoop_acc_1353_nl = nl_MultLoop_acc_1353_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_70_itm_1  =
      conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_1355_nl))) + conv_s2s_14_16(MultLoop_acc_785_itm_17_4)
      + conv_s2s_14_16(~ (data_rsci_idat[449:436])) + conv_s2s_14_16(readslicef_19_14_5((MultLoop_acc_1353_nl)));
  assign nl_MultLoop_acc_851_nl = conv_s2s_18_21(~ (data_rsci_idat[827:810])) + ({(data_rsci_idat[827:810])
      , 3'b001});
  assign MultLoop_acc_851_nl = nl_MultLoop_acc_851_nl[20:0];
  assign nl_MultLoop_acc_4074_nl =  -conv_s2s_13_14(data_rsci_idat[323:311]);
  assign MultLoop_acc_4074_nl = nl_MultLoop_acc_4074_nl[13:0];
  assign nl_MultLoop_acc_824_nl = conv_s2s_23_24({(~ (data_rsci_idat[323:306])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[323:306])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4074_nl)
      , (~ (data_rsci_idat[310:306]))});
  assign MultLoop_acc_824_nl = nl_MultLoop_acc_824_nl[23:0];
  assign nl_MultLoop_acc_2137_nl = conv_s2s_18_19(data_rsci_idat[287:270]) + conv_s2s_16_19({MultLoop_acc_4075_cse_1
      , (data_rsci_idat[275:273])});
  assign MultLoop_acc_2137_nl = nl_MultLoop_acc_2137_nl[18:0];
  assign nl_MultLoop_acc_822_nl = conv_s2u_19_21(MultLoop_acc_2137_nl) + ({(~ (data_rsci_idat[287:270]))
      , 3'b000});
  assign MultLoop_acc_822_nl = nl_MultLoop_acc_822_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_69_itm_1  =
      conv_s2s_15_16(readslicef_21_15_6((MultLoop_acc_851_nl))) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_824_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_822_nl)));
  assign nl_MultLoop_acc_2139_nl = conv_s2s_18_19(data_rsci_idat[755:738]) + conv_s2s_16_19({MultLoop_acc_4076_cse_1
      , (data_rsci_idat[743:741])});
  assign MultLoop_acc_2139_nl = nl_MultLoop_acc_2139_nl[18:0];
  assign nl_MultLoop_acc_847_nl = conv_s2u_19_21(MultLoop_acc_2139_nl) + ({(~ (data_rsci_idat[755:738]))
      , 3'b000});
  assign MultLoop_acc_847_nl = nl_MultLoop_acc_847_nl[20:0];
  assign nl_MultLoop_acc_2141_nl = ({(data_rsci_idat[683:666]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_816_18_7
      , (~ (data_rsci_idat[672:666]))});
  assign MultLoop_acc_2141_nl = nl_MultLoop_acc_2141_nl[20:0];
  assign nl_MultLoop_acc_4078_nl = conv_s2u_14_18(readslicef_21_14_7((MultLoop_acc_2141_nl)))
      + (~ (data_rsci_idat[683:666]));
  assign MultLoop_acc_4078_nl = nl_MultLoop_acc_4078_nl[17:0];
  assign nl_MultLoop_acc_2144_nl = ({(data_rsci_idat[557:540]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[557:540])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_700_18_7
      , (~ (data_rsci_idat[546:540]))});
  assign MultLoop_acc_2144_nl = nl_MultLoop_acc_2144_nl[21:0];
  assign nl_MultLoop_acc_4080_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_2144_nl)))
      + (~ (data_rsci_idat[557:540]));
  assign MultLoop_acc_4080_nl = nl_MultLoop_acc_4080_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_83_itm_1  =
      conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_847_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4078_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4080_nl))) + conv_s2s_15_17(MultLoop_acc_1350_itm_22_7[15:1]);
  assign nl_MultLoop_acc_4614_nl = conv_s2u_15_19(MultLoop_acc_2145_itm_20_5[15:1])
      + conv_s2u_18_19(data_rsci_idat[233:216]);
  assign MultLoop_acc_4614_nl = nl_MultLoop_acc_4614_nl[18:0];
  assign nl_MultLoop_acc_1348_nl = conv_s2u_12_19(data_rsci_idat[215:204]) + conv_s2u_18_19(data_rsci_idat[215:198]);
  assign MultLoop_acc_1348_nl = nl_MultLoop_acc_1348_nl[18:0];
  assign nl_MultLoop_acc_2147_nl = ({(~ (data_rsci_idat[179:162])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[179:162])
      + conv_s2s_15_20(data_rsci_idat[179:165]);
  assign MultLoop_acc_2147_nl = nl_MultLoop_acc_2147_nl[19:0];
  assign nl_MultLoop_acc_1347_nl = conv_s2u_20_22(MultLoop_acc_2147_nl) + ({(data_rsci_idat[179:162])
      , 4'b0100});
  assign MultLoop_acc_1347_nl = nl_MultLoop_acc_1347_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_82_itm_1  =
      conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4614_nl))) + conv_s2s_15_17(MultLoop_acc_579_itm_19_4[15:1])
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_1348_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1347_nl)));
  assign nl_MultLoop_acc_4081_nl =  -conv_s2s_15_16(data_rsci_idat[143:129]);
  assign MultLoop_acc_4081_nl = nl_MultLoop_acc_4081_nl[15:0];
  assign nl_MultLoop_acc_814_nl = conv_s2s_19_22({(MultLoop_acc_4081_nl) , (~ (data_rsci_idat[128:126]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[143:126])) , 3'b001});
  assign MultLoop_acc_814_nl = nl_MultLoop_acc_814_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_64_itm_1  =
      conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_814_nl))) + conv_s2s_15_16(MultLoop_acc_528_itm_24_10);
  assign nl_MultLoop_acc_2149_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_16_18(data_rsci_idat[53:38]);
  assign MultLoop_acc_2149_nl = nl_MultLoop_acc_2149_nl[17:0];
  assign nl_MultLoop_acc_1345_nl = conv_s2u_18_22(MultLoop_acc_2149_nl) + ({(data_rsci_idat[53:36])
      , 4'b0001});
  assign MultLoop_acc_1345_nl = nl_MultLoop_acc_1345_nl[21:0];
  assign nl_MultLoop_acc_4082_nl =  -conv_s2s_16_17(data_rsci_idat[35:20]);
  assign MultLoop_acc_4082_nl = nl_MultLoop_acc_4082_nl[16:0];
  assign nl_MultLoop_acc_808_nl = conv_s2s_19_21({(MultLoop_acc_4082_nl) , (~ (data_rsci_idat[19:18]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[35:18])) , 2'b01});
  assign MultLoop_acc_808_nl = nl_MultLoop_acc_808_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_63_itm_1  =
      conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_1345_nl))) + conv_s2s_15_16(readslicef_21_15_6((MultLoop_acc_808_nl)));
  assign nl_MultLoop_acc_4615_nl = conv_s2u_14_19(MultLoop_acc_1479_itm_18_3[15:2])
      + conv_s2u_18_19(data_rsci_idat[809:792]);
  assign MultLoop_acc_4615_nl = nl_MultLoop_acc_4615_nl[18:0];
  assign nl_MultLoop_acc_2154_nl = conv_s2s_20_21({(data_rsci_idat[791:774]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[791:774]) + conv_s2s_16_21({MultLoop_acc_4083_cse_1
      , (data_rsci_idat[780:777])});
  assign MultLoop_acc_2154_nl = nl_MultLoop_acc_2154_nl[20:0];
  assign nl_MultLoop_acc_849_nl = conv_s2u_21_22(MultLoop_acc_2154_nl) + ({(~ (data_rsci_idat[791:774]))
      , 4'b0000});
  assign MultLoop_acc_849_nl = nl_MultLoop_acc_849_nl[21:0];
  assign nl_MultLoop_acc_2155_nl = ({(data_rsci_idat[737:720]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[737:720]));
  assign MultLoop_acc_2155_nl = nl_MultLoop_acc_2155_nl[19:0];
  assign nl_MultLoop_acc_2156_nl = ({(~ (data_rsci_idat[737:720])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2155_nl);
  assign MultLoop_acc_2156_nl = nl_MultLoop_acc_2156_nl[21:0];
  assign nl_MultLoop_acc_846_nl = conv_s2s_22_24(MultLoop_acc_2156_nl) + ({(data_rsci_idat[737:720])
      , 6'b010000});
  assign MultLoop_acc_846_nl = nl_MultLoop_acc_846_nl[23:0];
  assign nl_MultLoop_acc_2158_nl = conv_s2s_18_19(data_rsci_idat[629:612]) + conv_s2s_16_19({MultLoop_acc_4084_cse_1
      , (data_rsci_idat[619:615])});
  assign MultLoop_acc_2158_nl = nl_MultLoop_acc_2158_nl[18:0];
  assign nl_MultLoop_acc_840_nl = conv_s2u_19_23(MultLoop_acc_2158_nl) + ({(~ (data_rsci_idat[629:612]))
      , 5'b00000});
  assign MultLoop_acc_840_nl = nl_MultLoop_acc_840_nl[22:0];
  assign nl_MultLoop_acc_2161_nl = ({(~ (data_rsci_idat[611:594])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[611:594])
      + conv_s2s_16_20({MultLoop_MultLoop_conc_776_15_4 , (data_rsci_idat[600:597])});
  assign MultLoop_acc_2161_nl = nl_MultLoop_acc_2161_nl[19:0];
  assign nl_MultLoop_acc_1357_nl = conv_s2u_20_23(MultLoop_acc_2161_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[611:594])) , 4'b0100});
  assign MultLoop_acc_1357_nl = nl_MultLoop_acc_1357_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_98_itm_1  =
      conv_s2s_16_18(MultLoop_acc_4593_itm_18_3) + conv_s2s_16_18(MultLoop_acc_2073_cse_1[18:3])
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4615_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_849_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_846_nl))) + conv_s2s_16_18(MultLoop_acc_4592_itm_18_3)
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_840_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1357_nl)));
  assign nl_MultLoop_acc_2170_nl = (~ (data_rsci_idat[305:288])) + conv_s2s_16_18({MultLoop_acc_3989_cse_1
      , (data_rsci_idat[295:291])});
  assign MultLoop_acc_2170_nl = nl_MultLoop_acc_2170_nl[17:0];
  assign nl_MultLoop_acc_2171_nl = ({(data_rsci_idat[305:288]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2170_nl);
  assign MultLoop_acc_2171_nl = nl_MultLoop_acc_2171_nl[19:0];
  assign nl_MultLoop_acc_823_nl = conv_s2u_20_23(MultLoop_acc_2171_nl) + ({(~ (data_rsci_idat[305:288]))
      , 5'b00000});
  assign MultLoop_acc_823_nl = nl_MultLoop_acc_823_nl[22:0];
  assign nl_MultLoop_acc_4086_nl =  -conv_s2s_11_12(data_rsci_idat[539:529]);
  assign MultLoop_acc_4086_nl = nl_MultLoop_acc_4086_nl[11:0];
  assign nl_MultLoop_acc_835_nl = conv_s2s_25_26({(~ (data_rsci_idat[539:522])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[539:522])) , 5'b00001}) +
      conv_s2s_19_26({(MultLoop_acc_4086_nl) , (~ (data_rsci_idat[528:522]))});
  assign MultLoop_acc_835_nl = nl_MultLoop_acc_835_nl[25:0];
  assign nl_MultLoop_acc_2165_nl = (~ (data_rsci_idat[485:468])) + conv_s2s_17_18({MultLoop_MultLoop_conc_860_16_4
      , (data_rsci_idat[473:470])});
  assign MultLoop_acc_2165_nl = nl_MultLoop_acc_2165_nl[17:0];
  assign nl_MultLoop_acc_1354_nl = conv_s2u_18_23(MultLoop_acc_2165_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[485:468])) , 4'b0001});
  assign MultLoop_acc_1354_nl = nl_MultLoop_acc_1354_nl[22:0];
  assign nl_MultLoop_acc_4088_nl = conv_s2s_11_12(data_rsci_idat[413:403]) + 12'b000000000001;
  assign MultLoop_acc_4088_nl = nl_MultLoop_acc_4088_nl[11:0];
  assign nl_MultLoop_acc_2168_nl = ({(~ (data_rsci_idat[413:396])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[413:396])
      + conv_s2s_16_20({(MultLoop_acc_4088_nl) , (data_rsci_idat[402:399])});
  assign MultLoop_acc_2168_nl = nl_MultLoop_acc_2168_nl[19:0];
  assign nl_MultLoop_acc_1351_nl = conv_s2u_20_23(MultLoop_acc_2168_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[413:396])) , 4'b0100});
  assign MultLoop_acc_1351_nl = nl_MultLoop_acc_1351_nl[22:0];
  assign nl_MultLoop_acc_1349_nl = conv_s2u_16_19(data_rsci_idat[341:326]) + conv_s2u_18_19(data_rsci_idat[341:324]);
  assign MultLoop_acc_1349_nl = nl_MultLoop_acc_1349_nl[18:0];
  assign nl_MultLoop_acc_4616_nl = conv_s2u_19_20(MultLoop_acc_1735_cse_1[20:2])
      + ({(data_rsci_idat[251:234]) , 2'b01});
  assign MultLoop_acc_4616_nl = nl_MultLoop_acc_4616_nl[19:0];
  assign nl_MultLoop_acc_1346_nl = conv_s2u_11_19(data_rsci_idat[125:115]) + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_1346_nl = nl_MultLoop_acc_1346_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_97_itm_1  =
      conv_s2s_16_18(MultLoop_acc_826_itm_25_10) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_823_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_835_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1354_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1351_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1349_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_4616_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1346_nl)));
  assign nl_MultLoop_acc_3207_nl = ({(~ (data_rsci_idat[557:540])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_788_cse_1);
  assign MultLoop_acc_3207_nl = nl_MultLoop_acc_3207_nl[22:0];
  assign nl_MultLoop_acc_317_nl = conv_s2s_23_25(MultLoop_acc_3207_nl) + ({(data_rsci_idat[557:540])
      , 7'b0100000});
  assign MultLoop_acc_317_nl = nl_MultLoop_acc_317_nl[24:0];
  assign nl_MultLoop_acc_3209_nl = ({(~ (data_rsci_idat[503:486])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2923_cse_1);
  assign MultLoop_acc_3209_nl = nl_MultLoop_acc_3209_nl[21:0];
  assign nl_MultLoop_acc_3210_nl = ({(data_rsci_idat[503:486]) , 6'b010000}) + conv_s2s_22_24(MultLoop_acc_3209_nl);
  assign MultLoop_acc_3210_nl = nl_MultLoop_acc_3210_nl[23:0];
  assign nl_MultLoop_acc_4401_nl = conv_s2u_16_19(readslicef_24_16_8((MultLoop_acc_3210_nl)))
      + conv_s2u_18_19(data_rsci_idat[503:486]);
  assign MultLoop_acc_4401_nl = nl_MultLoop_acc_4401_nl[18:0];
  assign nl_MultLoop_acc_4639_nl = conv_s2u_18_19(data_rsci_idat[233:216]) + conv_s2u_16_19(MultLoop_acc_2145_itm_20_5);
  assign MultLoop_acc_4639_nl = nl_MultLoop_acc_4639_nl[18:0];
  assign nl_MultLoop_acc_4402_nl = conv_s2u_16_19(readslicef_19_16_3((MultLoop_acc_4639_nl)))
      + conv_s2u_18_19(data_rsci_idat[233:216]);
  assign MultLoop_acc_4402_nl = nl_MultLoop_acc_4402_nl[18:0];
  assign nl_MultLoop_acc_4640_nl = conv_s2u_22_23({(~ (data_rsci_idat[251:234]))
      , 4'b0001}) + conv_s2u_19_23(MultLoop_acc_3213_itm_21_3_1);
  assign MultLoop_acc_4640_nl = nl_MultLoop_acc_4640_nl[22:0];
  assign nl_MultLoop_acc_4403_nl = conv_s2u_19_20(readslicef_23_19_4((MultLoop_acc_4640_nl)))
      + ({(data_rsci_idat[251:234]) , 2'b01});
  assign MultLoop_acc_4403_nl = nl_MultLoop_acc_4403_nl[19:0];
  assign nl_MultLoop_acc_3259_nl = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_317_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4401_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4402_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_4403_nl)));
  assign MultLoop_acc_3259_nl = nl_MultLoop_acc_3259_nl[17:0];
  assign nl_MultLoop_acc_4399_nl = conv_s2s_12_13(data_rsci_idat[269:258]) + 13'b0000000000001;
  assign MultLoop_acc_4399_nl = nl_MultLoop_acc_4399_nl[12:0];
  assign nl_MultLoop_acc_3200_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_15_18({(MultLoop_acc_4399_nl)
      , (data_rsci_idat[257:256])});
  assign MultLoop_acc_3200_nl = nl_MultLoop_acc_3200_nl[17:0];
  assign nl_MultLoop_acc_1180_nl = conv_s2u_18_21(MultLoop_acc_3200_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[269:252])) , 2'b01});
  assign MultLoop_acc_1180_nl = nl_MultLoop_acc_1180_nl[20:0];
  assign nl_MultLoop_acc_3204_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_15_18(data_rsci_idat[755:741]);
  assign MultLoop_acc_3204_nl = nl_MultLoop_acc_3204_nl[17:0];
  assign nl_MultLoop_acc_3205_nl = ({(data_rsci_idat[755:738]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_3204_nl);
  assign MultLoop_acc_3205_nl = nl_MultLoop_acc_3205_nl[20:0];
  assign nl_MultLoop_acc_1193_nl = conv_s2u_21_24(MultLoop_acc_3205_nl) + conv_s2u_23_24({(data_rsci_idat[755:738])
      , 5'b00000});
  assign MultLoop_acc_1193_nl = nl_MultLoop_acc_1193_nl[23:0];
  assign nl_MultLoop_acc_324_nl = conv_s2u_14_18(data_rsci_idat[683:670]) - (data_rsci_idat[683:666]);
  assign MultLoop_acc_324_nl = nl_MultLoop_acc_324_nl[17:0];
  assign nl_MultLoop_acc_4400_nl = conv_s2s_12_13(data_rsci_idat[161:150]) + 13'b0000000000001;
  assign MultLoop_acc_4400_nl = nl_MultLoop_acc_4400_nl[12:0];
  assign nl_MultLoop_acc_3202_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_17_18({(MultLoop_acc_4400_nl)
      , (data_rsci_idat[149:146])});
  assign MultLoop_acc_3202_nl = nl_MultLoop_acc_3202_nl[17:0];
  assign nl_MultLoop_acc_1178_nl = conv_s2u_18_23(MultLoop_acc_3202_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[161:144])) , 4'b0001});
  assign MultLoop_acc_1178_nl = nl_MultLoop_acc_1178_nl[22:0];
  assign nl_MultLoop_acc_3203_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_16_18(data_rsci_idat[107:92]);
  assign MultLoop_acc_3203_nl = nl_MultLoop_acc_3203_nl[17:0];
  assign nl_MultLoop_acc_1176_nl = conv_s2u_18_21(MultLoop_acc_3203_nl) + ({(data_rsci_idat[107:90])
      , 3'b001});
  assign MultLoop_acc_1176_nl = nl_MultLoop_acc_1176_nl[20:0];
  assign nl_MultLoop_acc_3264_itm_1  = (MultLoop_acc_3259_nl) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1180_nl)))
      + conv_s2s_16_18(MultLoop_acc_2057_cse_1[18:3]) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1193_nl)))
      + conv_s2s_16_18(MultLoop_acc_1753_itm_19_4) + conv_s2s_14_18(MultLoop_acc_334_itm_20_5[15:2])
      + conv_s2s_14_18(readslicef_18_14_4((MultLoop_acc_324_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1178_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1176_nl)));
  assign nl_MultLoop_acc_4641_nl = conv_s2u_13_19(MultLoop_acc_2412_cse_1[18:6])
      + conv_s2u_18_19(data_rsci_idat[125:108]);
  assign MultLoop_acc_4641_nl = nl_MultLoop_acc_4641_nl[18:0];
  assign nl_MultLoop_acc_3217_nl = ({(data_rsci_idat[143:126]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[143:126])) , 2'b01}) + conv_s2s_18_22(~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_3217_nl = nl_MultLoop_acc_3217_nl[21:0];
  assign nl_MultLoop_acc_4404_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_3217_nl)))
      + conv_s2u_18_19(data_rsci_idat[143:126]);
  assign MultLoop_acc_4404_nl = nl_MultLoop_acc_4404_nl[18:0];
  assign nl_MultLoop_acc_4642_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_1485_cse_1[20:2]);
  assign MultLoop_acc_4642_nl = nl_MultLoop_acc_4642_nl[19:0];
  assign nl_MultLoop_acc_4405_nl = conv_s2u_14_19(readslicef_20_14_6((MultLoop_acc_4642_nl)))
      + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_4405_nl = nl_MultLoop_acc_4405_nl[18:0];
  assign nl_MultLoop_acc_3220_nl = (~ (data_rsci_idat[71:54])) + conv_s2s_16_18(data_rsci_idat[71:56]);
  assign MultLoop_acc_3220_nl = nl_MultLoop_acc_3220_nl[17:0];
  assign nl_MultLoop_acc_3221_nl = conv_s2s_20_21({(~ (data_rsci_idat[71:54])) ,
      2'b01}) + conv_s2s_18_21(MultLoop_acc_3220_nl);
  assign MultLoop_acc_3221_nl = nl_MultLoop_acc_3221_nl[20:0];
  assign nl_MultLoop_acc_1175_nl = conv_s2u_21_22(MultLoop_acc_3221_nl) + ({(data_rsci_idat[71:54])
      , 4'b0100});
  assign MultLoop_acc_1175_nl = nl_MultLoop_acc_1175_nl[21:0];
  assign nl_MultLoop_acc_3258_itm_1  = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4641_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4404_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4405_nl)))
      + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1175_nl)));
  assign nl_MultLoop_acc_3161_nl = ({(data_rsci_idat[647:630]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_834_18_5
      , (~ (data_rsci_idat[634:630]))});
  assign MultLoop_acc_3161_nl = nl_MultLoop_acc_3161_nl[20:0];
  assign nl_MultLoop_acc_322_nl = conv_s2s_21_23(MultLoop_acc_3161_nl) + ({(~ (data_rsci_idat[647:630]))
      , 5'b00000});
  assign MultLoop_acc_322_nl = nl_MultLoop_acc_322_nl[22:0];
  assign nl_MultLoop_acc_308_nl = conv_s2s_18_23(~ (data_rsci_idat[377:360])) + ({(data_rsci_idat[377:360])
      , 5'b00001});
  assign MultLoop_acc_308_nl = nl_MultLoop_acc_308_nl[22:0];
  assign nl_MultLoop_acc_3162_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_14_18(data_rsci_idat[179:166]);
  assign MultLoop_acc_3162_nl = nl_MultLoop_acc_3162_nl[17:0];
  assign nl_MultLoop_acc_1179_nl = conv_s2u_18_20(MultLoop_acc_3162_nl) + ({(data_rsci_idat[179:162])
      , 2'b01});
  assign MultLoop_acc_1179_nl = nl_MultLoop_acc_1179_nl[19:0];
  assign nl_MultLoop_acc_310_nl = conv_s2u_15_18(data_rsci_idat[413:399]) - (data_rsci_idat[413:396]);
  assign MultLoop_acc_310_nl = nl_MultLoop_acc_310_nl[17:0];
  assign nl_MultLoop_acc_288_nl = (MultLoop_acc_3683_itm_18_3_1[15:8]) + 8'b00011111;
  assign MultLoop_acc_288_nl = nl_MultLoop_acc_288_nl[7:0];
  assign nl_MultLoop_acc_3233_itm_1  = conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_322_nl)))
      + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_308_nl))) + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_1179_nl)))
      + conv_s2s_11_16(readslicef_18_11_7((MultLoop_acc_310_nl))) + conv_s2s_11_16(data_rsci_idat[215:205])
      + conv_s2s_11_16({(MultLoop_acc_288_nl) , (MultLoop_acc_3683_itm_18_3_1[7:5])});
  assign nl_MultLoop_acc_3164_nl = ({(data_rsci_idat[773:756]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_688_18_7
      , (~ (data_rsci_idat[762:756]))});
  assign MultLoop_acc_3164_nl = nl_MultLoop_acc_3164_nl[19:0];
  assign nl_MultLoop_acc_4408_nl = conv_s2u_13_18(readslicef_20_13_7((MultLoop_acc_3164_nl)))
      + (~ (data_rsci_idat[773:756]));
  assign MultLoop_acc_4408_nl = nl_MultLoop_acc_4408_nl[17:0];
  assign nl_MultLoop_acc_3232_itm_1  = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4408_nl)))
      + conv_s2s_15_16(MultLoop_acc_1191_itm_21_7);
  assign nl_MultLoop_acc_3166_nl = ({(~ (data_rsci_idat[737:720])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2522_cse_1);
  assign MultLoop_acc_3166_nl = nl_MultLoop_acc_3166_nl[19:0];
  assign nl_MultLoop_acc_1192_nl = conv_s2u_20_22(MultLoop_acc_3166_nl) + ({(data_rsci_idat[737:720])
      , 4'b0100});
  assign MultLoop_acc_1192_nl = nl_MultLoop_acc_1192_nl[21:0];
  assign nl_MultLoop_acc_321_nl = conv_s2u_13_18(data_rsci_idat[629:617]) - (data_rsci_idat[629:612]);
  assign MultLoop_acc_321_nl = nl_MultLoop_acc_321_nl[17:0];
  assign nl_MultLoop_acc_3167_nl = ({(data_rsci_idat[539:522]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[539:522]));
  assign MultLoop_acc_3167_nl = nl_MultLoop_acc_3167_nl[19:0];
  assign nl_MultLoop_acc_3168_nl = ({(~ (data_rsci_idat[539:522])) , 5'b00000}) +
      conv_s2s_20_23(MultLoop_acc_3167_nl);
  assign MultLoop_acc_3168_nl = nl_MultLoop_acc_3168_nl[22:0];
  assign nl_MultLoop_acc_316_nl = conv_s2s_23_25(MultLoop_acc_3168_nl) + ({(data_rsci_idat[539:522])
      , 7'b0100000});
  assign MultLoop_acc_316_nl = nl_MultLoop_acc_316_nl[24:0];
  assign nl_MultLoop_acc_4643_nl = conv_s2u_17_19(MultLoop_acc_2967_cse_1[18:2])
      + conv_s2u_18_19(data_rsci_idat[521:504]);
  assign MultLoop_acc_4643_nl = nl_MultLoop_acc_4643_nl[18:0];
  assign nl_MultLoop_acc_3245_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1192_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_321_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_316_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4643_nl)));
  assign nl_MultLoop_acc_3174_nl = conv_s2s_20_21({(data_rsci_idat[845:828]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[845:828]) + conv_s2s_15_21(data_rsci_idat[845:831]);
  assign MultLoop_acc_3174_nl = nl_MultLoop_acc_3174_nl[20:0];
  assign nl_MultLoop_acc_1194_nl = conv_s2u_21_23(MultLoop_acc_3174_nl) + conv_s2u_22_23({(data_rsci_idat[845:828])
      , 4'b0000});
  assign MultLoop_acc_1194_nl = nl_MultLoop_acc_1194_nl[22:0];
  assign nl_MultLoop_acc_4409_nl =  -conv_s2s_15_16(data_rsci_idat[35:21]);
  assign MultLoop_acc_4409_nl = nl_MultLoop_acc_4409_nl[15:0];
  assign nl_MultLoop_acc_290_nl = conv_s2s_19_22({(MultLoop_acc_4409_nl) , (~ (data_rsci_idat[20:18]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[35:18])) , 3'b001});
  assign MultLoop_acc_290_nl = nl_MultLoop_acc_290_nl[21:0];
  assign nl_MultLoop_acc_4410_nl =  -conv_s2s_12_13(data_rsci_idat[827:816]);
  assign MultLoop_acc_4410_nl = nl_MultLoop_acc_4410_nl[12:0];
  assign nl_MultLoop_acc_3159_nl = ({(data_rsci_idat[827:810]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4410_nl)
      , (~ (data_rsci_idat[815:810]))});
  assign MultLoop_acc_3159_nl = nl_MultLoop_acc_3159_nl[19:0];
  assign nl_MultLoop_acc_4411_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_3159_nl)))
      + (~ (data_rsci_idat[827:810]));
  assign MultLoop_acc_4411_nl = nl_MultLoop_acc_4411_nl[17:0];
  assign nl_MultLoop_acc_4681_nl = conv_s2u_19_21(MultLoop_acc_1715_itm_20_2_1) +
      ({(data_rsci_idat[485:468]) , 3'b001});
  assign MultLoop_acc_4681_nl = nl_MultLoop_acc_4681_nl[20:0];
  assign nl_MultLoop_acc_3171_nl = conv_s2s_20_21({(~ (data_rsci_idat[197:180]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_3171_nl = nl_MultLoop_acc_3171_nl[20:0];
  assign nl_MultLoop_acc_299_nl = conv_s2s_21_25(MultLoop_acc_3171_nl) + ({(data_rsci_idat[197:180])
      , 7'b0000100});
  assign MultLoop_acc_299_nl = nl_MultLoop_acc_299_nl[24:0];
  assign nl_MultLoop_acc_3256_itm_1  = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1194_nl)))
      + conv_s2s_15_18(readslicef_22_15_7((MultLoop_acc_290_nl))) + conv_s2s_14_18(readslicef_18_14_4((MultLoop_acc_4411_nl)))
      + conv_s2s_15_18(readslicef_21_15_6((MultLoop_acc_4681_nl))) + conv_s2s_15_18(MultLoop_acc_1476_itm_18_2[16:2])
      + conv_s2s_15_18(MultLoop_acc_307_itm_21_7) + conv_s2s_15_18(readslicef_25_15_10((MultLoop_acc_299_nl)));
  assign nl_MultLoop_acc_3175_nl = ({(data_rsci_idat[791:774]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[791:774]));
  assign MultLoop_acc_3175_nl = nl_MultLoop_acc_3175_nl[21:0];
  assign nl_MultLoop_acc_330_nl = conv_s2s_22_25(MultLoop_acc_3175_nl) + conv_s2s_24_25({(data_rsci_idat[791:774])
      , 6'b000000});
  assign MultLoop_acc_330_nl = nl_MultLoop_acc_330_nl[24:0];
  assign nl_MultLoop_acc_3176_nl = conv_s2s_20_21({(~ (data_rsci_idat[809:792]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[809:792]));
  assign MultLoop_acc_3176_nl = nl_MultLoop_acc_3176_nl[20:0];
  assign nl_MultLoop_acc_331_nl = conv_s2s_21_26(MultLoop_acc_3176_nl) + ({(data_rsci_idat[809:792])
      , 8'b00000100});
  assign MultLoop_acc_331_nl = nl_MultLoop_acc_331_nl[25:0];
  assign nl_MultLoop_acc_325_nl = conv_s2s_25_26({(~ (data_rsci_idat[701:684])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[701:684])) , 5'b00100}) +
      conv_s2s_20_26({(~ (data_rsci_idat[701:684])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_828_18_7
      , (~ (data_rsci_idat[690:684]))});
  assign MultLoop_acc_325_nl = nl_MultLoop_acc_325_nl[25:0];
  assign nl_MultLoop_acc_4644_nl = conv_s2u_15_19(MultLoop_acc_2073_cse_1[18:4])
      + conv_s2u_18_19(data_rsci_idat[665:648]);
  assign MultLoop_acc_4644_nl = nl_MultLoop_acc_4644_nl[18:0];
  assign nl_MultLoop_acc_3255_itm_1  = conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_330_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_331_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_325_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4644_nl)));
  assign nl_MultLoop_acc_3183_nl = ({(~ (data_rsci_idat[611:594])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3182_cse_1);
  assign MultLoop_acc_3183_nl = nl_MultLoop_acc_3183_nl[21:0];
  assign nl_MultLoop_acc_1189_nl = conv_s2u_22_24(MultLoop_acc_3183_nl) + ({(data_rsci_idat[611:594])
      , 6'b010000});
  assign MultLoop_acc_1189_nl = nl_MultLoop_acc_1189_nl[23:0];
  assign nl_MultLoop_acc_3184_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_16_18(data_rsci_idat[575:560]);
  assign MultLoop_acc_3184_nl = nl_MultLoop_acc_3184_nl[17:0];
  assign nl_MultLoop_acc_3185_nl = conv_s2s_20_21({(~ (data_rsci_idat[575:558]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3184_nl);
  assign MultLoop_acc_3185_nl = nl_MultLoop_acc_3185_nl[20:0];
  assign nl_MultLoop_acc_1187_nl = conv_s2u_21_23(MultLoop_acc_3185_nl) + ({(data_rsci_idat[575:558])
      , 5'b00100});
  assign MultLoop_acc_1187_nl = nl_MultLoop_acc_1187_nl[22:0];
  assign nl_MultLoop_acc_1188_nl = conv_s2u_18_22(Result_acc_152_cse_1) + ({(data_rsci_idat[593:576])
      , 4'b0001});
  assign MultLoop_acc_1188_nl = nl_MultLoop_acc_1188_nl[21:0];
  assign nl_MultLoop_acc_3188_nl = ({(~ (data_rsci_idat[467:450])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_3187_cse_1);
  assign MultLoop_acc_3188_nl = nl_MultLoop_acc_3188_nl[19:0];
  assign nl_MultLoop_acc_1185_nl = conv_s2u_20_24(MultLoop_acc_3188_nl) + ({(data_rsci_idat[467:450])
      , 6'b000100});
  assign MultLoop_acc_1185_nl = nl_MultLoop_acc_1185_nl[23:0];
  assign nl_MultLoop_acc_3254_itm_1  = conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1189_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1187_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1188_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1185_nl)));
  assign nl_MultLoop_acc_4682_nl = conv_s2u_16_19(MultLoop_acc_3190_itm_19_4) + conv_s2u_18_19(data_rsci_idat[395:378]);
  assign MultLoop_acc_4682_nl = nl_MultLoop_acc_4682_nl[18:0];
  assign nl_MultLoop_acc_4683_nl = conv_s2u_15_19(MultLoop_acc_3062_itm_19_4[15:1])
      + conv_s2u_18_19(data_rsci_idat[341:324]);
  assign MultLoop_acc_4683_nl = nl_MultLoop_acc_4683_nl[18:0];
  assign nl_MultLoop_acc_3238_itm_1  = conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4682_nl)))
      + conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4683_nl)));
  assign nl_MultLoop_acc_3194_nl = conv_s2s_23_24({(~ (data_rsci_idat[305:288]))
      , 5'b00100}) + conv_s2s_21_24(MultLoop_acc_1480_cse_1);
  assign MultLoop_acc_3194_nl = nl_MultLoop_acc_3194_nl[23:0];
  assign nl_MultLoop_acc_304_nl = conv_s2s_24_26(MultLoop_acc_3194_nl) + ({(data_rsci_idat[305:288])
      , 8'b00100000});
  assign MultLoop_acc_304_nl = nl_MultLoop_acc_304_nl[25:0];
  assign nl_MultLoop_acc_3198_nl = conv_s2s_22_23({(data_rsci_idat[323:306]) , 4'b0000})
      + conv_s2s_20_23({(data_rsci_idat[323:306]) , 2'b00}) + conv_s2s_18_23(data_rsci_idat[323:306])
      + conv_s2s_17_23({MultLoop_MultLoop_conc_778_16_6 , (data_rsci_idat[313:308])});
  assign MultLoop_acc_3198_nl = nl_MultLoop_acc_3198_nl[22:0];
  assign nl_MultLoop_acc_4414_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3198_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_4414_nl = nl_MultLoop_acc_4414_nl[17:0];
  assign nl_MultLoop_acc_3237_itm_1  = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_304_nl)))
      + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4414_nl)));
  assign nl_MultLoop_acc_760_nl = conv_s2s_18_23(~ (data_rsci_idat[35:18])) + ({(data_rsci_idat[35:18])
      , 5'b00001});
  assign MultLoop_acc_760_nl = nl_MultLoop_acc_760_nl[22:0];
  assign nl_MultLoop_acc_2262_nl = conv_s2s_13_14(readslicef_23_13_10((MultLoop_acc_760_nl)))
      + 14'b00001011011001;
  assign MultLoop_acc_2262_nl = nl_MultLoop_acc_2262_nl[13:0];
  assign nl_MultLoop_acc_2261_nl = ({(~ (data_rsci_idat[17:0])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_1043_cse_1);
  assign MultLoop_acc_2261_nl = nl_MultLoop_acc_2261_nl[21:0];
  assign nl_MultLoop_acc_759_nl = conv_s2s_22_24(MultLoop_acc_2261_nl) + ({(data_rsci_idat[17:0])
      , 6'b010000});
  assign MultLoop_acc_759_nl = nl_MultLoop_acc_759_nl[23:0];
  assign nl_MultLoop_770_MultLoop_acc_3_nl = conv_s2s_14_16(MultLoop_acc_2262_nl)
      + (readslicef_24_16_8((MultLoop_acc_759_nl)));
  assign MultLoop_770_MultLoop_acc_3_nl = nl_MultLoop_770_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_762_nl = conv_s2s_25_26({(~ (data_rsci_idat[71:54])) , 7'b0010000})
      + conv_s2s_22_26({(~ (data_rsci_idat[71:54])) , 4'b0001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_786_18_7
      , (~ (data_rsci_idat[60:54]))});
  assign MultLoop_acc_762_nl = nl_MultLoop_acc_762_nl[25:0];
  assign nl_MultLoop_acc_1327_nl = conv_s2u_18_21(MultLoop_acc_2259_cse_1) + ({(data_rsci_idat[53:36])
      , 3'b001});
  assign MultLoop_acc_1327_nl = nl_MultLoop_acc_1327_nl[20:0];
  assign nl_MultLoop_772_MultLoop_acc_3_nl = conv_s2s_16_17(MultLoop_770_MultLoop_acc_3_nl)
      + conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_762_nl))) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1327_nl)));
  assign MultLoop_772_MultLoop_acc_3_nl = nl_MultLoop_772_MultLoop_acc_3_nl[16:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_131_itm_1 
      = conv_s2s_17_18(MultLoop_acc_1237_itm_20_4) + conv_s2s_17_18(MultLoop_772_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_2267_nl = ({(data_rsci_idat[89:72]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_804_18_7
      , (~ (data_rsci_idat[78:72]))});
  assign MultLoop_acc_2267_nl = nl_MultLoop_acc_2267_nl[19:0];
  assign nl_MultLoop_acc_2268_nl = ({(~ (data_rsci_idat[89:72])) , 5'b00000}) + conv_s2s_20_23(MultLoop_acc_2267_nl);
  assign MultLoop_acc_2268_nl = nl_MultLoop_acc_2268_nl[22:0];
  assign nl_MultLoop_acc_763_nl = conv_s2s_23_26(MultLoop_acc_2268_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[89:72])) , 7'b0100000});
  assign MultLoop_acc_763_nl = nl_MultLoop_acc_763_nl[25:0];
  assign nl_MultLoop_acc_4093_nl =  -conv_s2s_14_15(data_rsci_idat[413:400]);
  assign MultLoop_acc_4093_nl = nl_MultLoop_acc_4093_nl[14:0];
  assign nl_MultLoop_acc_2192_nl = ({(data_rsci_idat[413:396]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4093_nl)
      , (~ (data_rsci_idat[399:396]))});
  assign MultLoop_acc_2192_nl = nl_MultLoop_acc_2192_nl[19:0];
  assign nl_MultLoop_acc_780_nl = conv_s2s_20_22(MultLoop_acc_2192_nl) + ({(~ (data_rsci_idat[413:396]))
      , 4'b0000});
  assign MultLoop_acc_780_nl = nl_MultLoop_acc_780_nl[21:0];
  assign nl_MultLoop_acc_4092_nl =  -conv_s2s_16_17(data_rsci_idat[233:218]);
  assign MultLoop_acc_4092_nl = nl_MultLoop_acc_4092_nl[16:0];
  assign nl_MultLoop_acc_770_nl = conv_s2s_19_21({(MultLoop_acc_4092_nl) , (~ (data_rsci_idat[217:216]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[233:216])) , 2'b01});
  assign MultLoop_acc_770_nl = nl_MultLoop_acc_770_nl[20:0];
  assign nl_MultLoop_acc_1330_nl = conv_s2u_16_19(data_rsci_idat[197:182]) + conv_s2u_18_19(data_rsci_idat[197:180]);
  assign MultLoop_acc_1330_nl = nl_MultLoop_acc_1330_nl[18:0];
  assign nl_MultLoop_acc_779_nl = conv_s2u_13_18(data_rsci_idat[395:383]) - (data_rsci_idat[395:378]);
  assign MultLoop_acc_779_nl = nl_MultLoop_acc_779_nl[17:0];
  assign nl_MultLoop_acc_4617_nl = conv_s2u_17_19(Result_acc_111_cse_1[18:2]) + conv_s2u_18_19(data_rsci_idat[107:90]);
  assign MultLoop_acc_4617_nl = nl_MultLoop_acc_4617_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_130_itm_1_16_0
      = (readslicef_26_17_9((MultLoop_acc_763_nl))) + conv_s2s_14_17(readslicef_22_14_8((MultLoop_acc_780_nl)))
      + conv_s2s_13_17(readslicef_21_13_8((MultLoop_acc_770_nl))) + conv_s2s_13_17(readslicef_19_13_6((MultLoop_acc_1330_nl)))
      + conv_s2s_14_17(readslicef_18_14_4((MultLoop_acc_779_nl))) + conv_s2s_14_17(readslicef_19_14_5((MultLoop_acc_4617_nl)));
  assign nl_MultLoop_acc_2194_nl = conv_s2s_18_19(data_rsci_idat[827:810]) + conv_s2s_15_19(data_rsci_idat[827:813]);
  assign MultLoop_acc_2194_nl = nl_MultLoop_acc_2194_nl[18:0];
  assign nl_MultLoop_acc_1344_nl = conv_s2u_19_22(MultLoop_acc_2194_nl) + conv_s2u_21_22({(data_rsci_idat[827:810])
      , 3'b000});
  assign MultLoop_acc_1344_nl = nl_MultLoop_acc_1344_nl[21:0];
  assign nl_MultLoop_acc_792_nl = conv_s2u_12_18(data_rsci_idat[629:618]) - (data_rsci_idat[629:612]);
  assign MultLoop_acc_792_nl = nl_MultLoop_acc_792_nl[17:0];
  assign nl_MultLoop_acc_2196_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_17_18({MultLoop_acc_4094_cse_1
      , (data_rsci_idat[562:560])});
  assign MultLoop_acc_2196_nl = nl_MultLoop_acc_2196_nl[17:0];
  assign nl_MultLoop_acc_1338_nl = conv_s2u_18_22(MultLoop_acc_2196_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[575:558])) , 3'b001});
  assign MultLoop_acc_1338_nl = nl_MultLoop_acc_1338_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_129_itm_1 
      = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1344_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_792_nl)))
      + conv_s2s_15_17(MultLoop_acc_788_cse_1[19:5]) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1338_nl)));
  assign nl_MultLoop_acc_4095_nl =  -conv_s2s_13_14(data_rsci_idat[467:455]);
  assign MultLoop_acc_4095_nl = nl_MultLoop_acc_4095_nl[13:0];
  assign nl_MultLoop_acc_783_nl = conv_s2s_23_24({(~ (data_rsci_idat[467:450])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[467:450])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4095_nl)
      , (~ (data_rsci_idat[454:450]))});
  assign MultLoop_acc_783_nl = nl_MultLoop_acc_783_nl[23:0];
  assign nl_MultLoop_acc_2199_nl = ({(data_rsci_idat[431:414]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[431:414]));
  assign MultLoop_acc_2199_nl = nl_MultLoop_acc_2199_nl[20:0];
  assign nl_MultLoop_acc_781_nl = conv_s2s_21_25(MultLoop_acc_2199_nl) + conv_s2s_24_25({(data_rsci_idat[431:414])
      , 6'b000000});
  assign MultLoop_acc_781_nl = nl_MultLoop_acc_781_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_128_itm_1 
      = conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_783_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_781_nl)))
      + conv_s2s_15_17(MultLoop_acc_67_itm_17_3) + conv_s2s_15_17(MultLoop_acc_355_itm_20_6);
  assign nl_MultLoop_acc_2206_nl = ({(data_rsci_idat[863:846]) , 6'b010000}) + conv_s2s_22_24({(~
      (data_rsci_idat[863:846])) , 4'b0001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_728_18_8
      , (~ (data_rsci_idat[853:846]))});
  assign MultLoop_acc_2206_nl = nl_MultLoop_acc_2206_nl[23:0];
  assign nl_MultLoop_acc_4098_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_2206_nl)))
      + (~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_4098_nl = nl_MultLoop_acc_4098_nl[17:0];
  assign nl_MultLoop_acc_2201_nl = (~ (data_rsci_idat[287:270])) + conv_s2s_17_18({MultLoop_acc_4075_cse_1
      , (data_rsci_idat[275:272])});
  assign MultLoop_acc_2201_nl = nl_MultLoop_acc_2201_nl[17:0];
  assign nl_MultLoop_acc_2202_nl = conv_s2s_20_21({(~ (data_rsci_idat[287:270]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2201_nl);
  assign MultLoop_acc_2202_nl = nl_MultLoop_acc_2202_nl[20:0];
  assign nl_MultLoop_acc_1334_nl = conv_s2u_21_23(MultLoop_acc_2202_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[287:270])) , 4'b0100});
  assign MultLoop_acc_1334_nl = nl_MultLoop_acc_1334_nl[22:0];
  assign nl_MultLoop_acc_2203_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_16_18(data_rsci_idat[251:236]);
  assign MultLoop_acc_2203_nl = nl_MultLoop_acc_2203_nl[17:0];
  assign nl_MultLoop_acc_1332_nl = conv_s2u_18_22(MultLoop_acc_2203_nl) + ({(data_rsci_idat[251:234])
      , 4'b0001});
  assign MultLoop_acc_1332_nl = nl_MultLoop_acc_1332_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_127_itm_1 
      = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4098_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1334_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1332_nl)));
  assign nl_MultLoop_acc_2208_nl = ({(data_rsci_idat[809:792]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_690_18_6
      , (~ (data_rsci_idat[797:792]))});
  assign MultLoop_acc_2208_nl = nl_MultLoop_acc_2208_nl[19:0];
  assign nl_MultLoop_acc_2209_nl = ({(~ (data_rsci_idat[809:792])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2208_nl);
  assign MultLoop_acc_2209_nl = nl_MultLoop_acc_2209_nl[21:0];
  assign nl_MultLoop_acc_802_nl = conv_s2s_22_25(MultLoop_acc_2209_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[809:792])) , 6'b010000});
  assign MultLoop_acc_802_nl = nl_MultLoop_acc_802_nl[24:0];
  assign nl_MultLoop_acc_2212_nl = conv_s2s_20_21({(data_rsci_idat[791:774]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[791:774]) + conv_s2s_17_21({MultLoop_MultLoop_conc_740_16_4
      , (data_rsci_idat[779:776])});
  assign MultLoop_acc_2212_nl = nl_MultLoop_acc_2212_nl[20:0];
  assign nl_MultLoop_acc_801_nl = conv_s2u_21_22(MultLoop_acc_2212_nl) + ({(~ (data_rsci_idat[791:774]))
      , 4'b0000});
  assign MultLoop_acc_801_nl = nl_MultLoop_acc_801_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_126_itm_1 
      = conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_802_nl))) + conv_s2s_16_17(readslicef_22_16_6((MultLoop_acc_801_nl)));
  assign nl_MultLoop_acc_798_nl = conv_s2s_24_25({(~ (data_rsci_idat[737:720])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[737:720])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[737:720])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_830_18_6
      , (~ (data_rsci_idat[725:720]))});
  assign MultLoop_acc_798_nl = nl_MultLoop_acc_798_nl[24:0];
  assign nl_MultLoop_acc_2216_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_13_18(data_rsci_idat[755:743]);
  assign MultLoop_acc_2216_nl = nl_MultLoop_acc_2216_nl[17:0];
  assign nl_MultLoop_acc_1343_nl = conv_s2u_18_20(MultLoop_acc_2216_nl) + ({(data_rsci_idat[755:738])
      , 2'b01});
  assign MultLoop_acc_1343_nl = nl_MultLoop_acc_1343_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_125_itm_1 
      = conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_798_nl))) + conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_1343_nl)));
  assign nl_MultLoop_acc_2218_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_15_18({Result_acc_183_cse_1
      , (data_rsci_idat[690:688])});
  assign MultLoop_acc_2218_nl = nl_MultLoop_acc_2218_nl[17:0];
  assign nl_MultLoop_acc_1341_nl = conv_s2u_18_22(MultLoop_acc_2218_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[701:684])) , 3'b001});
  assign MultLoop_acc_1341_nl = nl_MultLoop_acc_1341_nl[21:0];
  assign nl_MultLoop_acc_2221_nl = ({(~ (data_rsci_idat[719:702])) , 3'b000}) + conv_s2s_19_21(MultLoop_acc_2220_cse_1);
  assign MultLoop_acc_2221_nl = nl_MultLoop_acc_2221_nl[20:0];
  assign nl_MultLoop_acc_1342_nl = conv_s2u_21_24(MultLoop_acc_2221_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[719:702])) , 5'b01000});
  assign MultLoop_acc_1342_nl = nl_MultLoop_acc_1342_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_124_itm_1 
      = conv_s2s_16_17(readslicef_22_16_6((MultLoop_acc_1341_nl))) + conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_1342_nl)));
  assign nl_MultLoop_acc_2224_nl = ({(data_rsci_idat[665:648]) , 6'b000100}) + conv_s2s_20_24({(~
      (data_rsci_idat[665:648])) , 2'b01}) + conv_s2s_19_24({MultLoop_MultLoop_conc_756_18_8
      , (~ (data_rsci_idat[655:648]))});
  assign MultLoop_acc_2224_nl = nl_MultLoop_acc_2224_nl[23:0];
  assign nl_MultLoop_acc_4105_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_2224_nl)))
      + (~ (data_rsci_idat[665:648]));
  assign MultLoop_acc_4105_nl = nl_MultLoop_acc_4105_nl[17:0];
  assign nl_MultLoop_acc_2227_nl = ({(data_rsci_idat[593:576]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[593:576])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_704_18_6
      , (~ (data_rsci_idat[581:576]))});
  assign MultLoop_acc_2227_nl = nl_MultLoop_acc_2227_nl[21:0];
  assign nl_MultLoop_acc_4107_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2227_nl)))
      + (~ (data_rsci_idat[593:576]));
  assign MultLoop_acc_4107_nl = nl_MultLoop_acc_4107_nl[17:0];
  assign nl_MultLoop_acc_4108_nl =  -conv_s2s_12_13(data_rsci_idat[611:600]);
  assign MultLoop_acc_4108_nl = nl_MultLoop_acc_4108_nl[12:0];
  assign nl_MultLoop_acc_2230_nl = ({(data_rsci_idat[611:594]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[611:594])) , 2'b01}) + conv_s2s_19_22({(MultLoop_acc_4108_nl)
      , (~ (data_rsci_idat[599:594]))});
  assign MultLoop_acc_2230_nl = nl_MultLoop_acc_2230_nl[21:0];
  assign nl_MultLoop_acc_4109_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2230_nl)))
      + (~ (data_rsci_idat[611:594]));
  assign MultLoop_acc_4109_nl = nl_MultLoop_acc_4109_nl[17:0];
  assign nl_MultLoop_acc_2232_nl = (~ (data_rsci_idat[539:522])) + conv_s2s_15_18({MultLoop_MultLoop_conc_732_14_2
      , (data_rsci_idat[527:526])});
  assign MultLoop_acc_2232_nl = nl_MultLoop_acc_2232_nl[17:0];
  assign nl_MultLoop_acc_1337_nl = conv_s2u_18_21(MultLoop_acc_2232_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[539:522])) , 2'b01});
  assign MultLoop_acc_1337_nl = nl_MultLoop_acc_1337_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_135_itm_1 
      = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4105_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4107_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4109_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1337_nl)));
  assign nl_MultLoop_acc_4618_nl = conv_s2u_16_19(MultLoop_acc_4663_itm_19_4) + conv_s2u_18_19(data_rsci_idat[485:468]);
  assign MultLoop_acc_4618_nl = nl_MultLoop_acc_4618_nl[18:0];
  assign nl_MultLoop_acc_4111_nl =  -conv_s2s_10_11(data_rsci_idat[449:440]);
  assign MultLoop_acc_4111_nl = nl_MultLoop_acc_4111_nl[10:0];
  assign nl_MultLoop_acc_2237_nl = ({(data_rsci_idat[449:432]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[449:432])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_4111_nl)
      , (~ (data_rsci_idat[439:432]))});
  assign MultLoop_acc_2237_nl = nl_MultLoop_acc_2237_nl[22:0];
  assign nl_MultLoop_acc_4112_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_2237_nl)))
      + (~ (data_rsci_idat[449:432]));
  assign MultLoop_acc_4112_nl = nl_MultLoop_acc_4112_nl[17:0];
  assign nl_MultLoop_acc_4113_nl =  -conv_s2s_10_11(data_rsci_idat[377:368]);
  assign MultLoop_acc_4113_nl = nl_MultLoop_acc_4113_nl[10:0];
  assign nl_MultLoop_acc_2239_nl = ({(data_rsci_idat[377:360]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_4113_nl)
      , (~ (data_rsci_idat[367:360]))});
  assign MultLoop_acc_2239_nl = nl_MultLoop_acc_2239_nl[21:0];
  assign nl_MultLoop_acc_2240_nl = conv_s2s_24_25({(data_rsci_idat[377:360]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_2239_nl);
  assign MultLoop_acc_2240_nl = nl_MultLoop_acc_2240_nl[24:0];
  assign nl_MultLoop_acc_4114_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_2240_nl)))
      + (~ (data_rsci_idat[377:360]));
  assign MultLoop_acc_4114_nl = nl_MultLoop_acc_4114_nl[17:0];
  assign nl_MultLoop_acc_2243_nl = conv_s2s_24_25({(~ (data_rsci_idat[305:288]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[305:288])) , 4'b0100}) +
      conv_s2s_21_25(MultLoop_acc_1480_cse_1);
  assign MultLoop_acc_2243_nl = nl_MultLoop_acc_2243_nl[24:0];
  assign nl_MultLoop_acc_774_nl = conv_s2s_25_26(MultLoop_acc_2243_nl) + ({(data_rsci_idat[305:288])
      , 8'b01000000});
  assign MultLoop_acc_774_nl = nl_MultLoop_acc_774_nl[25:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_134_itm_1 
      = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4618_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4112_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4114_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_774_nl)));
  assign nl_MultLoop_acc_2258_nl = ({(~ (data_rsci_idat[683:666])) , 4'b0000}) +
      conv_s2s_18_22(data_rsci_idat[683:666]) + conv_s2s_17_22({MultLoop_MultLoop_conc_784_16_6
      , (data_rsci_idat[673:668])});
  assign MultLoop_acc_2258_nl = nl_MultLoop_acc_2258_nl[21:0];
  assign nl_MultLoop_acc_1340_nl = conv_s2u_22_25(MultLoop_acc_2258_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[683:666])) , 6'b010000});
  assign MultLoop_acc_1340_nl = nl_MultLoop_acc_1340_nl[24:0];
  assign nl_MultLoop_acc_2254_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_16_18(data_rsci_idat[143:128]);
  assign MultLoop_acc_2254_nl = nl_MultLoop_acc_2254_nl[17:0];
  assign nl_MultLoop_acc_2255_nl = ({(data_rsci_idat[143:126]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_2254_nl);
  assign MultLoop_acc_2255_nl = nl_MultLoop_acc_2255_nl[20:0];
  assign nl_MultLoop_acc_1329_nl = conv_s2u_21_24(MultLoop_acc_2255_nl) + conv_s2u_23_24({(data_rsci_idat[143:126])
      , 5'b00000});
  assign MultLoop_acc_1329_nl = nl_MultLoop_acc_1329_nl[23:0];
  assign nl_MultLoop_acc_2244_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_16_18(data_rsci_idat[323:308]);
  assign MultLoop_acc_2244_nl = nl_MultLoop_acc_2244_nl[17:0];
  assign nl_MultLoop_acc_2246_nl = conv_s2s_22_23({(~ (data_rsci_idat[323:306]))
      , 4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[323:306])) , 2'b01}) + conv_s2s_18_23(MultLoop_acc_2244_nl);
  assign MultLoop_acc_2246_nl = nl_MultLoop_acc_2246_nl[22:0];
  assign nl_MultLoop_acc_1335_nl = conv_s2u_23_24(MultLoop_acc_2246_nl) + ({(data_rsci_idat[323:306])
      , 6'b010000});
  assign MultLoop_acc_1335_nl = nl_MultLoop_acc_1335_nl[23:0];
  assign nl_MultLoop_acc_4115_nl = conv_s2s_11_12(data_rsci_idat[269:259]) + 12'b000000000001;
  assign MultLoop_acc_4115_nl = nl_MultLoop_acc_4115_nl[11:0];
  assign nl_MultLoop_acc_2249_nl = ({(~ (data_rsci_idat[269:252])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[269:252])
      + conv_s2s_16_20({(MultLoop_acc_4115_nl) , (data_rsci_idat[258:255])});
  assign MultLoop_acc_2249_nl = nl_MultLoop_acc_2249_nl[19:0];
  assign nl_MultLoop_acc_1333_nl = conv_s2u_20_23(MultLoop_acc_2249_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[269:252])) , 4'b0100});
  assign MultLoop_acc_1333_nl = nl_MultLoop_acc_1333_nl[22:0];
  assign nl_MultLoop_acc_4116_nl = conv_s2s_11_12(data_rsci_idat[215:205]) + 12'b000000000001;
  assign MultLoop_acc_4116_nl = nl_MultLoop_acc_4116_nl[11:0];
  assign nl_MultLoop_acc_2251_nl = (~ (data_rsci_idat[215:198])) + conv_s2s_17_18({(MultLoop_acc_4116_nl)
      , (data_rsci_idat[204:200])});
  assign MultLoop_acc_2251_nl = nl_MultLoop_acc_2251_nl[17:0];
  assign nl_MultLoop_acc_1331_nl = conv_s2u_18_24(MultLoop_acc_2251_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[215:198])) , 5'b00001});
  assign MultLoop_acc_1331_nl = nl_MultLoop_acc_1331_nl[23:0];
  assign nl_MultLoop_acc_4117_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_15_18(MultLoop_acc_2252_itm_20_5[15:1]);
  assign MultLoop_acc_4117_nl = nl_MultLoop_acc_4117_nl[17:0];
  assign nl_MultLoop_acc_4118_nl = conv_s2u_18_20(MultLoop_acc_4117_nl) + ({(data_rsci_idat[125:108])
      , 2'b01});
  assign MultLoop_acc_4118_nl = nl_MultLoop_acc_4118_nl[19:0];
  assign nl_MultLoop_acc_1336_nl = conv_s2u_14_19(data_rsci_idat[521:508]) + conv_s2u_18_19(data_rsci_idat[521:504]);
  assign MultLoop_acc_1336_nl = nl_MultLoop_acc_1336_nl[18:0];
  assign nl_MultLoop_acc_767_nl = conv_s2u_15_18(data_rsci_idat[161:147]) - (data_rsci_idat[161:144]);
  assign MultLoop_acc_767_nl = nl_MultLoop_acc_767_nl[17:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_6_nl = ~((data_rsci_idat[170:162]!=9'b000000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl = conv_s2s_11_12(readslicef_18_11_7((MultLoop_acc_767_nl)))
      + conv_s2s_9_12(~ (data_rsci_idat[179:171])) + conv_u2s_1_12(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_6_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl[11:0];
  assign nl_MultLoop_acc_800_nl = conv_s2u_15_18(data_rsci_idat[773:759]) - (data_rsci_idat[773:756]);
  assign MultLoop_acc_800_nl = nl_MultLoop_acc_800_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_140_itm_1 
      = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1340_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1329_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1335_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1333_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1331_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_4118_nl)))
      + conv_s2s_13_18(data_rsci_idat[845:833]) + conv_s2s_13_18(readslicef_19_13_6((MultLoop_acc_1336_nl)))
      + conv_s2s_13_18(MultLoop_acc_785_itm_17_4[13:1]) + conv_s2s_12_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_103_nl)
      + conv_s2s_12_18(readslicef_18_12_6((MultLoop_acc_800_nl)));
  assign nl_MultLoop_acc_3096_nl = (~ (data_rsci_idat[665:648])) + conv_s2s_16_18(data_rsci_idat[665:650]);
  assign MultLoop_acc_3096_nl = nl_MultLoop_acc_3096_nl[17:0];
  assign nl_MultLoop_acc_3097_nl = conv_s2s_20_21({(~ (data_rsci_idat[665:648]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3096_nl);
  assign MultLoop_acc_3097_nl = nl_MultLoop_acc_3097_nl[20:0];
  assign nl_MultLoop_acc_1207_nl = conv_s2u_21_22(MultLoop_acc_3097_nl) + ({(data_rsci_idat[665:648])
      , 4'b0100});
  assign MultLoop_acc_1207_nl = nl_MultLoop_acc_1207_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_298_itm_1 
      = conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_1207_nl))) + conv_s2s_14_16(MultLoop_acc_1708_cse_1[18:5])
      + conv_s2s_14_16(MultLoop_acc_1204_itm_19_5[14:1]) + conv_s2s_14_16(MultLoop_acc_1200_itm_19_4[15:2]);
  assign nl_MultLoop_acc_4371_nl =  -conv_s2s_14_15(data_rsci_idat[377:364]);
  assign MultLoop_acc_4371_nl = nl_MultLoop_acc_4371_nl[14:0];
  assign nl_MultLoop_acc_356_nl = conv_s2s_19_23({(MultLoop_acc_4371_nl) , (~ (data_rsci_idat[363:360]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[377:360])) , 4'b0001});
  assign MultLoop_acc_356_nl = nl_MultLoop_acc_356_nl[22:0];
  assign nl_MultLoop_acc_4636_nl = conv_s2u_19_21(MultLoop_acc_3099_cse_1[21:3])
      + ({(data_rsci_idat[215:198]) , 3'b001});
  assign MultLoop_acc_4636_nl = nl_MultLoop_acc_4636_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_297_itm_1 
      = conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_356_nl))) + conv_s2s_14_16(MultLoop_acc_355_itm_20_6[14:1])
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_4636_nl))) + conv_s2s_13_16(MultLoop_acc_3283_cse[18:6]);
  assign nl_MultLoop_acc_3101_nl = ({(data_rsci_idat[845:828]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_696_18_7
      , (~ (data_rsci_idat[834:828]))});
  assign MultLoop_acc_3101_nl = nl_MultLoop_acc_3101_nl[21:0];
  assign nl_MultLoop_acc_4373_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_3101_nl)))
      + (~ (data_rsci_idat[845:828]));
  assign MultLoop_acc_4373_nl = nl_MultLoop_acc_4373_nl[17:0];
  assign nl_MultLoop_acc_1210_nl = conv_s2u_13_19(data_rsci_idat[863:851]) + conv_s2u_18_19(data_rsci_idat[863:846]);
  assign MultLoop_acc_1210_nl = nl_MultLoop_acc_1210_nl[18:0];
  assign nl_MultLoop_acc_4637_nl = conv_s2u_15_19(MultLoop_acc_2289_itm_20_5[15:1])
      + conv_s2u_18_19(data_rsci_idat[809:792]);
  assign MultLoop_acc_4637_nl = nl_MultLoop_acc_4637_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_311_itm_1 
      = conv_s2s_15_17(~ (data_rsci_idat[521:507])) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4373_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_1210_nl))) + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4637_nl)));
  assign nl_MultLoop_acc_4374_nl =  -conv_s2s_13_14(data_rsci_idat[755:743]);
  assign MultLoop_acc_4374_nl = nl_MultLoop_acc_4374_nl[13:0];
  assign nl_MultLoop_acc_3104_nl = ({(data_rsci_idat[755:738]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4374_nl)
      , (~ (data_rsci_idat[742:738]))});
  assign MultLoop_acc_3104_nl = nl_MultLoop_acc_3104_nl[20:0];
  assign nl_MultLoop_acc_376_nl = conv_s2s_21_23(MultLoop_acc_3104_nl) + ({(~ (data_rsci_idat[755:738]))
      , 5'b00000});
  assign MultLoop_acc_376_nl = nl_MultLoop_acc_376_nl[22:0];
  assign nl_MultLoop_acc_3106_nl = conv_s2s_20_21({(data_rsci_idat[485:468]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_3105_cse);
  assign MultLoop_acc_3106_nl = nl_MultLoop_acc_3106_nl[20:0];
  assign nl_MultLoop_acc_1201_nl = conv_s2u_21_23(MultLoop_acc_3106_nl) + conv_s2u_22_23({(data_rsci_idat[485:468])
      , 4'b0000});
  assign MultLoop_acc_1201_nl = nl_MultLoop_acc_1201_nl[22:0];
  assign nl_MultLoop_acc_4375_nl =  -conv_s2s_13_14(data_rsci_idat[413:401]);
  assign MultLoop_acc_4375_nl = nl_MultLoop_acc_4375_nl[13:0];
  assign nl_MultLoop_acc_3108_nl = ({(data_rsci_idat[413:396]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4375_nl)
      , (~ (data_rsci_idat[400:396]))});
  assign MultLoop_acc_3108_nl = nl_MultLoop_acc_3108_nl[20:0];
  assign nl_MultLoop_acc_358_nl = conv_s2s_21_23(MultLoop_acc_3108_nl) + ({(~ (data_rsci_idat[413:396]))
      , 5'b00000});
  assign MultLoop_acc_358_nl = nl_MultLoop_acc_358_nl[22:0];
  assign nl_MultLoop_acc_3109_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_16_18(data_rsci_idat[269:254]);
  assign MultLoop_acc_3109_nl = nl_MultLoop_acc_3109_nl[17:0];
  assign nl_MultLoop_acc_3110_nl = conv_s2s_20_21({(~ (data_rsci_idat[269:252]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_3109_nl);
  assign MultLoop_acc_3110_nl = nl_MultLoop_acc_3110_nl[20:0];
  assign nl_MultLoop_acc_1197_nl = conv_s2u_21_22(MultLoop_acc_3110_nl) + ({(data_rsci_idat[269:252])
      , 4'b0100});
  assign MultLoop_acc_1197_nl = nl_MultLoop_acc_1197_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_310_itm_1 
      = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_376_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1201_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_358_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1197_nl)));
  assign nl_MultLoop_acc_4376_nl =  -conv_s2s_15_16(data_rsci_idat[233:219]);
  assign MultLoop_acc_4376_nl = nl_MultLoop_acc_4376_nl[15:0];
  assign nl_MultLoop_acc_348_nl = conv_s2s_19_22({(MultLoop_acc_4376_nl) , (~ (data_rsci_idat[218:216]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[233:216])) , 3'b001});
  assign MultLoop_acc_348_nl = nl_MultLoop_acc_348_nl[21:0];
  assign nl_MultLoop_acc_3112_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_14_18(data_rsci_idat[107:94]);
  assign MultLoop_acc_3112_nl = nl_MultLoop_acc_3112_nl[17:0];
  assign nl_MultLoop_acc_1196_nl = conv_s2u_18_21(MultLoop_acc_3112_nl) + ({(data_rsci_idat[107:90])
      , 3'b001});
  assign MultLoop_acc_1196_nl = nl_MultLoop_acc_1196_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_309_itm_1 
      = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_348_nl))) + conv_s2s_15_17(MultLoop_acc_343_itm_19_5)
      + conv_s2s_15_17(MultLoop_acc_340_itm_17_3) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1196_nl)));
  assign nl_MultLoop_acc_4377_nl =  -conv_s2s_10_11(data_rsci_idat[791:782]);
  assign MultLoop_acc_4377_nl = nl_MultLoop_acc_4377_nl[10:0];
  assign nl_MultLoop_acc_3114_nl = ({(data_rsci_idat[791:774]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_4377_nl)
      , (~ (data_rsci_idat[781:774]))});
  assign MultLoop_acc_3114_nl = nl_MultLoop_acc_3114_nl[21:0];
  assign nl_MultLoop_acc_3115_nl = conv_s2s_24_25({(data_rsci_idat[791:774]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_3114_nl);
  assign MultLoop_acc_3115_nl = nl_MultLoop_acc_3115_nl[24:0];
  assign nl_MultLoop_acc_4378_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_3115_nl)))
      + (~ (data_rsci_idat[791:774]));
  assign MultLoop_acc_4378_nl = nl_MultLoop_acc_4378_nl[17:0];
  assign nl_MultLoop_acc_3119_nl = conv_s2s_22_23({(data_rsci_idat[719:702]) , 4'b0000})
      + conv_s2s_20_23({(data_rsci_idat[719:702]) , 2'b00}) + conv_s2s_18_23(data_rsci_idat[719:702])
      + conv_s2s_17_23({Result_acc_206_cse_1 , (data_rsci_idat[709:704])});
  assign MultLoop_acc_3119_nl = nl_MultLoop_acc_3119_nl[22:0];
  assign nl_MultLoop_acc_4380_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_3119_nl)))
      + (~ (data_rsci_idat[719:702]));
  assign MultLoop_acc_4380_nl = nl_MultLoop_acc_4380_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_308_itm_1 
      = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4378_nl))) + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4380_nl)));
  assign nl_MultLoop_acc_4381_nl =  -conv_s2s_10_11(data_rsci_idat[683:674]);
  assign MultLoop_acc_4381_nl = nl_MultLoop_acc_4381_nl[10:0];
  assign nl_MultLoop_acc_3121_nl = ({(data_rsci_idat[683:666]) , 4'b0001}) + conv_s2s_19_22({(MultLoop_acc_4381_nl)
      , (~ (data_rsci_idat[673:666]))});
  assign MultLoop_acc_3121_nl = nl_MultLoop_acc_3121_nl[21:0];
  assign nl_MultLoop_acc_3122_nl = conv_s2s_24_25({(data_rsci_idat[683:666]) , 6'b000000})
      + conv_s2s_22_25(MultLoop_acc_3121_nl);
  assign MultLoop_acc_3122_nl = nl_MultLoop_acc_3122_nl[24:0];
  assign nl_MultLoop_acc_4382_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_3122_nl)))
      + (~ (data_rsci_idat[683:666]));
  assign MultLoop_acc_4382_nl = nl_MultLoop_acc_4382_nl[17:0];
  assign nl_MultLoop_acc_3124_nl = conv_s2s_21_22({(data_rsci_idat[611:594]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[611:594]) + conv_s2s_16_22(data_rsci_idat[611:596]);
  assign MultLoop_acc_3124_nl = nl_MultLoop_acc_3124_nl[21:0];
  assign nl_MultLoop_acc_1205_nl = conv_s2u_22_24(MultLoop_acc_3124_nl) + conv_s2u_23_24({(data_rsci_idat[611:594])
      , 5'b00000});
  assign MultLoop_acc_1205_nl = nl_MultLoop_acc_1205_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_307_itm_1 
      = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4382_nl))) + conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_1205_nl)));
  assign nl_MultLoop_acc_3126_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_16_18({MultLoop_acc_4146_cse_1
      , (data_rsci_idat[547:543])});
  assign MultLoop_acc_3126_nl = nl_MultLoop_acc_3126_nl[17:0];
  assign nl_MultLoop_acc_3127_nl = ({(data_rsci_idat[557:540]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_3126_nl);
  assign MultLoop_acc_3127_nl = nl_MultLoop_acc_3127_nl[19:0];
  assign nl_MultLoop_acc_365_nl = conv_s2u_20_23(MultLoop_acc_3127_nl) + ({(~ (data_rsci_idat[557:540]))
      , 5'b00000});
  assign MultLoop_acc_365_nl = nl_MultLoop_acc_365_nl[22:0];
  assign nl_MultLoop_acc_366_nl = conv_s2s_18_25(~ (data_rsci_idat[575:558])) + ({(data_rsci_idat[575:558])
      , 7'b0000001});
  assign MultLoop_acc_366_nl = nl_MultLoop_acc_366_nl[24:0];
  assign nl_MultLoop_acc_3129_nl = ({(~ (data_rsci_idat[539:522])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_1962_cse_1);
  assign MultLoop_acc_3129_nl = nl_MultLoop_acc_3129_nl[19:0];
  assign nl_MultLoop_acc_1203_nl = conv_s2u_20_22(MultLoop_acc_3129_nl) + ({(data_rsci_idat[539:522])
      , 4'b0100});
  assign MultLoop_acc_1203_nl = nl_MultLoop_acc_1203_nl[21:0];
  assign nl_MultLoop_acc_3131_nl = conv_s2s_23_24({(~ (data_rsci_idat[449:432]))
      , 5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[449:432])) , 2'b01}) + conv_s2s_18_24(~
      (data_rsci_idat[449:432]));
  assign MultLoop_acc_3131_nl = nl_MultLoop_acc_3131_nl[23:0];
  assign nl_MultLoop_acc_360_nl = conv_s2s_24_25(MultLoop_acc_3131_nl) + ({(data_rsci_idat[449:432])
      , 7'b0100000});
  assign MultLoop_acc_360_nl = nl_MultLoop_acc_360_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_317_itm_1 
      = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_365_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_366_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1203_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_360_nl)));
  assign nl_MultLoop_acc_4384_nl =  -conv_s2s_14_15(data_rsci_idat[395:382]);
  assign MultLoop_acc_4384_nl = nl_MultLoop_acc_4384_nl[14:0];
  assign nl_MultLoop_acc_3133_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4384_nl)
      , (~ (data_rsci_idat[381:378]))});
  assign MultLoop_acc_3133_nl = nl_MultLoop_acc_3133_nl[19:0];
  assign nl_MultLoop_acc_357_nl = conv_s2s_20_22(MultLoop_acc_3133_nl) + ({(~ (data_rsci_idat[395:378]))
      , 4'b0000});
  assign MultLoop_acc_357_nl = nl_MultLoop_acc_357_nl[21:0];
  assign nl_MultLoop_acc_3135_nl = ({(data_rsci_idat[341:324]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_854_18_8
      , (~ (data_rsci_idat[331:324]))});
  assign MultLoop_acc_3135_nl = nl_MultLoop_acc_3135_nl[20:0];
  assign nl_MultLoop_acc_3136_nl = conv_s2s_23_24({(data_rsci_idat[341:324]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_3135_nl);
  assign MultLoop_acc_3136_nl = nl_MultLoop_acc_3136_nl[23:0];
  assign nl_MultLoop_acc_4386_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_3136_nl)))
      + (~ (data_rsci_idat[341:324]));
  assign MultLoop_acc_4386_nl = nl_MultLoop_acc_4386_nl[17:0];
  assign nl_MultLoop_acc_352_nl = conv_s2u_11_18(data_rsci_idat[305:295]) - (data_rsci_idat[305:288]);
  assign MultLoop_acc_352_nl = nl_MultLoop_acc_352_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_316_itm_1 
      = conv_s2s_16_18(MultLoop_acc_4587_itm_18_3) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_357_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4386_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_352_nl)));
  assign nl_MultLoop_acc_1198_nl = conv_s2u_14_19(data_rsci_idat[323:310]) + conv_s2u_18_19(data_rsci_idat[323:306]);
  assign MultLoop_acc_1198_nl = nl_MultLoop_acc_1198_nl[18:0];
  assign nl_MultLoop_acc_4638_nl = conv_s2u_14_19(MultLoop_acc_2836_itm_19_6) + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_4638_nl = nl_MultLoop_acc_4638_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_302_itm_1 
      = conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_1198_nl))) + conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4638_nl)));
  assign nl_MultLoop_acc_4387_nl =  -conv_s2s_11_12(data_rsci_idat[251:241]);
  assign MultLoop_acc_4387_nl = nl_MultLoop_acc_4387_nl[11:0];
  assign nl_MultLoop_acc_349_nl = conv_s2s_25_26({(~ (data_rsci_idat[251:234])) ,
      7'b0000100}) + conv_s2s_20_26({(~ (data_rsci_idat[251:234])) , 2'b01}) + conv_s2s_19_26({(MultLoop_acc_4387_nl)
      , (~ (data_rsci_idat[240:234]))});
  assign MultLoop_acc_349_nl = nl_MultLoop_acc_349_nl[25:0];
  assign nl_MultLoop_acc_346_nl = conv_s2s_25_26({(~ (data_rsci_idat[197:180])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[197:180])) , 5'b01000}) +
      conv_s2s_21_26({(~ (data_rsci_idat[197:180])) , 3'b001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_698_18_7
      , (~ (data_rsci_idat[186:180]))});
  assign MultLoop_acc_346_nl = nl_MultLoop_acc_346_nl[25:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_301_itm_1 
      = conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_349_nl))) + conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_346_nl)));
  assign nl_MultLoop_acc_3144_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_15_19({MultLoop_acc_4162_cse_1
      , (data_rsci_idat[150:148])});
  assign MultLoop_acc_3144_nl = nl_MultLoop_acc_3144_nl[18:0];
  assign nl_MultLoop_acc_344_nl = conv_s2u_19_21(MultLoop_acc_3144_nl) + ({(~ (data_rsci_idat[161:144]))
      , 3'b000});
  assign MultLoop_acc_344_nl = nl_MultLoop_acc_344_nl[20:0];
  assign nl_MultLoop_acc_342_nl = conv_s2s_25_26({(~ (data_rsci_idat[125:108])) ,
      7'b0000100}) + conv_s2s_20_26({(~ (data_rsci_idat[125:108])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_832_18_7
      , (~ (data_rsci_idat[114:108]))});
  assign MultLoop_acc_342_nl = nl_MultLoop_acc_342_nl[25:0];
  assign nl_MultLoop_acc_4392_nl = (MultLoop_acc_335_itm_21_9[12:1]) + 12'b000001110001;
  assign MultLoop_acc_4392_nl = nl_MultLoop_acc_4392_nl[11:0];
  assign nl_MultLoop_acc_4393_nl =  -conv_s2s_13_14(data_rsci_idat[35:23]);
  assign MultLoop_acc_4393_nl = nl_MultLoop_acc_4393_nl[13:0];
  assign nl_MultLoop_acc_337_nl = conv_s2s_19_24({(MultLoop_acc_4393_nl) , (~ (data_rsci_idat[22:18]))})
      + conv_s2s_23_24({(~ (data_rsci_idat[35:18])) , 5'b00001});
  assign MultLoop_acc_337_nl = nl_MultLoop_acc_337_nl[23:0];
  assign nl_MultLoop_338_MultLoop_acc_3_nl = conv_s2s_13_14({(MultLoop_acc_4392_nl)
      , (MultLoop_acc_335_itm_21_9[0])}) + (readslicef_24_14_10((MultLoop_acc_337_nl)));
  assign MultLoop_338_MultLoop_acc_3_nl = nl_MultLoop_338_MultLoop_acc_3_nl[13:0];
  assign nl_MultLoop_acc_3154_nl = conv_s2s_14_15(MultLoop_338_MultLoop_acc_3_nl)
      + conv_s2s_14_15(MultLoop_acc_4594_itm_18_2[16:3]);
  assign MultLoop_acc_3154_nl = nl_MultLoop_acc_3154_nl[14:0];
  assign nl_MultLoop_acc_3153_nl = conv_s2s_21_22({(~ (data_rsci_idat[71:54])) ,
      3'b001}) + conv_s2s_18_22(MultLoop_acc_1636_cse_1);
  assign MultLoop_acc_3153_nl = nl_MultLoop_acc_3153_nl[21:0];
  assign nl_MultLoop_acc_1195_nl = conv_s2u_22_24(MultLoop_acc_3153_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[71:54])) , 5'b01000});
  assign MultLoop_acc_1195_nl = nl_MultLoop_acc_1195_nl[23:0];
  assign nl_MultLoop_340_MultLoop_acc_3_nl = conv_s2s_15_16(MultLoop_acc_3154_nl)
      + (readslicef_24_16_8((MultLoop_acc_1195_nl)));
  assign MultLoop_340_MultLoop_acc_3_nl = nl_MultLoop_340_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_4395_nl = conv_s2s_14_15(data_rsci_idat[179:166]) + 15'b000000000000001;
  assign MultLoop_acc_4395_nl = nl_MultLoop_acc_4395_nl[14:0];
  assign nl_MultLoop_acc_3094_nl = conv_s2s_18_19(data_rsci_idat[179:162]) + conv_s2s_17_19({(MultLoop_acc_4395_nl)
      , (data_rsci_idat[165:164])});
  assign MultLoop_acc_3094_nl = nl_MultLoop_acc_3094_nl[18:0];
  assign nl_MultLoop_acc_345_nl = conv_s2u_19_20(MultLoop_acc_3094_nl) + ({(~ (data_rsci_idat[179:162]))
      , 2'b00});
  assign MultLoop_acc_345_nl = nl_MultLoop_acc_345_nl[19:0];
  assign nl_MultLoop_acc_4396_nl =  -conv_s2s_16_17(data_rsci_idat[647:632]);
  assign MultLoop_acc_4396_nl = nl_MultLoop_acc_4396_nl[16:0];
  assign nl_MultLoop_acc_370_nl = conv_s2s_19_21({(MultLoop_acc_4396_nl) , (~ (data_rsci_idat[631:630]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[647:630])) , 2'b01});
  assign MultLoop_acc_370_nl = nl_MultLoop_acc_370_nl[20:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl = ~((data_rsci_idat[818:810]!=9'b000000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl = (readslicef_21_12_9((MultLoop_acc_370_nl)))
      + conv_s2s_9_12(~ (data_rsci_idat[827:819])) + conv_u2s_1_12(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_2_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl[11:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl = ~((data_rsci_idat[506:504]!=3'b000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl = conv_s2s_13_14(readslicef_20_13_7((MultLoop_acc_345_nl)))
      + conv_s2s_12_14(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_284_nl)
      + conv_u2s_1_14(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_1_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl[13:0];
  assign nl_MultLoop_acc_3095_nl = (~ (data_rsci_idat[773:756])) + conv_s2s_15_18(data_rsci_idat[773:759]);
  assign MultLoop_acc_3095_nl = nl_MultLoop_acc_3095_nl[17:0];
  assign nl_MultLoop_acc_1209_nl = conv_s2u_18_21(MultLoop_acc_3095_nl) + ({(data_rsci_idat[773:756])
      , 3'b001});
  assign MultLoop_acc_1209_nl = nl_MultLoop_acc_1209_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_314_itm_1 
      = conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_344_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_342_nl)))
      + conv_s2s_16_18(MultLoop_340_MultLoop_acc_3_nl) + conv_s2s_14_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_285_nl)
      + conv_s2s_14_18(readslicef_21_14_7((MultLoop_acc_1209_nl)));
  assign nl_MultLoop_acc_375_nl = conv_s2s_19_27({MultLoop_MultLoop_conc_820_18_8
      , (~ (data_rsci_idat[727:720]))}) + conv_s2s_26_27({(~ (data_rsci_idat[737:720]))
      , 8'b00000001});
  assign MultLoop_acc_375_nl = nl_MultLoop_acc_375_nl[26:0];
  assign nl_MultLoop_acc_4398_nl = conv_s2s_10_11(data_rsci_idat[701:692]) + 11'b00000000001;
  assign MultLoop_acc_4398_nl = nl_MultLoop_acc_4398_nl[10:0];
  assign nl_MultLoop_acc_3157_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_14_18({(MultLoop_acc_4398_nl)
      , (data_rsci_idat[691:689])});
  assign MultLoop_acc_3157_nl = nl_MultLoop_acc_3157_nl[17:0];
  assign nl_MultLoop_acc_1208_nl = conv_s2u_18_22(MultLoop_acc_3157_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[701:684])) , 3'b001});
  assign MultLoop_acc_1208_nl = nl_MultLoop_acc_1208_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_313_itm_1 
      = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_375_nl))) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1208_nl)));
  assign nl_MultLoop_acc_2344_nl = ({(~ (data_rsci_idat[341:324])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[341:324])
      + conv_s2s_17_20({MultLoop_acc_4122_cse_1 , (data_rsci_idat[331:326])});
  assign MultLoop_acc_2344_nl = nl_MultLoop_acc_2344_nl[19:0];
  assign nl_MultLoop_acc_1319_nl = conv_s2u_20_25(MultLoop_acc_2344_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[341:324])) , 6'b000100});
  assign MultLoop_acc_1319_nl = nl_MultLoop_acc_1319_nl[24:0];
  assign nl_MultLoop_acc_4123_nl = conv_s2s_12_13(data_rsci_idat[323:312]) + 13'b0000000000001;
  assign MultLoop_acc_4123_nl = nl_MultLoop_acc_4123_nl[12:0];
  assign nl_MultLoop_acc_2346_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_16_18({(MultLoop_acc_4123_nl)
      , (data_rsci_idat[311:309])});
  assign MultLoop_acc_2346_nl = nl_MultLoop_acc_2346_nl[17:0];
  assign nl_MultLoop_acc_1318_nl = conv_s2u_18_22(MultLoop_acc_2346_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[323:306])) , 3'b001});
  assign MultLoop_acc_1318_nl = nl_MultLoop_acc_1318_nl[21:0];
  assign nl_MultLoop_acc_724_nl = conv_s2s_25_26({(~ (data_rsci_idat[233:216])) ,
      7'b0010000}) + conv_s2s_22_26({(~ (data_rsci_idat[233:216])) , 4'b0001}) +
      conv_s2s_19_26({MultLoop_MultLoop_conc_730_18_7 , (~ (data_rsci_idat[222:216]))});
  assign MultLoop_acc_724_nl = nl_MultLoop_acc_724_nl[25:0];
  assign nl_MultLoop_acc_712_nl = (MultLoop_acc_713_itm_23_8[15:2]) + 14'b00000000110111;
  assign MultLoop_acc_712_nl = nl_MultLoop_acc_712_nl[13:0];
  assign nl_MultLoop_acc_727_nl = conv_s2s_24_25({(~ (data_rsci_idat[287:270])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[287:270])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_752_18_6
      , (~ (data_rsci_idat[275:270]))});
  assign MultLoop_acc_727_nl = nl_MultLoop_acc_727_nl[24:0];
  assign nl_MultLoop_acc_748_nl = conv_s2s_22_23({(~ (data_rsci_idat[683:666])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[683:666])) , 2'b01}) + conv_s2s_19_23({MultLoop_MultLoop_conc_838_18_4
      , (~ (data_rsci_idat[669:666]))});
  assign MultLoop_acc_748_nl = nl_MultLoop_acc_748_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl = (readslicef_25_15_10((MultLoop_acc_727_nl)))
      + conv_s2s_13_15(readslicef_23_13_10((MultLoop_acc_748_nl))) + conv_s2s_13_15(MultLoop_acc_3105_cse[18:6]);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl[14:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_184_itm_1 
      = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1319_nl))) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1318_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_724_nl))) + conv_s2s_16_18({(MultLoop_acc_712_nl)
      , (MultLoop_acc_713_itm_23_8[1:0])}) + conv_s2s_15_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_153_nl);
  assign nl_MultLoop_acc_4125_nl =  -conv_s2s_10_11(data_rsci_idat[143:134]);
  assign MultLoop_acc_4125_nl = nl_MultLoop_acc_4125_nl[10:0];
  assign nl_MultLoop_acc_720_nl = conv_s2s_26_27({(~ (data_rsci_idat[143:126])) ,
      8'b00001000}) + conv_s2s_21_27({(~ (data_rsci_idat[143:126])) , 3'b001}) +
      conv_s2s_19_27({(MultLoop_acc_4125_nl) , (~ (data_rsci_idat[133:126]))});
  assign MultLoop_acc_720_nl = nl_MultLoop_acc_720_nl[26:0];
  assign nl_MultLoop_acc_716_nl = conv_s2s_18_21(~ (data_rsci_idat[71:54])) + ({(data_rsci_idat[71:54])
      , 3'b001});
  assign MultLoop_acc_716_nl = nl_MultLoop_acc_716_nl[20:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_5_nl = ~((data_rsci_idat[203:198]!=6'b000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl = conv_s2s_13_14(readslicef_21_13_8((MultLoop_acc_716_nl)))
      + conv_s2s_12_14(~ (data_rsci_idat[215:204])) + conv_u2s_1_14(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_5_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl[13:0];
  assign nl_MultLoop_acc_1326_nl = conv_s2u_18_21(MultLoop_acc_2035_cse_1) + ({(data_rsci_idat[791:774])
      , 3'b001});
  assign MultLoop_acc_1326_nl = nl_MultLoop_acc_1326_nl[20:0];
  assign nl_MultLoop_acc_4126_nl =  -conv_s2s_13_14(data_rsci_idat[737:725]);
  assign MultLoop_acc_4126_nl = nl_MultLoop_acc_4126_nl[13:0];
  assign nl_MultLoop_acc_751_nl = conv_s2s_23_24({(~ (data_rsci_idat[737:720])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[737:720])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4126_nl)
      , (~ (data_rsci_idat[724:720]))});
  assign MultLoop_acc_751_nl = nl_MultLoop_acc_751_nl[23:0];
  assign nl_MultLoop_acc_4127_nl = conv_s2s_12_13(data_rsci_idat[593:582]) + 13'b0000000000001;
  assign MultLoop_acc_4127_nl = nl_MultLoop_acc_4127_nl[12:0];
  assign nl_MultLoop_acc_2276_nl = (~ (data_rsci_idat[593:576])) + conv_s2s_17_18({(MultLoop_acc_4127_nl)
      , (data_rsci_idat[581:578])});
  assign MultLoop_acc_2276_nl = nl_MultLoop_acc_2276_nl[17:0];
  assign nl_MultLoop_acc_2277_nl = ({(data_rsci_idat[593:576]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2276_nl);
  assign MultLoop_acc_2277_nl = nl_MultLoop_acc_2277_nl[19:0];
  assign nl_MultLoop_acc_743_nl = conv_s2u_20_22(MultLoop_acc_2277_nl) + ({(~ (data_rsci_idat[593:576]))
      , 4'b0000});
  assign MultLoop_acc_743_nl = nl_MultLoop_acc_743_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_159_itm_1 
      = conv_s2s_14_16(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_146_nl)
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1326_nl))) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_751_nl)))
      + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_743_nl)));
  assign nl_MultLoop_acc_4128_nl =  -conv_s2s_16_17(data_rsci_idat[539:524]);
  assign MultLoop_acc_4128_nl = nl_MultLoop_acc_4128_nl[16:0];
  assign nl_MultLoop_acc_740_nl = conv_s2s_19_21({(MultLoop_acc_4128_nl) , (~ (data_rsci_idat[523:522]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[539:522])) , 2'b01});
  assign MultLoop_acc_740_nl = nl_MultLoop_acc_740_nl[20:0];
  assign nl_MultLoop_acc_4129_nl = conv_s2s_14_15(data_rsci_idat[413:400]) + 15'b000000000000001;
  assign MultLoop_acc_4129_nl = nl_MultLoop_acc_4129_nl[14:0];
  assign nl_MultLoop_acc_2280_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_17_19({(MultLoop_acc_4129_nl)
      , (data_rsci_idat[399:398])});
  assign MultLoop_acc_2280_nl = nl_MultLoop_acc_2280_nl[18:0];
  assign nl_MultLoop_acc_733_nl = conv_s2u_19_20(MultLoop_acc_2280_nl) + ({(~ (data_rsci_idat[413:396]))
      , 2'b00});
  assign MultLoop_acc_733_nl = nl_MultLoop_acc_733_nl[19:0];
  assign nl_MultLoop_acc_728_nl = conv_s2s_19_24({MultLoop_MultLoop_conc_674_18_5
      , (~ (data_rsci_idat[292:288]))}) + conv_s2s_23_24({(~ (data_rsci_idat[305:288]))
      , 5'b00001});
  assign MultLoop_acc_728_nl = nl_MultLoop_acc_728_nl[23:0];
  assign nl_MultLoop_acc_4669_nl = ({(data_rsci_idat[197:180]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_1816_itm_20_2_1);
  assign MultLoop_acc_4669_nl = nl_MultLoop_acc_4669_nl[19:0];
  assign nl_MultLoop_acc_4132_nl = conv_s2u_16_18(readslicef_20_16_4((MultLoop_acc_4669_nl)))
      + (~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_4132_nl = nl_MultLoop_acc_4132_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_158_itm_1 
      = conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_740_nl))) + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_733_nl)))
      + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_728_nl))) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4132_nl)));
  assign nl_MultLoop_acc_2287_nl = ({(data_rsci_idat[827:810]) , 2'b01}) + conv_s2s_19_20({MultLoop_acc_4133_itm
      , (~ (data_rsci_idat[816:810]))});
  assign MultLoop_acc_2287_nl = nl_MultLoop_acc_2287_nl[19:0];
  assign nl_MultLoop_acc_2288_nl = conv_s2s_22_23({(data_rsci_idat[827:810]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2287_nl);
  assign MultLoop_acc_2288_nl = nl_MultLoop_acc_2288_nl[22:0];
  assign nl_MultLoop_acc_4134_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_2288_nl)))
      + (~ (data_rsci_idat[827:810]));
  assign MultLoop_acc_4134_nl = nl_MultLoop_acc_4134_nl[17:0];
  assign nl_MultLoop_acc_2285_nl = conv_s2s_21_22({(~ (data_rsci_idat[125:108]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_2285_nl = nl_MultLoop_acc_2285_nl[21:0];
  assign nl_MultLoop_acc_719_nl = conv_s2s_22_24(MultLoop_acc_2285_nl) + ({(data_rsci_idat[125:108])
      , 6'b001000});
  assign MultLoop_acc_719_nl = nl_MultLoop_acc_719_nl[23:0];
  assign nl_MultLoop_acc_2269_nl = conv_s2s_20_21({(~ (data_rsci_idat[719:702]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[719:702]));
  assign MultLoop_acc_2269_nl = nl_MultLoop_acc_2269_nl[20:0];
  assign nl_MultLoop_acc_750_nl = conv_s2s_21_22(MultLoop_acc_2269_nl) + ({(data_rsci_idat[719:702])
      , 4'b0100});
  assign MultLoop_acc_750_nl = nl_MultLoop_acc_750_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_157_itm_1 
      = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4134_nl))) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_719_nl)))
      + conv_s2s_13_16(readslicef_22_13_9((MultLoop_acc_750_nl)));
  assign nl_MultLoop_acc_4619_nl = conv_s2u_16_19(MultLoop_acc_2289_itm_20_5) + conv_s2u_18_19(data_rsci_idat[809:792]);
  assign MultLoop_acc_4619_nl = nl_MultLoop_acc_4619_nl[18:0];
  assign nl_MultLoop_acc_2291_nl = ({(data_rsci_idat[611:594]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_750_18_7
      , (~ (data_rsci_idat[600:594]))});
  assign MultLoop_acc_2291_nl = nl_MultLoop_acc_2291_nl[19:0];
  assign nl_MultLoop_acc_2292_nl = conv_s2s_22_23({(data_rsci_idat[611:594]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2291_nl);
  assign MultLoop_acc_2292_nl = nl_MultLoop_acc_2292_nl[22:0];
  assign nl_MultLoop_acc_4136_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_2292_nl)))
      + (~ (data_rsci_idat[611:594]));
  assign MultLoop_acc_4136_nl = nl_MultLoop_acc_4136_nl[17:0];
  assign nl_MultLoop_acc_2294_nl = ({(~ (data_rsci_idat[575:558])) , 3'b000}) + conv_s2s_19_21(Result_acc_127_cse_1);
  assign MultLoop_acc_2294_nl = nl_MultLoop_acc_2294_nl[20:0];
  assign nl_MultLoop_acc_1323_nl = conv_s2u_21_23(MultLoop_acc_2294_nl) + ({(data_rsci_idat[575:558])
      , 5'b01000});
  assign MultLoop_acc_1323_nl = nl_MultLoop_acc_1323_nl[22:0];
  assign nl_MultLoop_acc_735_nl = conv_s2s_19_24({MultLoop_MultLoop_conc_806_18_5
      , (~ (data_rsci_idat[436:432]))}) + conv_s2s_23_24({(~ (data_rsci_idat[449:432]))
      , 5'b00001});
  assign MultLoop_acc_735_nl = nl_MultLoop_acc_735_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_172_itm_1 
      = conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4619_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4136_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1323_nl))) + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_735_nl)));
  assign nl_MultLoop_acc_4139_nl = conv_s2s_13_14(data_rsci_idat[845:833]) + 14'b00000000000001;
  assign MultLoop_acc_4139_nl = nl_MultLoop_acc_4139_nl[13:0];
  assign nl_MultLoop_acc_2303_nl = conv_s2s_18_19(data_rsci_idat[845:828]) + conv_s2s_16_19({(MultLoop_acc_4139_nl)
      , (data_rsci_idat[832:831])});
  assign MultLoop_acc_2303_nl = nl_MultLoop_acc_2303_nl[18:0];
  assign nl_MultLoop_acc_757_nl = conv_s2u_19_20(MultLoop_acc_2303_nl) + ({(~ (data_rsci_idat[845:828]))
      , 2'b00});
  assign MultLoop_acc_757_nl = nl_MultLoop_acc_757_nl[19:0];
  assign nl_MultLoop_acc_4138_nl = conv_s2s_13_14(data_rsci_idat[377:365]) + 14'b00000000000001;
  assign MultLoop_acc_4138_nl = nl_MultLoop_acc_4138_nl[13:0];
  assign nl_MultLoop_acc_2297_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_16_18({(MultLoop_acc_4138_nl)
      , (data_rsci_idat[364:363])});
  assign MultLoop_acc_2297_nl = nl_MultLoop_acc_2297_nl[17:0];
  assign nl_MultLoop_acc_1320_nl = conv_s2u_18_21(MultLoop_acc_2297_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[377:360])) , 2'b01});
  assign MultLoop_acc_1320_nl = nl_MultLoop_acc_1320_nl[20:0];
  assign nl_MultLoop_acc_2299_nl = conv_s2s_23_24({(~ (data_rsci_idat[359:342]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[359:342])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[359:342]));
  assign MultLoop_acc_2299_nl = nl_MultLoop_acc_2299_nl[23:0];
  assign nl_MultLoop_acc_731_nl = conv_s2s_24_25(MultLoop_acc_2299_nl) + ({(data_rsci_idat[359:342])
      , 7'b0100000});
  assign MultLoop_acc_731_nl = nl_MultLoop_acc_731_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_171_itm_1 
      = conv_s2s_16_17(readslicef_20_16_4((MultLoop_acc_757_nl))) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1320_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_731_nl)));
  assign nl_MultLoop_acc_2304_nl = ({(data_rsci_idat[863:846]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[863:846]));
  assign MultLoop_acc_2304_nl = nl_MultLoop_acc_2304_nl[20:0];
  assign nl_MultLoop_acc_4140_nl = conv_s2u_14_19(readslicef_21_14_7((MultLoop_acc_2304_nl)))
      + conv_s2u_18_19(data_rsci_idat[863:846]);
  assign MultLoop_acc_4140_nl = nl_MultLoop_acc_4140_nl[18:0];
  assign nl_MultLoop_acc_4620_nl = conv_s2u_14_18(Result_acc_163_cse_1[18:5]) + (~
      (data_rsci_idat[755:738]));
  assign MultLoop_acc_4620_nl = nl_MultLoop_acc_4620_nl[17:0];
  assign nl_MultLoop_acc_1325_nl = conv_s2u_18_20(MultLoop_acc_2307_cse_1) + ({(data_rsci_idat[773:756])
      , 2'b01});
  assign MultLoop_acc_1325_nl = nl_MultLoop_acc_1325_nl[19:0];
  assign nl_MultLoop_acc_2310_nl = ({(data_rsci_idat[701:684]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[701:684])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_782_18_8
      , (~ (data_rsci_idat[691:684]))});
  assign MultLoop_acc_2310_nl = nl_MultLoop_acc_2310_nl[22:0];
  assign nl_MultLoop_acc_4143_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_2310_nl)))
      + (~ (data_rsci_idat[701:684]));
  assign MultLoop_acc_4143_nl = nl_MultLoop_acc_4143_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_181_itm_1 
      = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4140_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4620_nl)))
      + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1325_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4143_nl)));
  assign nl_MultLoop_acc_4144_nl =  -conv_s2s_16_17(data_rsci_idat[665:650]);
  assign MultLoop_acc_4144_nl = nl_MultLoop_acc_4144_nl[16:0];
  assign nl_MultLoop_acc_747_nl = conv_s2s_19_21({(MultLoop_acc_4144_nl) , (~ (data_rsci_idat[649:648]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[665:648])) , 2'b01});
  assign MultLoop_acc_747_nl = nl_MultLoop_acc_747_nl[20:0];
  assign nl_MultLoop_acc_4145_nl = conv_s2s_11_12(data_rsci_idat[629:619]) + 12'b000000000001;
  assign MultLoop_acc_4145_nl = nl_MultLoop_acc_4145_nl[11:0];
  assign nl_MultLoop_acc_2314_nl = conv_s2s_20_21({(data_rsci_idat[629:612]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[629:612]) + conv_s2s_17_21({(MultLoop_acc_4145_nl)
      , (data_rsci_idat[618:614])});
  assign MultLoop_acc_2314_nl = nl_MultLoop_acc_2314_nl[20:0];
  assign nl_MultLoop_acc_745_nl = conv_s2u_21_23(MultLoop_acc_2314_nl) + ({(~ (data_rsci_idat[629:612]))
      , 5'b00000});
  assign MultLoop_acc_745_nl = nl_MultLoop_acc_745_nl[22:0];
  assign nl_MultLoop_acc_2316_nl = conv_s2s_18_19(data_rsci_idat[557:540]) + conv_s2s_13_19({MultLoop_acc_4146_cse_1
      , (data_rsci_idat[547:546])});
  assign MultLoop_acc_2316_nl = nl_MultLoop_acc_2316_nl[18:0];
  assign nl_MultLoop_acc_741_nl = conv_s2u_19_20(MultLoop_acc_2316_nl) + ({(~ (data_rsci_idat[557:540]))
      , 2'b00});
  assign MultLoop_acc_741_nl = nl_MultLoop_acc_741_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_180_itm_1 
      = conv_s2s_16_18(MultLoop_acc_1324_itm_22_7) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_747_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_745_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_741_nl)));
  assign nl_MultLoop_acc_4621_nl = conv_s2u_15_19(MultLoop_acc_2317_itm_20_5[15:1])
      + conv_s2u_18_19(data_rsci_idat[503:486]);
  assign MultLoop_acc_4621_nl = nl_MultLoop_acc_4621_nl[18:0];
  assign nl_MultLoop_acc_1322_nl = conv_s2u_11_19(data_rsci_idat[521:511]) + conv_s2u_18_19(data_rsci_idat[521:504]);
  assign MultLoop_acc_1322_nl = nl_MultLoop_acc_1322_nl[18:0];
  assign nl_MultLoop_acc_2319_nl = ({(data_rsci_idat[467:450]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_678_18_7
      , (~ (data_rsci_idat[456:450]))});
  assign MultLoop_acc_2319_nl = nl_MultLoop_acc_2319_nl[19:0];
  assign nl_MultLoop_acc_2320_nl = conv_s2s_23_24({(data_rsci_idat[467:450]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_2319_nl);
  assign MultLoop_acc_2320_nl = nl_MultLoop_acc_2320_nl[23:0];
  assign nl_MultLoop_acc_4148_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_2320_nl)))
      + (~ (data_rsci_idat[467:450]));
  assign MultLoop_acc_4148_nl = nl_MultLoop_acc_4148_nl[17:0];
  assign nl_MultLoop_acc_734_nl = conv_s2s_23_24({(~ (data_rsci_idat[431:414])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[431:414])) , 3'b001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_788_18_5
      , (~ (data_rsci_idat[418:414]))});
  assign MultLoop_acc_734_nl = nl_MultLoop_acc_734_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_179_itm_1 
      = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4621_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1322_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4148_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_734_nl)));
  assign nl_MultLoop_acc_2334_nl = (~ (data_rsci_idat[89:72])) + conv_s2s_16_18({MultLoop_acc_3925_cse_1
      , (data_rsci_idat[78:75])});
  assign MultLoop_acc_2334_nl = nl_MultLoop_acc_2334_nl[17:0];
  assign nl_MultLoop_acc_1316_nl = conv_s2u_18_23(MultLoop_acc_2334_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[89:72])) , 4'b0001});
  assign MultLoop_acc_1316_nl = nl_MultLoop_acc_1316_nl[22:0];
  assign nl_MultLoop_acc_718_nl = conv_s2s_19_25({MultLoop_MultLoop_conc_792_18_6
      , (~ (data_rsci_idat[95:90]))}) + conv_s2s_24_25({(~ (data_rsci_idat[107:90]))
      , 6'b000001});
  assign MultLoop_acc_718_nl = nl_MultLoop_acc_718_nl[24:0];
  assign nl_MultLoop_acc_2324_nl = (~ (data_rsci_idat[269:252])) + conv_s2s_17_18({MultLoop_acc_4150_cse_1
      , (data_rsci_idat[259:254])});
  assign MultLoop_acc_2324_nl = nl_MultLoop_acc_2324_nl[17:0];
  assign nl_MultLoop_acc_2325_nl = ({(data_rsci_idat[269:252]) , 4'b0001}) + conv_s2s_18_22(MultLoop_acc_2324_nl);
  assign MultLoop_acc_2325_nl = nl_MultLoop_acc_2325_nl[21:0];
  assign nl_MultLoop_acc_4151_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2325_nl)))
      + (~ (data_rsci_idat[269:252]));
  assign MultLoop_acc_4151_nl = nl_MultLoop_acc_4151_nl[17:0];
  assign nl_MultLoop_acc_4152_nl = conv_s2s_12_13(data_rsci_idat[251:240]) + 13'b0000000000001;
  assign MultLoop_acc_4152_nl = nl_MultLoop_acc_4152_nl[12:0];
  assign nl_MultLoop_acc_2327_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_15_18({(MultLoop_acc_4152_nl)
      , (data_rsci_idat[239:238])});
  assign MultLoop_acc_2327_nl = nl_MultLoop_acc_2327_nl[17:0];
  assign nl_MultLoop_acc_1317_nl = conv_s2u_18_21(MultLoop_acc_2327_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[251:234])) , 2'b01});
  assign MultLoop_acc_1317_nl = nl_MultLoop_acc_1317_nl[20:0];
  assign nl_MultLoop_acc_2329_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_17_18({MultLoop_acc_4153_cse_1
      , (data_rsci_idat[151:146])});
  assign MultLoop_acc_2329_nl = nl_MultLoop_acc_2329_nl[17:0];
  assign nl_MultLoop_acc_2330_nl = ({(data_rsci_idat[161:144]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_2329_nl);
  assign MultLoop_acc_2330_nl = nl_MultLoop_acc_2330_nl[20:0];
  assign nl_MultLoop_acc_4154_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_2330_nl)))
      + (~ (data_rsci_idat[161:144]));
  assign MultLoop_acc_4154_nl = nl_MultLoop_acc_4154_nl[17:0];
  assign nl_MultLoop_acc_2332_nl = conv_s2s_23_24({(~ (data_rsci_idat[179:162]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[179:162])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[179:162]));
  assign MultLoop_acc_2332_nl = nl_MultLoop_acc_2332_nl[23:0];
  assign nl_MultLoop_acc_722_nl = conv_s2s_24_25(MultLoop_acc_2332_nl) + ({(data_rsci_idat[179:162])
      , 7'b0100000});
  assign MultLoop_acc_722_nl = nl_MultLoop_acc_722_nl[24:0];
  assign nl_MultLoop_acc_2338_nl = conv_s2s_20_21({(data_rsci_idat[53:36]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_2337_cse_1);
  assign MultLoop_acc_2338_nl = nl_MultLoop_acc_2338_nl[20:0];
  assign nl_MultLoop_acc_715_nl = conv_s2u_21_23(MultLoop_acc_2338_nl) + ({(~ (data_rsci_idat[53:36]))
      , 5'b00000});
  assign MultLoop_acc_715_nl = nl_MultLoop_acc_715_nl[22:0];
  assign nl_MultLoop_acc_4670_nl = conv_s2u_18_19(data_rsci_idat[35:18]) + conv_s2u_15_19(MultLoop_acc_2340_itm_19_4[15:1]);
  assign MultLoop_acc_4670_nl = nl_MultLoop_acc_4670_nl[18:0];
  assign nl_MultLoop_acc_4159_nl = conv_s2u_16_18(readslicef_19_16_3((MultLoop_acc_4670_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_4159_nl = nl_MultLoop_acc_4159_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_185_itm_1 
      = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1316_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_718_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4151_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1317_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4154_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_722_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_715_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4159_nl)));
  assign nl_MultLoop_acc_407_nl = conv_s2s_26_27({(~ (data_rsci_idat[485:468])) ,
      8'b00000100}) + conv_s2s_20_27({(~ (data_rsci_idat[485:468])) , 2'b01}) + conv_s2s_19_27({MultLoop_MultLoop_conc_796_18_8
      , (~ (data_rsci_idat[475:468]))});
  assign MultLoop_acc_407_nl = nl_MultLoop_acc_407_nl[26:0];
  assign nl_MultLoop_acc_404_nl = conv_s2s_23_24({(~ (data_rsci_idat[431:414])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[431:414])) , 2'b01}) + conv_s2s_19_24({MultLoop_MultLoop_conc_788_18_5
      , (~ (data_rsci_idat[418:414]))});
  assign MultLoop_acc_404_nl = nl_MultLoop_acc_404_nl[23:0];
  assign nl_MultLoop_acc_3087_nl = ({(data_rsci_idat[395:378]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_818_18_7
      , (~ (data_rsci_idat[384:378]))});
  assign MultLoop_acc_3087_nl = nl_MultLoop_acc_3087_nl[19:0];
  assign nl_MultLoop_acc_3088_nl = ({(~ (data_rsci_idat[395:378])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_3087_nl);
  assign MultLoop_acc_3088_nl = nl_MultLoop_acc_3088_nl[21:0];
  assign nl_MultLoop_acc_402_nl = conv_s2s_22_26(MultLoop_acc_3088_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[395:378])) , 7'b0010000});
  assign MultLoop_acc_402_nl = nl_MultLoop_acc_402_nl[25:0];
  assign nl_MultLoop_acc_4350_nl =  -conv_s2s_15_16(data_rsci_idat[323:309]);
  assign MultLoop_acc_4350_nl = nl_MultLoop_acc_4350_nl[15:0];
  assign nl_MultLoop_acc_398_nl = conv_s2s_19_22({(MultLoop_acc_4350_nl) , (~ (data_rsci_idat[308:306]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[323:306])) , 3'b001});
  assign MultLoop_acc_398_nl = nl_MultLoop_acc_398_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_407_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_404_nl))) + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_402_nl)))
      + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_398_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl[17:0];
  assign nl_MultLoop_acc_419_nl = conv_s2s_26_27({(~ (data_rsci_idat[701:684])) ,
      8'b00100000}) + conv_s2s_23_27({(~ (data_rsci_idat[701:684])) , 5'b00100})
      + conv_s2s_20_27({(~ (data_rsci_idat[701:684])) , 2'b01}) + conv_s2s_19_27({MultLoop_MultLoop_conc_782_18_8
      , (~ (data_rsci_idat[691:684]))});
  assign MultLoop_acc_419_nl = nl_MultLoop_acc_419_nl[26:0];
  assign nl_MultLoop_acc_414_nl = conv_s2s_26_27({(~ (data_rsci_idat[611:594])) ,
      8'b01000000}) + conv_s2s_24_27({(~ (data_rsci_idat[611:594])) , 6'b000100})
      + conv_s2s_21_27(Result_acc_129_cse_1);
  assign MultLoop_acc_414_nl = nl_MultLoop_acc_414_nl[26:0];
  assign nl_MultLoop_acc_3078_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_16_18({MultLoop_acc_4094_cse_1
      , (data_rsci_idat[562:561])});
  assign MultLoop_acc_3078_nl = nl_MultLoop_acc_3078_nl[17:0];
  assign nl_MultLoop_acc_1219_nl = conv_s2u_18_21(MultLoop_acc_3078_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[575:558])) , 2'b01});
  assign MultLoop_acc_1219_nl = nl_MultLoop_acc_1219_nl[20:0];
  assign nl_MultLoop_acc_409_nl = conv_s2s_25_26({(~ (data_rsci_idat[521:504])) ,
      7'b0010000}) + conv_s2s_22_26({(~ (data_rsci_idat[521:504])) , 4'b0100}) +
      conv_s2s_20_26({(~ (data_rsci_idat[521:504])) , 2'b01}) + conv_s2s_19_26({MultLoop_MultLoop_conc_726_18_7
      , (~ (data_rsci_idat[510:504]))});
  assign MultLoop_acc_409_nl = nl_MultLoop_acc_409_nl[25:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_281_itm_1 
      = (nnet_product_input_t_config2_weight_t_config2_accum_t_acc_276_nl) + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_419_nl)))
      + conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_414_nl))) + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1219_nl)))
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_409_nl)));
  assign nl_MultLoop_acc_3091_nl = (~ (data_rsci_idat[287:270])) + conv_s2s_15_18({MultLoop_acc_3976_cse_1
      , (data_rsci_idat[277:274])});
  assign MultLoop_acc_3091_nl = nl_MultLoop_acc_3091_nl[17:0];
  assign nl_MultLoop_acc_1215_nl = conv_s2u_18_23(MultLoop_acc_3091_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[287:270])) , 4'b0001});
  assign MultLoop_acc_1215_nl = nl_MultLoop_acc_1215_nl[22:0];
  assign nl_MultLoop_acc_389_nl = conv_s2u_16_18(data_rsci_idat[143:128]) - (data_rsci_idat[143:126]);
  assign MultLoop_acc_389_nl = nl_MultLoop_acc_389_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_245_itm_1 
      = conv_s2s_14_15(MultLoop_acc_1227_itm_21_5[16:3]) + conv_s2s_13_15(MultLoop_acc_400_itm_22_7[15:3])
      + conv_s2s_13_15(readslicef_18_13_5((MultLoop_acc_389_nl)));
  assign nl_MultLoop_acc_3026_nl = ({(data_rsci_idat[791:774]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_676_18_6
      , (~ (data_rsci_idat[779:774]))});
  assign MultLoop_acc_3026_nl = nl_MultLoop_acc_3026_nl[21:0];
  assign nl_MultLoop_acc_4353_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_3026_nl)))
      + (~ (data_rsci_idat[791:774]));
  assign MultLoop_acc_4353_nl = nl_MultLoop_acc_4353_nl[17:0];
  assign nl_MultLoop_acc_4679_nl = conv_s2u_18_19(data_rsci_idat[755:738]) + conv_s2u_16_19(MultLoop_acc_2906_itm_19_4);
  assign MultLoop_acc_4679_nl = nl_MultLoop_acc_4679_nl[18:0];
  assign nl_MultLoop_acc_4355_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_4679_nl)))
      + (~ (data_rsci_idat[755:738]));
  assign MultLoop_acc_4355_nl = nl_MultLoop_acc_4355_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_244_itm_1 
      = conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_4353_nl))) + conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_4355_nl)));
  assign nl_MultLoop_acc_405_nl = conv_s2s_18_24(~ (data_rsci_idat[449:432])) + ({(data_rsci_idat[449:432])
      , 6'b000001});
  assign MultLoop_acc_405_nl = nl_MultLoop_acc_405_nl[23:0];
  assign nl_MultLoop_acc_3031_nl = ({(data_rsci_idat[305:288]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_674_18_5
      , (~ (data_rsci_idat[292:288]))});
  assign MultLoop_acc_3031_nl = nl_MultLoop_acc_3031_nl[20:0];
  assign nl_MultLoop_acc_397_nl = conv_s2s_21_23(MultLoop_acc_3031_nl) + ({(~ (data_rsci_idat[305:288]))
      , 5'b00000});
  assign MultLoop_acc_397_nl = nl_MultLoop_acc_397_nl[22:0];
  assign nl_MultLoop_acc_4357_nl = conv_s2s_13_14(data_rsci_idat[179:167]) + 14'b00000000000001;
  assign MultLoop_acc_4357_nl = nl_MultLoop_acc_4357_nl[13:0];
  assign nl_MultLoop_acc_3033_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_17_18({(MultLoop_acc_4357_nl)
      , (data_rsci_idat[166:164])});
  assign MultLoop_acc_3033_nl = nl_MultLoop_acc_3033_nl[17:0];
  assign nl_MultLoop_acc_1212_nl = conv_s2u_18_22(MultLoop_acc_3033_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[179:162])) , 3'b001});
  assign MultLoop_acc_1212_nl = nl_MultLoop_acc_1212_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_253_itm_1 
      = conv_s2s_14_16(data_rsci_idat[215:202]) + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_405_nl)))
      + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_397_nl))) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_1212_nl)));
  assign nl_MultLoop_acc_1226_nl = conv_s2u_13_19(data_rsci_idat[737:725]) + conv_s2u_18_19(data_rsci_idat[737:720]);
  assign MultLoop_acc_1226_nl = nl_MultLoop_acc_1226_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_252_itm_1 
      = conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_1226_nl))) + conv_s2s_15_16(MultLoop_acc_1191_itm_21_7);
  assign nl_MultLoop_acc_3034_nl = (~ (data_rsci_idat[665:648])) + conv_s2s_15_18(data_rsci_idat[665:651]);
  assign MultLoop_acc_3034_nl = nl_MultLoop_acc_3034_nl[17:0];
  assign nl_MultLoop_acc_1223_nl = conv_s2u_18_22(MultLoop_acc_3034_nl) + ({(data_rsci_idat[665:648])
      , 4'b0001});
  assign MultLoop_acc_1223_nl = nl_MultLoop_acc_1223_nl[21:0];
  assign nl_MultLoop_acc_3035_nl = (~ (data_rsci_idat[683:666])) + conv_s2s_16_18(data_rsci_idat[683:668]);
  assign MultLoop_acc_3035_nl = nl_MultLoop_acc_3035_nl[17:0];
  assign nl_MultLoop_acc_1224_nl = conv_s2u_18_21(MultLoop_acc_3035_nl) + ({(data_rsci_idat[683:666])
      , 3'b001});
  assign MultLoop_acc_1224_nl = nl_MultLoop_acc_1224_nl[20:0];
  assign nl_MultLoop_acc_3036_nl = (~ (data_rsci_idat[629:612])) + conv_s2s_13_18(data_rsci_idat[629:617]);
  assign MultLoop_acc_3036_nl = nl_MultLoop_acc_3036_nl[17:0];
  assign nl_MultLoop_acc_1221_nl = conv_s2u_18_20(MultLoop_acc_3036_nl) + ({(data_rsci_idat[629:612])
      , 2'b01});
  assign MultLoop_acc_1221_nl = nl_MultLoop_acc_1221_nl[19:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_263_itm_1 
      = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1223_nl))) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1224_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1221_nl))) + conv_s2s_15_17(MultLoop_acc_408_itm_23_9);
  assign nl_MultLoop_acc_3038_nl = conv_s2s_18_19(data_rsci_idat[413:396]) + conv_s2s_17_19({MultLoop_acc_4032_cse_1
      , (data_rsci_idat[400:398])});
  assign MultLoop_acc_3038_nl = nl_MultLoop_acc_3038_nl[18:0];
  assign nl_MultLoop_acc_403_nl = conv_s2u_19_21(MultLoop_acc_3038_nl) + ({(~ (data_rsci_idat[413:396]))
      , 3'b000});
  assign MultLoop_acc_403_nl = nl_MultLoop_acc_403_nl[20:0];
  assign nl_MultLoop_acc_3040_nl = conv_s2s_23_24({(~ (data_rsci_idat[233:216]))
      , 5'b01000}) + conv_s2s_22_24(MultLoop_acc_2592_cse_1);
  assign MultLoop_acc_3040_nl = nl_MultLoop_acc_3040_nl[23:0];
  assign nl_MultLoop_acc_393_nl = conv_s2s_24_25(MultLoop_acc_3040_nl) + ({(data_rsci_idat[233:216])
      , 7'b0100000});
  assign MultLoop_acc_393_nl = nl_MultLoop_acc_393_nl[24:0];
  assign nl_MultLoop_acc_4359_nl = conv_s2s_14_15(data_rsci_idat[197:184]) + 15'b000000000000001;
  assign MultLoop_acc_4359_nl = nl_MultLoop_acc_4359_nl[14:0];
  assign nl_MultLoop_acc_3042_nl = (~ (data_rsci_idat[197:180])) + conv_s2s_17_18({(MultLoop_acc_4359_nl)
      , (data_rsci_idat[183:182])});
  assign MultLoop_acc_3042_nl = nl_MultLoop_acc_3042_nl[17:0];
  assign nl_MultLoop_acc_1213_nl = conv_s2u_18_21(MultLoop_acc_3042_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[197:180])) , 2'b01});
  assign MultLoop_acc_1213_nl = nl_MultLoop_acc_1213_nl[20:0];
  assign nl_MultLoop_acc_3044_nl = conv_s2s_18_19(data_rsci_idat[161:144]) + conv_s2s_16_19({MultLoop_acc_4162_cse_1
      , (data_rsci_idat[150:147])});
  assign MultLoop_acc_3044_nl = nl_MultLoop_acc_3044_nl[18:0];
  assign nl_MultLoop_acc_390_nl = conv_s2u_19_22(MultLoop_acc_3044_nl) + ({(~ (data_rsci_idat[161:144]))
      , 4'b0000});
  assign MultLoop_acc_390_nl = nl_MultLoop_acc_390_nl[21:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_262_itm_1 
      = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_403_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_393_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1213_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_390_nl)));
  assign nl_MultLoop_acc_3053_nl = conv_s2s_20_21({(~ (data_rsci_idat[845:828]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2604_cse_1);
  assign MultLoop_acc_3053_nl = nl_MultLoop_acc_3053_nl[20:0];
  assign nl_MultLoop_acc_1228_nl = conv_s2u_21_24(MultLoop_acc_3053_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[845:828])) , 5'b00100});
  assign MultLoop_acc_1228_nl = nl_MultLoop_acc_1228_nl[23:0];
  assign nl_MultLoop_acc_3046_nl = ({(data_rsci_idat[125:108]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_832_18_7
      , (~ (data_rsci_idat[114:108]))});
  assign MultLoop_acc_3046_nl = nl_MultLoop_acc_3046_nl[19:0];
  assign nl_MultLoop_acc_3047_nl = conv_s2s_23_24({(data_rsci_idat[125:108]) , 5'b00000})
      + conv_s2s_20_24(MultLoop_acc_3046_nl);
  assign MultLoop_acc_3047_nl = nl_MultLoop_acc_3047_nl[23:0];
  assign nl_MultLoop_acc_4362_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_3047_nl)))
      + (~ (data_rsci_idat[125:108]));
  assign MultLoop_acc_4362_nl = nl_MultLoop_acc_4362_nl[17:0];
  assign nl_MultLoop_acc_3049_nl = ({(data_rsci_idat[17:0]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_708_18_6
      , (~ (data_rsci_idat[5:0]))});
  assign MultLoop_acc_3049_nl = nl_MultLoop_acc_3049_nl[19:0];
  assign nl_MultLoop_acc_3050_nl = ({(~ (data_rsci_idat[17:0])) , 4'b0000}) + conv_s2s_20_22(MultLoop_acc_3049_nl);
  assign MultLoop_acc_3050_nl = nl_MultLoop_acc_3050_nl[21:0];
  assign nl_MultLoop_acc_382_nl = conv_s2s_22_25(MultLoop_acc_3050_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[17:0])) , 6'b010000});
  assign MultLoop_acc_382_nl = nl_MultLoop_acc_382_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_261_itm_1 
      = conv_s2s_16_17(readslicef_24_16_8((MultLoop_acc_1228_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4362_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_382_nl)));
  assign nl_MultLoop_acc_3055_nl = ({(data_rsci_idat[827:810]) , 3'b001}) + conv_s2s_19_21({MultLoop_acc_4133_itm
      , (~ (data_rsci_idat[816:810]))});
  assign MultLoop_acc_3055_nl = nl_MultLoop_acc_3055_nl[20:0];
  assign nl_MultLoop_acc_4366_nl = conv_s2u_14_18(readslicef_21_14_7((MultLoop_acc_3055_nl)))
      + (~ (data_rsci_idat[827:810]));
  assign MultLoop_acc_4366_nl = nl_MultLoop_acc_4366_nl[17:0];
  assign nl_MultLoop_acc_3057_nl = conv_s2s_20_21({(~ (data_rsci_idat[593:576]))
      , 2'b01}) + conv_s2s_18_21(Result_acc_152_cse_1);
  assign MultLoop_acc_3057_nl = nl_MultLoop_acc_3057_nl[20:0];
  assign nl_MultLoop_acc_1220_nl = conv_s2u_21_23(MultLoop_acc_3057_nl) + ({(data_rsci_idat[593:576])
      , 5'b00100});
  assign MultLoop_acc_1220_nl = nl_MultLoop_acc_1220_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_260_itm_1 
      = conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4366_nl))) + conv_s2s_16_17(readslicef_23_16_7((MultLoop_acc_1220_nl)));
  assign nl_MultLoop_acc_1218_nl = conv_s2u_12_19(data_rsci_idat[557:546]) + conv_s2u_18_19(data_rsci_idat[557:540]);
  assign MultLoop_acc_1218_nl = nl_MultLoop_acc_1218_nl[18:0];
  assign nl_MultLoop_acc_3059_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_17_18({MultLoop_MultLoop_conc_736_16_5
      , (data_rsci_idat[366:362])});
  assign MultLoop_acc_3059_nl = nl_MultLoop_acc_3059_nl[17:0];
  assign nl_MultLoop_acc_3060_nl = ({(data_rsci_idat[377:360]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_3059_nl);
  assign MultLoop_acc_3060_nl = nl_MultLoop_acc_3060_nl[20:0];
  assign nl_MultLoop_acc_401_nl = conv_s2u_21_23(MultLoop_acc_3060_nl) + ({(~ (data_rsci_idat[377:360]))
      , 5'b00000});
  assign MultLoop_acc_401_nl = nl_MultLoop_acc_401_nl[22:0];
  assign nl_MultLoop_acc_4680_nl = conv_s2u_16_19(MultLoop_acc_3062_itm_19_4) + conv_s2u_18_19(data_rsci_idat[341:324]);
  assign MultLoop_acc_4680_nl = nl_MultLoop_acc_4680_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_272_itm_1 
      = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1218_nl))) + conv_s2s_16_18(MultLoop_acc_1200_itm_19_4)
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_401_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4680_nl)));
  assign nl_MultLoop_acc_423_nl = conv_s2s_26_27({(~ (data_rsci_idat[773:756])) ,
      8'b00100000}) + conv_s2s_23_27({(~ (data_rsci_idat[773:756])) , 5'b01000})
      + conv_s2s_21_27({(~ (data_rsci_idat[773:756])) , 3'b001}) + conv_s2s_19_27({MultLoop_MultLoop_conc_846_18_8
      , (~ (data_rsci_idat[763:756]))});
  assign MultLoop_acc_423_nl = nl_MultLoop_acc_423_nl[26:0];
  assign nl_MultLoop_acc_3066_nl = ({(data_rsci_idat[35:18]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_780_18_8
      , (~ (data_rsci_idat[25:18]))});
  assign MultLoop_acc_3066_nl = nl_MultLoop_acc_3066_nl[20:0];
  assign nl_MultLoop_acc_3067_nl = conv_s2s_24_25({(data_rsci_idat[35:18]) , 6'b000000})
      + conv_s2s_21_25(MultLoop_acc_3066_nl);
  assign MultLoop_acc_3067_nl = nl_MultLoop_acc_3067_nl[24:0];
  assign nl_MultLoop_acc_4369_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_3067_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_4369_nl = nl_MultLoop_acc_4369_nl[17:0];
  assign nl_MultLoop_acc_1214_nl = conv_s2u_18_23(MultLoop_acc_3063_cse_1) + ({(data_rsci_idat[269:252])
      , 5'b00001});
  assign MultLoop_acc_1214_nl = nl_MultLoop_acc_1214_nl[22:0];
  assign nl_MultLoop_acc_4635_nl = conv_s2u_16_19(MultLoop_acc_2802_itm_19_4) + conv_s2u_18_19(data_rsci_idat[251:234]);
  assign MultLoop_acc_4635_nl = nl_MultLoop_acc_4635_nl[18:0];
  assign nl_MultLoop_acc_385_nl = conv_s2u_13_18(data_rsci_idat[53:41]) - (data_rsci_idat[53:36]);
  assign MultLoop_acc_385_nl = nl_MultLoop_acc_385_nl[17:0];
  assign nl_MultLoop_acc_428_nl = conv_s2u_14_18(data_rsci_idat[863:850]) - (data_rsci_idat[863:846]);
  assign MultLoop_acc_428_nl = nl_MultLoop_acc_428_nl[17:0];
  assign nl_MultLoop_acc_1222_nl = conv_s2u_15_19(data_rsci_idat[647:633]) + conv_s2u_18_19(data_rsci_idat[647:630]);
  assign MultLoop_acc_1222_nl = nl_MultLoop_acc_1222_nl[18:0];
  assign nl_MultLoop_acc_386_nl = conv_s2u_15_18(data_rsci_idat[71:57]) - (data_rsci_idat[71:54]);
  assign MultLoop_acc_386_nl = nl_MultLoop_acc_386_nl[17:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl = ~((data_rsci_idat[97:90]!=8'b00000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl = conv_s2s_10_11(~
      (data_rsci_idat[107:98])) + conv_u2s_9_11({8'b10001110 , (nnet_product_input_t_config2_weight_t_config2_accum_t_nor_3_nl)});
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl[10:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_278_itm_1 
      = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_423_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4369_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1214_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4635_nl)))
      + conv_s2s_16_18(MultLoop_acc_1211_itm_23_8) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_385_nl)))
      + conv_s2s_13_18(readslicef_18_13_5((MultLoop_acc_428_nl))) + conv_s2s_13_18(readslicef_19_13_6((MultLoop_acc_1222_nl)))
      + conv_s2s_13_18(MultLoop_acc_410_itm_20_7[13:1]) + conv_s2s_12_18(readslicef_18_12_6((MultLoop_acc_386_nl)))
      + conv_s2s_11_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_237_nl);
  assign nl_MultLoop_acc_2411_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_17_18({MultLoop_acc_4162_cse_1
      , (data_rsci_idat[150:146])});
  assign MultLoop_acc_2411_nl = nl_MultLoop_acc_2411_nl[17:0];
  assign nl_MultLoop_acc_1307_nl = conv_s2u_18_24(MultLoop_acc_2411_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[161:144])) , 5'b00001});
  assign MultLoop_acc_1307_nl = nl_MultLoop_acc_1307_nl[23:0];
  assign nl_MultLoop_acc_2413_nl = conv_s2s_20_21({(data_rsci_idat[125:108]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_2412_cse_1);
  assign MultLoop_acc_2413_nl = nl_MultLoop_acc_2413_nl[20:0];
  assign nl_MultLoop_acc_1305_nl = conv_s2u_21_23(MultLoop_acc_2413_nl) + conv_s2u_22_23({(data_rsci_idat[125:108])
      , 4'b0000});
  assign MultLoop_acc_1305_nl = nl_MultLoop_acc_1305_nl[22:0];
  assign nl_MultLoop_acc_2406_nl = (~ (data_rsci_idat[431:414])) + conv_s2s_17_18({MultLoop_MultLoop_conc_680_16_6
      , (data_rsci_idat[421:416])});
  assign MultLoop_acc_2406_nl = nl_MultLoop_acc_2406_nl[17:0];
  assign nl_MultLoop_acc_2408_nl = ({(data_rsci_idat[431:414]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[431:414])) , 2'b01}) + conv_s2s_18_22(MultLoop_acc_2406_nl);
  assign MultLoop_acc_2408_nl = nl_MultLoop_acc_2408_nl[21:0];
  assign nl_MultLoop_acc_4161_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2408_nl)))
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_4161_nl = nl_MultLoop_acc_4161_nl[17:0];
  assign nl_MultLoop_acc_4671_nl = conv_s2u_19_24(MultLoop_acc_2409_itm_20_2_1) +
      ({(data_rsci_idat[377:360]) , 6'b000001});
  assign MultLoop_acc_4671_nl = nl_MultLoop_acc_4671_nl[23:0];
  assign nl_MultLoop_acc_682_nl = conv_s2s_18_25(~ (data_rsci_idat[341:324])) + ({(data_rsci_idat[341:324])
      , 7'b0000001});
  assign MultLoop_acc_682_nl = nl_MultLoop_acc_682_nl[24:0];
  assign nl_MultLoop_acc_2415_nl = ({(~ (data_rsci_idat[143:126])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[143:126])
      + conv_s2s_16_20(data_rsci_idat[143:128]);
  assign MultLoop_acc_2415_nl = nl_MultLoop_acc_2415_nl[19:0];
  assign nl_MultLoop_acc_2416_nl = conv_s2s_22_23({(~ (data_rsci_idat[143:126]))
      , 4'b0100}) + conv_s2s_20_23(MultLoop_acc_2415_nl);
  assign MultLoop_acc_2416_nl = nl_MultLoop_acc_2416_nl[22:0];
  assign nl_MultLoop_acc_1306_nl = conv_s2u_23_24(MultLoop_acc_2416_nl) + ({(data_rsci_idat[143:126])
      , 6'b010000});
  assign MultLoop_acc_1306_nl = nl_MultLoop_acc_1306_nl[23:0];
  assign nl_MultLoop_acc_2418_nl = ({(data_rsci_idat[107:90]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_822_18_7
      , (~ (data_rsci_idat[96:90]))});
  assign MultLoop_acc_2418_nl = nl_MultLoop_acc_2418_nl[21:0];
  assign nl_MultLoop_acc_4164_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_2418_nl)))
      + (~ (data_rsci_idat[107:90]));
  assign MultLoop_acc_4164_nl = nl_MultLoop_acc_4164_nl[17:0];
  assign nl_MultLoop_acc_2470_itm_1  = conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1307_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1305_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4161_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_4671_nl))) + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_682_nl)))
      + conv_s2s_16_18(MultLoop_acc_400_itm_22_7) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1306_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4164_nl)));
  assign nl_MultLoop_acc_2425_nl = ({(~ (data_rsci_idat[539:522])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2424_cse_1);
  assign MultLoop_acc_2425_nl = nl_MultLoop_acc_2425_nl[19:0];
  assign nl_MultLoop_acc_1310_nl = conv_s2u_20_24(MultLoop_acc_2425_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[539:522])) , 5'b00100});
  assign MultLoop_acc_1310_nl = nl_MultLoop_acc_1310_nl[23:0];
  assign nl_MultLoop_acc_4168_nl = conv_s2u_15_19(MultLoop_acc_1730_itm_22_7[15:1])
      + conv_s2u_18_19(data_rsci_idat[395:378]);
  assign MultLoop_acc_4168_nl = nl_MultLoop_acc_4168_nl[18:0];
  assign nl_MultLoop_acc_2427_nl = ({(data_rsci_idat[251:234]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[251:234]));
  assign MultLoop_acc_2427_nl = nl_MultLoop_acc_2427_nl[20:0];
  assign nl_MultLoop_acc_677_nl = conv_s2s_21_25(MultLoop_acc_2427_nl) + conv_s2s_24_25({(data_rsci_idat[251:234])
      , 6'b000000});
  assign MultLoop_acc_677_nl = nl_MultLoop_acc_677_nl[24:0];
  assign nl_MultLoop_acc_1303_nl = conv_s2u_18_22(MultLoop_acc_2259_cse_1) + ({(data_rsci_idat[53:36])
      , 4'b0001});
  assign MultLoop_acc_1303_nl = nl_MultLoop_acc_1303_nl[21:0];
  assign nl_MultLoop_acc_2421_nl = ({(data_rsci_idat[71:54]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_758_18_6
      , (~ (data_rsci_idat[59:54]))});
  assign MultLoop_acc_2421_nl = nl_MultLoop_acc_2421_nl[19:0];
  assign nl_MultLoop_acc_2422_nl = conv_s2s_22_23({(data_rsci_idat[71:54]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2421_nl);
  assign MultLoop_acc_2422_nl = nl_MultLoop_acc_2422_nl[22:0];
  assign nl_MultLoop_acc_4166_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2422_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_4166_nl = nl_MultLoop_acc_4166_nl[17:0];
  assign nl_MultLoop_acc_2469_itm_1  = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1310_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4168_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_677_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1303_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4166_nl)));
  assign nl_MultLoop_acc_4169_nl =  -conv_s2s_10_11(data_rsci_idat[17:8]);
  assign MultLoop_acc_4169_nl = nl_MultLoop_acc_4169_nl[10:0];
  assign nl_MultLoop_acc_663_nl = conv_s2s_26_27({(~ (data_rsci_idat[17:0])) , 8'b00010000})
      + conv_s2s_22_27({(~ (data_rsci_idat[17:0])) , 4'b0001}) + conv_s2s_19_27({(MultLoop_acc_4169_nl)
      , (~ (data_rsci_idat[7:0]))});
  assign MultLoop_acc_663_nl = nl_MultLoop_acc_663_nl[26:0];
  assign nl_MultLoop_acc_694_nl = conv_s2u_13_18(data_rsci_idat[557:545]) - (data_rsci_idat[557:540]);
  assign MultLoop_acc_694_nl = nl_MultLoop_acc_694_nl[17:0];
  assign nl_MultLoop_acc_4170_nl = conv_s2s_13_14(data_rsci_idat[35:23]) + 14'b00000000000001;
  assign MultLoop_acc_4170_nl = nl_MultLoop_acc_4170_nl[13:0];
  assign nl_MultLoop_acc_2353_nl = conv_s2s_18_19(data_rsci_idat[35:18]) + conv_s2s_16_19({(MultLoop_acc_4170_nl)
      , (data_rsci_idat[22:21])});
  assign MultLoop_acc_2353_nl = nl_MultLoop_acc_2353_nl[18:0];
  assign nl_MultLoop_acc_665_nl = conv_s2u_19_20(MultLoop_acc_2353_nl) + ({(~ (data_rsci_idat[35:18]))
      , 2'b00});
  assign MultLoop_acc_665_nl = nl_MultLoop_acc_665_nl[19:0];
  assign nl_MultLoop_acc_698_nl = conv_s2u_16_18(data_rsci_idat[629:614]) - (data_rsci_idat[629:612]);
  assign MultLoop_acc_698_nl = nl_MultLoop_acc_698_nl[17:0];
  assign nl_MultLoop_acc_2355_nl = ({(data_rsci_idat[233:216]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_702_18_6
      , (~ (data_rsci_idat[221:216]))});
  assign MultLoop_acc_2355_nl = nl_MultLoop_acc_2355_nl[20:0];
  assign nl_MultLoop_acc_4172_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_2355_nl)))
      + (~ (data_rsci_idat[233:216]));
  assign MultLoop_acc_4172_nl = nl_MultLoop_acc_4172_nl[17:0];
  assign nl_MultLoop_acc_1304_nl = conv_s2u_13_19(data_rsci_idat[89:77]) + conv_s2u_18_19(data_rsci_idat[89:72]);
  assign MultLoop_acc_1304_nl = nl_MultLoop_acc_1304_nl[18:0];
  assign nl_MultLoop_acc_2458_itm_1  = (readslicef_27_17_10((MultLoop_acc_663_nl)))
      + conv_s2s_14_17(readslicef_18_14_4((MultLoop_acc_694_nl))) + conv_s2s_13_17(readslicef_20_13_7((MultLoop_acc_665_nl)))
      + conv_s2s_12_17(readslicef_18_12_6((MultLoop_acc_698_nl))) + conv_s2s_14_17(readslicef_18_14_4((MultLoop_acc_4172_nl)))
      + conv_s2s_14_17(readslicef_19_14_5((MultLoop_acc_1304_nl)));
  assign nl_MultLoop_acc_2356_nl = (~ (data_rsci_idat[809:792])) + conv_s2s_16_18(data_rsci_idat[809:794]);
  assign MultLoop_acc_2356_nl = nl_MultLoop_acc_2356_nl[17:0];
  assign nl_MultLoop_acc_2357_nl = ({(data_rsci_idat[809:792]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2356_nl);
  assign MultLoop_acc_2357_nl = nl_MultLoop_acc_2357_nl[19:0];
  assign nl_MultLoop_acc_1314_nl = conv_s2u_20_23(MultLoop_acc_2357_nl) + conv_s2u_22_23({(data_rsci_idat[809:792])
      , 4'b0000});
  assign MultLoop_acc_1314_nl = nl_MultLoop_acc_1314_nl[22:0];
  assign nl_MultLoop_acc_2359_nl = ({(data_rsci_idat[737:720]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_830_18_6
      , (~ (data_rsci_idat[725:720]))});
  assign MultLoop_acc_2359_nl = nl_MultLoop_acc_2359_nl[19:0];
  assign nl_MultLoop_acc_2360_nl = ({(~ (data_rsci_idat[737:720])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2359_nl);
  assign MultLoop_acc_2360_nl = nl_MultLoop_acc_2360_nl[21:0];
  assign nl_MultLoop_acc_703_nl = conv_s2s_22_25(MultLoop_acc_2360_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[737:720])) , 6'b010000});
  assign MultLoop_acc_703_nl = nl_MultLoop_acc_703_nl[24:0];
  assign nl_MultLoop_acc_2362_nl = conv_s2s_18_19(data_rsci_idat[755:738]) + conv_s2s_15_19({MultLoop_acc_4076_cse_1
      , (data_rsci_idat[743:742])});
  assign MultLoop_acc_2362_nl = nl_MultLoop_acc_2362_nl[18:0];
  assign nl_MultLoop_acc_704_nl = conv_s2u_19_20(MultLoop_acc_2362_nl) + ({(~ (data_rsci_idat[755:738]))
      , 2'b00});
  assign MultLoop_acc_704_nl = nl_MultLoop_acc_704_nl[19:0];
  assign nl_MultLoop_acc_2457_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1314_nl)))
      + conv_s2s_15_17(MultLoop_acc_471_itm_21_7) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_703_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_704_nl)));
  assign nl_MultLoop_acc_690_nl = conv_s2s_24_25({(~ (data_rsci_idat[485:468])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[485:468])) , 4'b0100}) + conv_s2s_20_25({(~
      (data_rsci_idat[485:468])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_724_18_6
      , (~ (data_rsci_idat[473:468]))});
  assign MultLoop_acc_690_nl = nl_MultLoop_acc_690_nl[24:0];
  assign nl_MultLoop_acc_2366_nl = conv_s2s_21_22({(~ (data_rsci_idat[305:288]))
      , 3'b001}) + conv_s2s_18_22(~ (data_rsci_idat[305:288]));
  assign MultLoop_acc_2366_nl = nl_MultLoop_acc_2366_nl[21:0];
  assign nl_MultLoop_acc_680_nl = conv_s2s_22_24(MultLoop_acc_2366_nl) + ({(data_rsci_idat[305:288])
      , 6'b001000});
  assign MultLoop_acc_680_nl = nl_MultLoop_acc_680_nl[23:0];
  assign nl_MultLoop_acc_2438_itm_1  = conv_s2s_15_16(readslicef_25_15_10((MultLoop_acc_690_nl)))
      + conv_s2s_15_16(readslicef_24_15_9((MultLoop_acc_680_nl)));
  assign nl_MultLoop_acc_4176_nl =  -conv_s2s_12_13(data_rsci_idat[323:312]);
  assign MultLoop_acc_4176_nl = nl_MultLoop_acc_4176_nl[12:0];
  assign nl_MultLoop_acc_2368_nl = ({(data_rsci_idat[323:306]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4176_nl)
      , (~ (data_rsci_idat[311:306]))});
  assign MultLoop_acc_2368_nl = nl_MultLoop_acc_2368_nl[19:0];
  assign nl_MultLoop_acc_2369_nl = ({(~ (data_rsci_idat[323:306])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2368_nl);
  assign MultLoop_acc_2369_nl = nl_MultLoop_acc_2369_nl[21:0];
  assign nl_MultLoop_acc_681_nl = conv_s2s_22_25(MultLoop_acc_2369_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[323:306])) , 6'b010000});
  assign MultLoop_acc_681_nl = nl_MultLoop_acc_681_nl[24:0];
  assign nl_MultLoop_acc_4622_nl = conv_s2u_16_19(MultLoop_acc_2057_cse_1[18:3])
      + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_4622_nl = nl_MultLoop_acc_4622_nl[18:0];
  assign nl_MultLoop_acc_2437_itm_1  = conv_s2s_15_16(readslicef_25_15_10((MultLoop_acc_681_nl)))
      + conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_4622_nl)));
  assign nl_MultLoop_acc_2372_nl = ({(data_rsci_idat[197:180]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_862_18_6
      , (~ (data_rsci_idat[185:180]))});
  assign MultLoop_acc_2372_nl = nl_MultLoop_acc_2372_nl[19:0];
  assign nl_MultLoop_acc_2373_nl = conv_s2s_22_23({(data_rsci_idat[197:180]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2372_nl);
  assign MultLoop_acc_2373_nl = nl_MultLoop_acc_2373_nl[22:0];
  assign nl_MultLoop_acc_4178_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2373_nl)))
      + (~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_4178_nl = nl_MultLoop_acc_4178_nl[17:0];
  assign nl_MultLoop_acc_675_nl = conv_s2u_14_18(data_rsci_idat[215:202]) - (data_rsci_idat[215:198]);
  assign MultLoop_acc_675_nl = nl_MultLoop_acc_675_nl[17:0];
  assign nl_MultLoop_acc_673_nl = conv_s2u_13_18(data_rsci_idat[179:167]) - (data_rsci_idat[179:162]);
  assign MultLoop_acc_673_nl = nl_MultLoop_acc_673_nl[17:0];
  assign nl_MultLoop_acc_4179_nl = conv_s2s_10_11(data_rsci_idat[647:638]) + 11'b11111001011;
  assign MultLoop_acc_4179_nl = nl_MultLoop_acc_4179_nl[10:0];
  assign nl_MultLoop_acc_4180_nl =  -conv_s2s_16_17(data_rsci_idat[269:254]);
  assign MultLoop_acc_4180_nl = nl_MultLoop_acc_4180_nl[16:0];
  assign nl_MultLoop_acc_678_nl = conv_s2s_19_21({(MultLoop_acc_4180_nl) , (~ (data_rsci_idat[253:252]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[269:252])) , 2'b01});
  assign MultLoop_acc_678_nl = nl_MultLoop_acc_678_nl[20:0];
  assign nl_MultLoop_acc_2455_itm_1  = conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4178_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_675_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_673_nl)))
      + conv_s2s_13_17({(MultLoop_acc_4179_nl) , (data_rsci_idat[637:636])}) + conv_s2s_13_17(readslicef_21_13_8((MultLoop_acc_678_nl)));
  assign nl_MultLoop_acc_2376_nl = ({(data_rsci_idat[845:828]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2375_cse_1);
  assign MultLoop_acc_2376_nl = nl_MultLoop_acc_2376_nl[19:0];
  assign nl_MultLoop_acc_709_nl = conv_s2u_20_22(MultLoop_acc_2376_nl) + ({(~ (data_rsci_idat[845:828]))
      , 4'b0000});
  assign MultLoop_acc_709_nl = nl_MultLoop_acc_709_nl[21:0];
  assign nl_MultLoop_acc_708_nl = conv_s2u_13_18(data_rsci_idat[827:815]) - (data_rsci_idat[827:810]);
  assign MultLoop_acc_708_nl = nl_MultLoop_acc_708_nl[17:0];
  assign nl_MultLoop_acc_4182_nl = conv_s2s_10_11(data_rsci_idat[791:782]) + 11'b00000000001;
  assign MultLoop_acc_4182_nl = nl_MultLoop_acc_4182_nl[10:0];
  assign nl_MultLoop_acc_2378_nl = (~ (data_rsci_idat[791:774])) + conv_s2s_15_18({(MultLoop_acc_4182_nl)
      , (data_rsci_idat[781:778])});
  assign MultLoop_acc_2378_nl = nl_MultLoop_acc_2378_nl[17:0];
  assign nl_MultLoop_acc_2379_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2378_nl);
  assign MultLoop_acc_2379_nl = nl_MultLoop_acc_2379_nl[19:0];
  assign nl_MultLoop_acc_706_nl = conv_s2u_20_22(MultLoop_acc_2379_nl) + ({(~ (data_rsci_idat[791:774]))
      , 4'b0000});
  assign MultLoop_acc_706_nl = nl_MultLoop_acc_706_nl[21:0];
  assign nl_MultLoop_acc_2466_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_709_nl)))
      + conv_s2s_16_18(MultLoop_acc_1315_itm_19_4) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_708_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_706_nl)));
  assign nl_MultLoop_acc_2380_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_15_18(data_rsci_idat[701:687]);
  assign MultLoop_acc_2380_nl = nl_MultLoop_acc_2380_nl[17:0];
  assign nl_MultLoop_acc_1313_nl = conv_s2u_18_21(MultLoop_acc_2380_nl) + ({(data_rsci_idat[701:684])
      , 3'b001});
  assign MultLoop_acc_1313_nl = nl_MultLoop_acc_1313_nl[20:0];
  assign nl_MultLoop_acc_702_nl = conv_s2s_25_26({(~ (data_rsci_idat[719:702])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[719:702])) , 5'b01000}) +
      conv_s2s_21_26({(~ (data_rsci_idat[719:702])) , 3'b001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_840_18_7
      , (~ (data_rsci_idat[708:702]))});
  assign MultLoop_acc_702_nl = nl_MultLoop_acc_702_nl[25:0];
  assign nl_MultLoop_acc_2452_itm_1  = conv_s2s_16_17(readslicef_21_16_5((MultLoop_acc_1313_nl)))
      + conv_s2s_16_17(readslicef_26_16_10((MultLoop_acc_702_nl)));
  assign nl_MultLoop_acc_4623_nl = conv_s2u_16_19(MultLoop_acc_2073_cse_1[18:3])
      + conv_s2u_18_19(data_rsci_idat[665:648]);
  assign MultLoop_acc_4623_nl = nl_MultLoop_acc_4623_nl[18:0];
  assign nl_MultLoop_acc_2386_nl = conv_s2s_23_24({(~ (data_rsci_idat[683:666]))
      , 5'b00100}) + conv_s2s_21_24(MultLoop_acc_2385_cse_1);
  assign MultLoop_acc_2386_nl = nl_MultLoop_acc_2386_nl[23:0];
  assign nl_MultLoop_acc_700_nl = conv_s2s_24_25(MultLoop_acc_2386_nl) + ({(data_rsci_idat[683:666])
      , 7'b0100000});
  assign MultLoop_acc_700_nl = nl_MultLoop_acc_700_nl[24:0];
  assign nl_MultLoop_acc_2451_itm_1  = conv_s2s_16_17(readslicef_19_16_3((MultLoop_acc_4623_nl)))
      + conv_s2s_16_17(readslicef_25_16_9((MultLoop_acc_700_nl)));
  assign nl_MultLoop_acc_2389_nl = conv_s2s_24_25({(~ (data_rsci_idat[593:576]))
      , 6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[593:576])) , 4'b0100}) +
      conv_s2s_21_25(MultLoop_acc_2387_cse_1);
  assign MultLoop_acc_2389_nl = nl_MultLoop_acc_2389_nl[24:0];
  assign nl_MultLoop_acc_696_nl = conv_s2s_25_26(MultLoop_acc_2389_nl) + ({(data_rsci_idat[593:576])
      , 8'b01000000});
  assign MultLoop_acc_696_nl = nl_MultLoop_acc_696_nl[25:0];
  assign nl_MultLoop_acc_2391_nl = ({(~ (data_rsci_idat[575:558])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_2390_cse_1);
  assign MultLoop_acc_2391_nl = nl_MultLoop_acc_2391_nl[22:0];
  assign nl_MultLoop_acc_695_nl = conv_s2s_23_26(MultLoop_acc_2391_nl) + ({(data_rsci_idat[575:558])
      , 8'b00100000});
  assign MultLoop_acc_695_nl = nl_MultLoop_acc_695_nl[25:0];
  assign nl_MultLoop_acc_2394_nl = conv_s2s_21_22({(data_rsci_idat[521:504]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[521:504]) + conv_s2s_16_22({MultLoop_acc_3987_cse_1
      , (data_rsci_idat[511:507])});
  assign MultLoop_acc_2394_nl = nl_MultLoop_acc_2394_nl[21:0];
  assign nl_MultLoop_acc_692_nl = conv_s2u_22_23(MultLoop_acc_2394_nl) + ({(~ (data_rsci_idat[521:504]))
      , 5'b00000});
  assign MultLoop_acc_692_nl = nl_MultLoop_acc_692_nl[22:0];
  assign nl_MultLoop_acc_2464_itm_1  = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_696_nl)))
      + conv_s2s_16_18(MultLoop_acc_1154_itm_21_6) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_695_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_692_nl)));
  assign nl_MultLoop_acc_691_nl = conv_s2s_19_26({MultLoop_MultLoop_conc_716_18_7
      , (~ (data_rsci_idat[492:486]))}) + conv_s2s_25_26({(~ (data_rsci_idat[503:486]))
      , 7'b0000001});
  assign MultLoop_acc_691_nl = nl_MultLoop_acc_691_nl[25:0];
  assign nl_MultLoop_acc_2397_nl = (~ (data_rsci_idat[449:432])) + conv_s2s_17_18({MultLoop_acc_4186_cse_1
      , (data_rsci_idat[439:434])});
  assign MultLoop_acc_2397_nl = nl_MultLoop_acc_2397_nl[17:0];
  assign nl_MultLoop_acc_2398_nl = ({(data_rsci_idat[449:432]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2397_nl);
  assign MultLoop_acc_2398_nl = nl_MultLoop_acc_2398_nl[19:0];
  assign nl_MultLoop_acc_2399_nl = conv_s2s_22_23({(data_rsci_idat[449:432]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2398_nl);
  assign MultLoop_acc_2399_nl = nl_MultLoop_acc_2399_nl[22:0];
  assign nl_MultLoop_acc_4187_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2399_nl)))
      + (~ (data_rsci_idat[449:432]));
  assign MultLoop_acc_4187_nl = nl_MultLoop_acc_4187_nl[17:0];
  assign nl_MultLoop_acc_2402_nl = conv_s2s_20_21({(data_rsci_idat[467:450]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[467:450]) + conv_s2s_16_21({MultLoop_acc_4030_cse_1
      , (data_rsci_idat[457:453])});
  assign MultLoop_acc_2402_nl = nl_MultLoop_acc_2402_nl[20:0];
  assign nl_MultLoop_acc_689_nl = conv_s2u_21_23(MultLoop_acc_2402_nl) + ({(~ (data_rsci_idat[467:450]))
      , 5'b00000});
  assign MultLoop_acc_689_nl = nl_MultLoop_acc_689_nl[22:0];
  assign nl_MultLoop_acc_2404_nl = ({(data_rsci_idat[413:396]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2403_cse_1);
  assign MultLoop_acc_2404_nl = nl_MultLoop_acc_2404_nl[19:0];
  assign nl_MultLoop_acc_1309_nl = conv_s2u_20_23(MultLoop_acc_2404_nl) + conv_s2u_22_23({(data_rsci_idat[413:396])
      , 4'b0000});
  assign MultLoop_acc_1309_nl = nl_MultLoop_acc_1309_nl[22:0];
  assign nl_MultLoop_acc_2463_itm_1  = conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_691_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4187_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_689_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1309_nl)));
  assign nl_MultLoop_acc_465_nl = conv_s2s_19_27({MultLoop_MultLoop_conc_756_18_8
      , (~ (data_rsci_idat[655:648]))}) + conv_s2s_26_27({(~ (data_rsci_idat[665:648]))
      , 8'b00000001});
  assign MultLoop_acc_465_nl = nl_MultLoop_acc_465_nl[26:0];
  assign nl_MultLoop_acc_4634_nl = ({(data_rsci_idat[557:540]) , 3'b001}) + conv_s2u_19_21(MultLoop_acc_2669_itm_20_2_1);
  assign MultLoop_acc_4634_nl = nl_MultLoop_acc_4634_nl[20:0];
  assign nl_MultLoop_acc_4314_nl = conv_s2u_15_19(readslicef_21_15_6((MultLoop_acc_4634_nl)))
      + conv_s2u_18_19(data_rsci_idat[557:540]);
  assign MultLoop_acc_4314_nl = nl_MultLoop_acc_4314_nl[18:0];
  assign nl_MultLoop_acc_2968_nl = ({(~ (data_rsci_idat[521:504])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2967_cse_1);
  assign MultLoop_acc_2968_nl = nl_MultLoop_acc_2968_nl[19:0];
  assign nl_MultLoop_acc_2969_nl = ({(data_rsci_idat[521:504]) , 4'b0100}) + conv_s2s_20_22(MultLoop_acc_2968_nl);
  assign MultLoop_acc_2969_nl = nl_MultLoop_acc_2969_nl[21:0];
  assign nl_MultLoop_acc_1234_nl = conv_s2u_22_25(MultLoop_acc_2969_nl) + conv_s2u_24_25({(data_rsci_idat[521:504])
      , 6'b000000});
  assign MultLoop_acc_1234_nl = nl_MultLoop_acc_1234_nl[24:0];
  assign nl_MultLoop_acc_4315_nl =  -conv_s2s_14_15(data_rsci_idat[485:472]);
  assign MultLoop_acc_4315_nl = nl_MultLoop_acc_4315_nl[14:0];
  assign nl_MultLoop_acc_455_nl = conv_s2s_19_23({(MultLoop_acc_4315_nl) , (~ (data_rsci_idat[471:468]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[485:468])) , 4'b0001});
  assign MultLoop_acc_455_nl = nl_MultLoop_acc_455_nl[22:0];
  assign nl_MultLoop_acc_3018_itm_1  = conv_s2s_17_18(readslicef_27_17_10((MultLoop_acc_465_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4314_nl))) + conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1234_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_455_nl)));
  assign nl_MultLoop_acc_4316_nl = conv_s2s_11_12(data_rsci_idat[35:25]) + 12'b000000000001;
  assign MultLoop_acc_4316_nl = nl_MultLoop_acc_4316_nl[11:0];
  assign nl_MultLoop_acc_2973_nl = conv_s2s_20_21({(data_rsci_idat[35:18]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[35:18]) + conv_s2s_17_21({(MultLoop_acc_4316_nl)
      , (data_rsci_idat[24:20])});
  assign MultLoop_acc_2973_nl = nl_MultLoop_acc_2973_nl[20:0];
  assign nl_MultLoop_acc_430_nl = conv_s2u_21_23(MultLoop_acc_2973_nl) + ({(~ (data_rsci_idat[35:18]))
      , 5'b00000});
  assign MultLoop_acc_430_nl = nl_MultLoop_acc_430_nl[22:0];
  assign nl_MultLoop_acc_2976_nl = conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_430_nl)))
      + 16'b0000000011111101;
  assign MultLoop_acc_2976_nl = nl_MultLoop_acc_2976_nl[15:0];
  assign nl_MultLoop_acc_4317_nl =  -conv_s2s_11_12(data_rsci_idat[17:7]);
  assign MultLoop_acc_4317_nl = nl_MultLoop_acc_4317_nl[11:0];
  assign nl_MultLoop_acc_429_nl = conv_s2s_25_26({(~ (data_rsci_idat[17:0])) , 7'b0001000})
      + conv_s2s_21_26({(~ (data_rsci_idat[17:0])) , 3'b001}) + conv_s2s_19_26({(MultLoop_acc_4317_nl)
      , (~ (data_rsci_idat[6:0]))});
  assign MultLoop_acc_429_nl = nl_MultLoop_acc_429_nl[25:0];
  assign nl_MultLoop_434_MultLoop_acc_3_nl = conv_s2s_16_17(MultLoop_acc_2976_nl)
      + (readslicef_26_17_9((MultLoop_acc_429_nl)));
  assign MultLoop_434_MultLoop_acc_3_nl = nl_MultLoop_434_MultLoop_acc_3_nl[16:0];
  assign nl_MultLoop_acc_2979_nl = ({(~ (data_rsci_idat[53:36])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2337_cse_1);
  assign MultLoop_acc_2979_nl = nl_MultLoop_acc_2979_nl[19:0];
  assign nl_MultLoop_acc_1229_nl = conv_s2u_20_24(MultLoop_acc_2979_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[53:36])) , 5'b00100});
  assign MultLoop_acc_1229_nl = nl_MultLoop_acc_1229_nl[23:0];
  assign nl_MultLoop_acc_3008_itm_1  = conv_s2s_17_18(MultLoop_434_MultLoop_acc_3_nl)
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1229_nl)));
  assign nl_MultLoop_acc_4320_nl = conv_s2u_14_18(MultLoop_acc_2906_itm_19_4[15:2])
      + (~ (data_rsci_idat[755:738]));
  assign MultLoop_acc_4320_nl = nl_MultLoop_acc_4320_nl[17:0];
  assign nl_MultLoop_acc_4321_nl =  -conv_s2s_12_13(data_rsci_idat[719:708]);
  assign MultLoop_acc_4321_nl = nl_MultLoop_acc_4321_nl[12:0];
  assign nl_MultLoop_acc_2909_nl = ({(data_rsci_idat[719:702]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[719:702])) , 2'b01}) + conv_s2s_19_22({(MultLoop_acc_4321_nl)
      , (~ (data_rsci_idat[707:702]))});
  assign MultLoop_acc_2909_nl = nl_MultLoop_acc_2909_nl[21:0];
  assign nl_MultLoop_acc_4322_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2909_nl)))
      + (~ (data_rsci_idat[719:702]));
  assign MultLoop_acc_4322_nl = nl_MultLoop_acc_4322_nl[17:0];
  assign nl_MultLoop_acc_2984_itm_1  = conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_4320_nl)))
      + conv_s2s_14_15(readslicef_18_14_4((MultLoop_acc_4322_nl)));
  assign nl_MultLoop_acc_2912_nl = conv_s2s_20_21({(data_rsci_idat[611:594]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[611:594]) + conv_s2s_17_21({MultLoop_MultLoop_conc_774_16_4
      , (data_rsci_idat[599:596])});
  assign MultLoop_acc_2912_nl = nl_MultLoop_acc_2912_nl[20:0];
  assign nl_MultLoop_acc_462_nl = conv_s2u_21_22(MultLoop_acc_2912_nl) + ({(~ (data_rsci_idat[611:594]))
      , 4'b0000});
  assign MultLoop_acc_462_nl = nl_MultLoop_acc_462_nl[21:0];
  assign nl_MultLoop_acc_2983_itm_1  = conv_s2s_14_15(readslicef_22_14_8((MultLoop_acc_462_nl)))
      + conv_s2s_14_15(MultLoop_acc_410_itm_20_7);
  assign nl_MultLoop_acc_474_nl = conv_s2u_14_18(data_rsci_idat[827:814]) - (data_rsci_idat[827:810]);
  assign MultLoop_acc_474_nl = nl_MultLoop_acc_474_nl[17:0];
  assign nl_MultLoop_acc_2913_nl = (~ (data_rsci_idat[251:234])) + conv_s2s_15_18(data_rsci_idat[251:237]);
  assign MultLoop_acc_2913_nl = nl_MultLoop_acc_2913_nl[17:0];
  assign nl_MultLoop_acc_1231_nl = conv_s2u_18_21(MultLoop_acc_2913_nl) + ({(data_rsci_idat[251:234])
      , 3'b001});
  assign MultLoop_acc_1231_nl = nl_MultLoop_acc_1231_nl[20:0];
  assign nl_MultLoop_acc_4324_nl = conv_s2s_12_13(data_rsci_idat[215:204]) + 13'b0000000000001;
  assign MultLoop_acc_4324_nl = nl_MultLoop_acc_4324_nl[12:0];
  assign nl_MultLoop_acc_2915_nl = conv_s2s_18_19(data_rsci_idat[215:198]) + conv_s2s_16_19({(MultLoop_acc_4324_nl)
      , (data_rsci_idat[203:201])});
  assign MultLoop_acc_2915_nl = nl_MultLoop_acc_2915_nl[18:0];
  assign nl_MultLoop_acc_440_nl = conv_s2u_19_21(MultLoop_acc_2915_nl) + ({(~ (data_rsci_idat[215:198]))
      , 3'b000});
  assign MultLoop_acc_440_nl = nl_MultLoop_acc_440_nl[20:0];
  assign nl_MultLoop_acc_2993_itm_1  = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_474_nl)))
      + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1231_nl))) + conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_440_nl)));
  assign nl_MultLoop_acc_4325_nl =  -conv_s2s_13_14(data_rsci_idat[791:779]);
  assign MultLoop_acc_4325_nl = nl_MultLoop_acc_4325_nl[13:0];
  assign nl_MultLoop_acc_2917_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_19_20({(MultLoop_acc_4325_nl)
      , (~ (data_rsci_idat[778:774]))});
  assign MultLoop_acc_2917_nl = nl_MultLoop_acc_2917_nl[19:0];
  assign nl_MultLoop_acc_472_nl = conv_s2s_20_23(MultLoop_acc_2917_nl) + ({(~ (data_rsci_idat[791:774]))
      , 5'b00000});
  assign MultLoop_acc_472_nl = nl_MultLoop_acc_472_nl[22:0];
  assign nl_MultLoop_acc_4326_nl = conv_s2s_12_13(data_rsci_idat[737:726]) + 13'b0000000000001;
  assign MultLoop_acc_4326_nl = nl_MultLoop_acc_4326_nl[12:0];
  assign nl_MultLoop_acc_2919_nl = (~ (data_rsci_idat[737:720])) + conv_s2s_16_18({(MultLoop_acc_4326_nl)
      , (data_rsci_idat[725:723])});
  assign MultLoop_acc_2919_nl = nl_MultLoop_acc_2919_nl[17:0];
  assign nl_MultLoop_acc_1238_nl = conv_s2u_18_22(MultLoop_acc_2919_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[737:720])) , 3'b001});
  assign MultLoop_acc_1238_nl = nl_MultLoop_acc_1238_nl[21:0];
  assign nl_MultLoop_acc_2921_nl = ({(~ (data_rsci_idat[701:684])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_1940_cse_1);
  assign MultLoop_acc_2921_nl = nl_MultLoop_acc_2921_nl[21:0];
  assign nl_MultLoop_acc_467_nl = conv_s2s_22_25(MultLoop_acc_2921_nl) + ({(data_rsci_idat[701:684])
      , 7'b0010000});
  assign MultLoop_acc_467_nl = nl_MultLoop_acc_467_nl[24:0];
  assign nl_MultLoop_acc_3006_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_472_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1238_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_467_nl)))
      + conv_s2s_15_17(MultLoop_acc_1204_itm_19_5);
  assign nl_MultLoop_acc_460_nl = conv_s2s_19_25({MultLoop_MultLoop_conc_686_18_6
      , (~ (data_rsci_idat[563:558]))}) + conv_s2s_24_25({(~ (data_rsci_idat[575:558]))
      , 6'b000001});
  assign MultLoop_acc_460_nl = nl_MultLoop_acc_460_nl[24:0];
  assign nl_MultLoop_acc_456_nl = conv_s2s_24_25({(data_rsci_idat[503:486]) , 6'b000000})
      + conv_s2s_22_25({(data_rsci_idat[503:486]) , 4'b0000}) + conv_s2s_20_25(MultLoop_acc_2923_cse_1);
  assign MultLoop_acc_456_nl = nl_MultLoop_acc_456_nl[24:0];
  assign nl_MultLoop_acc_2926_nl = conv_s2s_23_24({(~ (data_rsci_idat[395:378]))
      , 5'b01000}) + conv_s2s_22_24(MultLoop_acc_2781_cse_1);
  assign MultLoop_acc_2926_nl = nl_MultLoop_acc_2926_nl[23:0];
  assign nl_MultLoop_acc_450_nl = conv_s2s_24_25(MultLoop_acc_2926_nl) + ({(data_rsci_idat[395:378])
      , 7'b0100000});
  assign MultLoop_acc_450_nl = nl_MultLoop_acc_450_nl[24:0];
  assign nl_MultLoop_acc_2927_nl = ({(data_rsci_idat[323:306]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[323:306]));
  assign MultLoop_acc_2927_nl = nl_MultLoop_acc_2927_nl[20:0];
  assign nl_MultLoop_acc_446_nl = conv_s2s_21_25(MultLoop_acc_2927_nl) + conv_s2s_24_25({(data_rsci_idat[323:306])
      , 6'b000000});
  assign MultLoop_acc_446_nl = nl_MultLoop_acc_446_nl[24:0];
  assign nl_MultLoop_acc_3005_itm_1  = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_460_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_456_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_450_nl)))
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_446_nl)));
  assign nl_MultLoop_acc_4328_nl = conv_s2s_12_13(data_rsci_idat[197:186]) + 13'b0000000000001;
  assign MultLoop_acc_4328_nl = nl_MultLoop_acc_4328_nl[12:0];
  assign nl_MultLoop_acc_2929_nl = (~ (data_rsci_idat[197:180])) + conv_s2s_17_18({(MultLoop_acc_4328_nl)
      , (data_rsci_idat[185:182])});
  assign MultLoop_acc_2929_nl = nl_MultLoop_acc_2929_nl[17:0];
  assign nl_MultLoop_acc_1230_nl = conv_s2u_18_23(MultLoop_acc_2929_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[197:180])) , 4'b0001});
  assign MultLoop_acc_1230_nl = nl_MultLoop_acc_1230_nl[22:0];
  assign nl_MultLoop_acc_2930_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[161:144]));
  assign MultLoop_acc_2930_nl = nl_MultLoop_acc_2930_nl[19:0];
  assign nl_MultLoop_acc_437_nl = conv_s2s_20_23(MultLoop_acc_2930_nl) + conv_s2s_22_23({(data_rsci_idat[161:144])
      , 4'b0000});
  assign MultLoop_acc_437_nl = nl_MultLoop_acc_437_nl[22:0];
  assign nl_MultLoop_acc_2932_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_850_18_6
      , (~ (data_rsci_idat[167:162]))});
  assign MultLoop_acc_2932_nl = nl_MultLoop_acc_2932_nl[19:0];
  assign nl_MultLoop_acc_2933_nl = ({(~ (data_rsci_idat[179:162])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2932_nl);
  assign MultLoop_acc_2933_nl = nl_MultLoop_acc_2933_nl[21:0];
  assign nl_MultLoop_acc_438_nl = conv_s2s_22_25(MultLoop_acc_2933_nl) + conv_s2s_24_25({(~
      (data_rsci_idat[179:162])) , 6'b010000});
  assign MultLoop_acc_438_nl = nl_MultLoop_acc_438_nl[24:0];
  assign nl_MultLoop_acc_3004_itm_1  = conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1230_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_437_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_438_nl)))
      + conv_s2s_15_17(MultLoop_acc_2252_itm_20_5[15:1]);
  assign nl_MultLoop_acc_2934_nl = conv_s2s_22_23({(~ (data_rsci_idat[143:126]))
      , 4'b0001}) + conv_s2s_18_23(~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_2934_nl = nl_MultLoop_acc_2934_nl[22:0];
  assign nl_MultLoop_acc_436_nl = conv_s2s_23_25(MultLoop_acc_2934_nl) + ({(data_rsci_idat[143:126])
      , 7'b0010000});
  assign MultLoop_acc_436_nl = nl_MultLoop_acc_436_nl[24:0];
  assign nl_MultLoop_acc_3003_itm_1  = conv_s2s_16_17(MultLoop_acc_334_itm_20_5)
      + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_436_nl))) + conv_s2s_15_17(MultLoop_acc_434_itm_22_7[15:1]);
  assign nl_MultLoop_acc_2944_nl = (~ (data_rsci_idat[467:450])) + conv_s2s_14_18(data_rsci_idat[467:454]);
  assign MultLoop_acc_2944_nl = nl_MultLoop_acc_2944_nl[17:0];
  assign nl_MultLoop_acc_2945_nl = conv_s2s_20_21({(~ (data_rsci_idat[467:450]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2944_nl);
  assign MultLoop_acc_2945_nl = nl_MultLoop_acc_2945_nl[20:0];
  assign nl_MultLoop_acc_1233_nl = conv_s2u_21_22(MultLoop_acc_2945_nl) + ({(data_rsci_idat[467:450])
      , 4'b0100});
  assign MultLoop_acc_1233_nl = nl_MultLoop_acc_1233_nl[21:0];
  assign nl_MultLoop_acc_2947_nl = ({(data_rsci_idat[413:396]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_722_18_8
      , (~ (data_rsci_idat[403:396]))});
  assign MultLoop_acc_2947_nl = nl_MultLoop_acc_2947_nl[21:0];
  assign nl_MultLoop_acc_4333_nl = conv_s2u_14_18(readslicef_22_14_8((MultLoop_acc_2947_nl)))
      + (~ (data_rsci_idat[413:396]));
  assign MultLoop_acc_4333_nl = nl_MultLoop_acc_4333_nl[17:0];
  assign nl_MultLoop_acc_2937_nl = ({(data_rsci_idat[809:792]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_858_18_7
      , (~ (data_rsci_idat[798:792]))});
  assign MultLoop_acc_2937_nl = nl_MultLoop_acc_2937_nl[20:0];
  assign nl_MultLoop_acc_2938_nl = ({(~ (data_rsci_idat[809:792])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_2937_nl);
  assign MultLoop_acc_2938_nl = nl_MultLoop_acc_2938_nl[22:0];
  assign nl_MultLoop_acc_473_nl = conv_s2s_23_26(MultLoop_acc_2938_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[809:792])) , 7'b0100000});
  assign MultLoop_acc_473_nl = nl_MultLoop_acc_473_nl[25:0];
  assign nl_MultLoop_acc_2939_nl = (~ (data_rsci_idat[629:612])) + conv_s2s_16_18(data_rsci_idat[629:614]);
  assign MultLoop_acc_2939_nl = nl_MultLoop_acc_2939_nl[17:0];
  assign nl_MultLoop_acc_2940_nl = conv_s2s_21_22({(~ (data_rsci_idat[629:612]))
      , 3'b001}) + conv_s2s_18_22(MultLoop_acc_2939_nl);
  assign MultLoop_acc_2940_nl = nl_MultLoop_acc_2940_nl[21:0];
  assign nl_MultLoop_acc_1236_nl = conv_s2u_22_24(MultLoop_acc_2940_nl) + ({(data_rsci_idat[629:612])
      , 6'b001000});
  assign MultLoop_acc_1236_nl = nl_MultLoop_acc_1236_nl[23:0];
  assign nl_MultLoop_acc_2943_nl = conv_s2s_21_22({(data_rsci_idat[449:432]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[449:432]) + conv_s2s_16_22({MultLoop_acc_4186_cse_1
      , (data_rsci_idat[439:435])});
  assign MultLoop_acc_2943_nl = nl_MultLoop_acc_2943_nl[21:0];
  assign nl_MultLoop_acc_453_nl = conv_s2u_22_23(MultLoop_acc_2943_nl) + ({(~ (data_rsci_idat[449:432]))
      , 5'b00000});
  assign MultLoop_acc_453_nl = nl_MultLoop_acc_453_nl[22:0];
  assign nl_MultLoop_acc_452_nl = conv_s2u_15_18(data_rsci_idat[431:417]) - (data_rsci_idat[431:414]);
  assign MultLoop_acc_452_nl = nl_MultLoop_acc_452_nl[17:0];
  assign nl_MultLoop_acc_2948_nl = ({(data_rsci_idat[377:360]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[377:360]));
  assign MultLoop_acc_2948_nl = nl_MultLoop_acc_2948_nl[21:0];
  assign nl_MultLoop_acc_4334_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_2948_nl)))
      + conv_s2u_18_19(data_rsci_idat[377:360]);
  assign MultLoop_acc_4334_nl = nl_MultLoop_acc_4334_nl[18:0];
  assign nl_MultLoop_acc_3020_itm_1  = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1233_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4333_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_473_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1236_nl))) + conv_s2s_16_18(MultLoop_acc_1237_itm_20_4[16:1])
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_453_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_452_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4334_nl)));
  assign nl_MultLoop_acc_448_nl = conv_s2u_12_18(data_rsci_idat[359:348]) - (data_rsci_idat[359:342]);
  assign MultLoop_acc_448_nl = nl_MultLoop_acc_448_nl[17:0];
  assign nl_MultLoop_acc_445_nl = conv_s2s_25_26({(~ (data_rsci_idat[305:288])) ,
      7'b0001000}) + conv_s2s_21_26({(~ (data_rsci_idat[305:288])) , 3'b001}) + conv_s2s_19_26({MultLoop_MultLoop_conc_734_18_7
      , (~ (data_rsci_idat[294:288]))});
  assign MultLoop_acc_445_nl = nl_MultLoop_acc_445_nl[25:0];
  assign nl_MultLoop_acc_2952_nl = ({(~ (data_rsci_idat[269:252])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[269:252])
      + conv_s2s_15_20(data_rsci_idat[269:255]);
  assign MultLoop_acc_2952_nl = nl_MultLoop_acc_2952_nl[19:0];
  assign nl_MultLoop_acc_1232_nl = conv_s2u_20_23(MultLoop_acc_2952_nl) + ({(data_rsci_idat[269:252])
      , 5'b00100});
  assign MultLoop_acc_1232_nl = nl_MultLoop_acc_1232_nl[22:0];
  assign nl_MultLoop_acc_2954_nl = ({(data_rsci_idat[287:270]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_814_18_8
      , (~ (data_rsci_idat[277:270]))});
  assign MultLoop_acc_2954_nl = nl_MultLoop_acc_2954_nl[19:0];
  assign nl_MultLoop_acc_2955_nl = conv_s2s_24_25({(data_rsci_idat[287:270]) , 6'b000000})
      + conv_s2s_20_25(MultLoop_acc_2954_nl);
  assign MultLoop_acc_2955_nl = nl_MultLoop_acc_2955_nl[24:0];
  assign nl_MultLoop_acc_4337_nl = conv_s2u_17_18(readslicef_25_17_8((MultLoop_acc_2955_nl)))
      + (~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_4337_nl = nl_MultLoop_acc_4337_nl[17:0];
  assign nl_MultLoop_acc_3012_itm_1  = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_448_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_445_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1232_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4337_nl)));
  assign nl_MultLoop_acc_2958_nl = conv_s2s_21_22({(data_rsci_idat[233:216]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[233:216]) + conv_s2s_16_22({MultLoop_acc_3974_cse_1
      , (data_rsci_idat[223:219])});
  assign MultLoop_acc_2958_nl = nl_MultLoop_acc_2958_nl[21:0];
  assign nl_MultLoop_acc_441_nl = conv_s2u_22_23(MultLoop_acc_2958_nl) + ({(~ (data_rsci_idat[233:216]))
      , 5'b00000});
  assign MultLoop_acc_441_nl = nl_MultLoop_acc_441_nl[22:0];
  assign nl_MultLoop_acc_2961_nl = conv_s2s_20_21({(data_rsci_idat[89:72]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_1503_cse_1);
  assign MultLoop_acc_2961_nl = nl_MultLoop_acc_2961_nl[20:0];
  assign nl_MultLoop_acc_433_nl = conv_s2u_21_23(MultLoop_acc_2961_nl) + ({(~ (data_rsci_idat[89:72]))
      , 5'b00000});
  assign MultLoop_acc_433_nl = nl_MultLoop_acc_433_nl[22:0];
  assign nl_MultLoop_acc_2963_nl = ({(data_rsci_idat[71:54]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_758_18_6
      , (~ (data_rsci_idat[59:54]))});
  assign MultLoop_acc_2963_nl = nl_MultLoop_acc_2963_nl[20:0];
  assign nl_MultLoop_acc_4341_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_2963_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_4341_nl = nl_MultLoop_acc_4341_nl[17:0];
  assign nl_MultLoop_acc_4342_nl = conv_s2s_13_14(data_rsci_idat[683:671]) + 14'b00000000000001;
  assign MultLoop_acc_4342_nl = nl_MultLoop_acc_4342_nl[13:0];
  assign nl_MultLoop_acc_2904_nl = conv_s2s_18_19(data_rsci_idat[683:666]) + conv_s2s_16_19({(MultLoop_acc_4342_nl)
      , (data_rsci_idat[670:669])});
  assign MultLoop_acc_2904_nl = nl_MultLoop_acc_2904_nl[18:0];
  assign nl_MultLoop_acc_466_nl = conv_s2u_19_20(MultLoop_acc_2904_nl) + ({(~ (data_rsci_idat[683:666]))
      , 2'b00});
  assign MultLoop_acc_466_nl = nl_MultLoop_acc_466_nl[19:0];
  assign nl_MultLoop_acc_3011_itm_1  = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_441_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_433_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4341_nl)))
      + conv_s2s_13_18(MultLoop_acc_4590_itm_20_5[15:3]) + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_466_nl)))
      + conv_s2s_13_18(MultLoop_acc_447_itm_20_7[13:1]) + conv_s2s_12_18(MultLoop_acc_471_itm_21_7[14:3]);
  assign nl_MultLoop_acc_2551_nl = ({(~ (data_rsci_idat[341:324])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[341:324])
      + conv_s2s_16_20({MultLoop_acc_4122_cse_1 , (data_rsci_idat[331:327])});
  assign MultLoop_acc_2551_nl = nl_MultLoop_acc_2551_nl[19:0];
  assign nl_MultLoop_acc_1293_nl = conv_s2u_20_24(MultLoop_acc_2551_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[341:324])) , 5'b00100});
  assign MultLoop_acc_1293_nl = nl_MultLoop_acc_1293_nl[23:0];
  assign nl_MultLoop_acc_2554_nl = ({(~ (data_rsci_idat[269:252])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[269:252])
      + conv_s2s_16_21({MultLoop_acc_4150_cse_1 , (data_rsci_idat[259:255])});
  assign MultLoop_acc_2554_nl = nl_MultLoop_acc_2554_nl[20:0];
  assign nl_MultLoop_acc_1292_nl = conv_s2u_21_24(MultLoop_acc_2554_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[269:252])) , 5'b01000});
  assign MultLoop_acc_1292_nl = nl_MultLoop_acc_1292_nl[23:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_222_itm_1 
      = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1293_nl))) + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1292_nl)));
  assign nl_MultLoop_acc_2557_nl = ({(~ (data_rsci_idat[197:180])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[197:180])
      + conv_s2s_16_20({MultLoop_acc_4191_cse_1 , (data_rsci_idat[187:183])});
  assign MultLoop_acc_2557_nl = nl_MultLoop_acc_2557_nl[19:0];
  assign nl_MultLoop_acc_1291_nl = conv_s2u_20_24(MultLoop_acc_2557_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[197:180])) , 5'b00100});
  assign MultLoop_acc_1291_nl = nl_MultLoop_acc_1291_nl[23:0];
  assign nl_MultLoop_acc_4192_nl = conv_s2s_13_14(data_rsci_idat[791:779]) + 14'b00000000000001;
  assign MultLoop_acc_4192_nl = nl_MultLoop_acc_4192_nl[13:0];
  assign nl_MultLoop_acc_2480_nl = conv_s2s_18_19(data_rsci_idat[791:774]) + conv_s2s_17_19({(MultLoop_acc_4192_nl)
      , (data_rsci_idat[778:776])});
  assign MultLoop_acc_2480_nl = nl_MultLoop_acc_2480_nl[18:0];
  assign nl_MultLoop_acc_659_nl = conv_s2u_19_21(MultLoop_acc_2480_nl) + ({(~ (data_rsci_idat[791:774]))
      , 3'b000});
  assign MultLoop_acc_659_nl = nl_MultLoop_acc_659_nl[20:0];
  assign nl_MultLoop_acc_2481_nl = ({(data_rsci_idat[701:684]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[701:684]));
  assign MultLoop_acc_2481_nl = nl_MultLoop_acc_2481_nl[20:0];
  assign nl_MultLoop_acc_654_nl = conv_s2s_21_24(MultLoop_acc_2481_nl) + conv_s2s_23_24({(data_rsci_idat[701:684])
      , 5'b00000});
  assign MultLoop_acc_654_nl = nl_MultLoop_acc_654_nl[23:0];
  assign nl_MultLoop_acc_2483_nl = (~ (data_rsci_idat[719:702])) + conv_s2s_17_18({MultLoop_acc_3916_cse_1
      , (data_rsci_idat[707:704])});
  assign MultLoop_acc_2483_nl = nl_MultLoop_acc_2483_nl[17:0];
  assign nl_MultLoop_acc_2484_nl = ({(data_rsci_idat[719:702]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2483_nl);
  assign MultLoop_acc_2484_nl = nl_MultLoop_acc_2484_nl[19:0];
  assign nl_MultLoop_acc_655_nl = conv_s2u_20_22(MultLoop_acc_2484_nl) + ({(~ (data_rsci_idat[719:702]))
      , 4'b0000});
  assign MultLoop_acc_655_nl = nl_MultLoop_acc_655_nl[21:0];
  assign nl_MultLoop_acc_4194_nl =  -conv_s2s_14_15(data_rsci_idat[521:508]);
  assign MultLoop_acc_4194_nl = nl_MultLoop_acc_4194_nl[14:0];
  assign nl_MultLoop_acc_644_nl = conv_s2s_19_23({(MultLoop_acc_4194_nl) , (~ (data_rsci_idat[507:504]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[521:504])) , 4'b0001});
  assign MultLoop_acc_644_nl = nl_MultLoop_acc_644_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl = conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_659_nl)))
      + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_654_nl))) + conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_655_nl)))
      + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_644_nl)));
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl[15:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_221_itm_1_16_0
      = (readslicef_24_17_7((MultLoop_acc_1291_nl))) + conv_s2s_16_17(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_208_nl);
  assign nl_MultLoop_acc_645_nl = conv_s2u_12_18(data_rsci_idat[539:528]) - (data_rsci_idat[539:522]);
  assign MultLoop_acc_645_nl = nl_MultLoop_acc_645_nl[17:0];
  assign nl_MultLoop_acc_4195_nl =  -conv_s2s_14_15(data_rsci_idat[431:418]);
  assign MultLoop_acc_4195_nl = nl_MultLoop_acc_4195_nl[14:0];
  assign nl_MultLoop_acc_639_nl = conv_s2s_19_23({(MultLoop_acc_4195_nl) , (~ (data_rsci_idat[417:414]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[431:414])) , 4'b0001});
  assign MultLoop_acc_639_nl = nl_MultLoop_acc_639_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_207_itm_1 
      = conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_645_nl))) + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_639_nl)))
      + conv_s2s_14_16(MultLoop_acc_1128_itm_21_7[14:1]) + conv_s2s_14_16(MultLoop_acc_150_itm_17_4);
  assign nl_MultLoop_acc_1301_nl = conv_s2u_14_19(data_rsci_idat[845:832]) + conv_s2u_18_19(data_rsci_idat[845:828]);
  assign MultLoop_acc_1301_nl = nl_MultLoop_acc_1301_nl[18:0];
  assign nl_MultLoop_acc_4672_nl = conv_s2u_19_23(MultLoop_acc_2030_cse_1[20:2])
      + conv_s2u_22_23({(~ (data_rsci_idat[809:792])) , 4'b0001});
  assign MultLoop_acc_4672_nl = nl_MultLoop_acc_4672_nl[22:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_206_itm_1 
      = conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_1301_nl))) + conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_4672_nl)));
  assign nl_MultLoop_acc_4197_nl = conv_s2s_11_12(data_rsci_idat[755:745]) + 12'b000000000001;
  assign MultLoop_acc_4197_nl = nl_MultLoop_acc_4197_nl[11:0];
  assign nl_MultLoop_acc_2491_nl = conv_s2s_21_22({(data_rsci_idat[755:738]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[755:738]) + conv_s2s_17_22({(MultLoop_acc_4197_nl)
      , (data_rsci_idat[744:740])});
  assign MultLoop_acc_2491_nl = nl_MultLoop_acc_2491_nl[21:0];
  assign nl_MultLoop_acc_657_nl = conv_s2u_22_23(MultLoop_acc_2491_nl) + ({(~ (data_rsci_idat[755:738]))
      , 5'b00000});
  assign MultLoop_acc_657_nl = nl_MultLoop_acc_657_nl[22:0];
  assign nl_MultLoop_acc_4673_nl = conv_s2u_18_21(MultLoop_asn_1479) + ({(data_rsci_idat[683:666])
      , 3'b001});
  assign MultLoop_acc_4673_nl = nl_MultLoop_acc_4673_nl[20:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_205_itm_1 
      = conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_657_nl))) + conv_s2s_15_16(readslicef_21_15_6((MultLoop_acc_4673_nl)));
  assign nl_MultLoop_acc_2495_nl = conv_s2s_23_24({(~ (data_rsci_idat[611:594]))
      , 5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[611:594])) , 3'b001}) + conv_s2s_18_24(~
      (data_rsci_idat[611:594]));
  assign MultLoop_acc_2495_nl = nl_MultLoop_acc_2495_nl[23:0];
  assign nl_MultLoop_acc_649_nl = conv_s2s_24_25(MultLoop_acc_2495_nl) + ({(data_rsci_idat[611:594])
      , 7'b0100000});
  assign MultLoop_acc_649_nl = nl_MultLoop_acc_649_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_204_itm_1 
      = conv_s2s_15_16(MultLoop_acc_1097_itm_18_4) + conv_s2s_15_16(readslicef_25_15_10((MultLoop_acc_649_nl)));
  assign nl_MultLoop_acc_643_nl = conv_s2s_24_25({(~ (data_rsci_idat[503:486])) ,
      6'b000100}) + conv_s2s_20_25({(~ (data_rsci_idat[503:486])) , 2'b01}) + conv_s2s_19_25({MultLoop_MultLoop_conc_742_18_6
      , (~ (data_rsci_idat[491:486]))});
  assign MultLoop_acc_643_nl = nl_MultLoop_acc_643_nl[24:0];
  assign nl_MultLoop_acc_2499_nl = conv_s2s_21_22({(~ (data_rsci_idat[413:396]))
      , 3'b001}) + conv_s2s_18_22(MultLoop_acc_2403_cse_1);
  assign MultLoop_acc_2499_nl = nl_MultLoop_acc_2499_nl[21:0];
  assign nl_MultLoop_acc_1296_nl = conv_s2u_22_23(MultLoop_acc_2499_nl) + ({(data_rsci_idat[413:396])
      , 5'b01000});
  assign MultLoop_acc_1296_nl = nl_MultLoop_acc_1296_nl[22:0];
  assign nl_MultLoop_acc_2501_nl = ({(~ (data_rsci_idat[377:360])) , 3'b000}) + conv_s2s_19_21(MultLoop_acc_2500_cse_1);
  assign MultLoop_acc_2501_nl = nl_MultLoop_acc_2501_nl[20:0];
  assign nl_MultLoop_acc_1295_nl = conv_s2u_21_23(MultLoop_acc_2501_nl) + ({(data_rsci_idat[377:360])
      , 5'b01000});
  assign MultLoop_acc_1295_nl = nl_MultLoop_acc_1295_nl[22:0];
  assign nl_MultLoop_acc_2503_nl = conv_s2s_22_23({(~ (data_rsci_idat[395:378]))
      , 4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[395:378])) , 2'b01}) + conv_s2s_18_23(~
      (data_rsci_idat[395:378]));
  assign MultLoop_acc_2503_nl = nl_MultLoop_acc_2503_nl[22:0];
  assign nl_MultLoop_acc_637_nl = conv_s2s_23_25(MultLoop_acc_2503_nl) + ({(data_rsci_idat[395:378])
      , 7'b0010000});
  assign MultLoop_acc_637_nl = nl_MultLoop_acc_637_nl[24:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_218_itm_1 
      = conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_643_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1296_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1295_nl))) + conv_s2s_15_17(readslicef_25_15_10((MultLoop_acc_637_nl)));
  assign nl_MultLoop_acc_2505_nl = conv_s2s_18_19(data_rsci_idat[305:288]) + conv_s2s_17_19({MultLoop_MultLoop_conc_706_16_4
      , (data_rsci_idat[293:290])});
  assign MultLoop_acc_2505_nl = nl_MultLoop_acc_2505_nl[18:0];
  assign nl_MultLoop_acc_632_nl = conv_s2u_19_22(MultLoop_acc_2505_nl) + ({(~ (data_rsci_idat[305:288]))
      , 4'b0000});
  assign MultLoop_acc_632_nl = nl_MultLoop_acc_632_nl[21:0];
  assign nl_MultLoop_acc_2507_nl = (~ (data_rsci_idat[125:108])) + conv_s2s_17_18({Result_acc_187_cse_1
      , (data_rsci_idat[114:110])});
  assign MultLoop_acc_2507_nl = nl_MultLoop_acc_2507_nl[17:0];
  assign nl_MultLoop_acc_2508_nl = ({(data_rsci_idat[125:108]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_2507_nl);
  assign MultLoop_acc_2508_nl = nl_MultLoop_acc_2508_nl[20:0];
  assign nl_MultLoop_acc_622_nl = conv_s2u_21_23(MultLoop_acc_2508_nl) + ({(~ (data_rsci_idat[125:108]))
      , 5'b00000});
  assign MultLoop_acc_622_nl = nl_MultLoop_acc_622_nl[22:0];
  assign nl_MultLoop_acc_2509_nl = conv_s2s_18_19(data_rsci_idat[143:126]) + conv_s2s_14_19(data_rsci_idat[143:130]);
  assign MultLoop_acc_2509_nl = nl_MultLoop_acc_2509_nl[18:0];
  assign nl_MultLoop_acc_1289_nl = conv_s2u_19_21(MultLoop_acc_2509_nl) + conv_s2u_20_21({(data_rsci_idat[143:126])
      , 2'b00});
  assign MultLoop_acc_1289_nl = nl_MultLoop_acc_1289_nl[20:0];
  assign nl_MultLoop_acc_4201_nl =  -conv_s2s_12_13(data_rsci_idat[53:42]);
  assign MultLoop_acc_4201_nl = nl_MultLoop_acc_4201_nl[12:0];
  assign nl_MultLoop_acc_2512_nl = ({(data_rsci_idat[53:36]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[53:36])) , 2'b01}) + conv_s2s_19_22({(MultLoop_acc_4201_nl)
      , (~ (data_rsci_idat[41:36]))});
  assign MultLoop_acc_2512_nl = nl_MultLoop_acc_2512_nl[21:0];
  assign nl_MultLoop_acc_4202_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2512_nl)))
      + (~ (data_rsci_idat[53:36]));
  assign MultLoop_acc_4202_nl = nl_MultLoop_acc_4202_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_217_itm_1 
      = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_632_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_622_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1289_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4202_nl)));
  assign nl_MultLoop_acc_2514_nl = ({(data_rsci_idat[71:54]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_786_18_7
      , (~ (data_rsci_idat[60:54]))});
  assign MultLoop_acc_2514_nl = nl_MultLoop_acc_2514_nl[20:0];
  assign nl_MultLoop_acc_2515_nl = conv_s2s_23_24({(data_rsci_idat[71:54]) , 5'b00000})
      + conv_s2s_21_24(MultLoop_acc_2514_nl);
  assign MultLoop_acc_2515_nl = nl_MultLoop_acc_2515_nl[23:0];
  assign nl_MultLoop_acc_4204_nl = conv_s2u_17_18(readslicef_24_17_7((MultLoop_acc_2515_nl)))
      + (~ (data_rsci_idat[71:54]));
  assign MultLoop_acc_4204_nl = nl_MultLoop_acc_4204_nl[17:0];
  assign nl_MultLoop_acc_2518_nl = conv_s2s_20_21({(data_rsci_idat[17:0]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_1531_cse_1);
  assign MultLoop_acc_2518_nl = nl_MultLoop_acc_2518_nl[20:0];
  assign nl_MultLoop_acc_616_nl = conv_s2u_21_23(MultLoop_acc_2518_nl) + ({(~ (data_rsci_idat[17:0]))
      , 5'b00000});
  assign MultLoop_acc_616_nl = nl_MultLoop_acc_616_nl[22:0];
  assign nl_MultLoop_625_MultLoop_acc_3_nl = (readslicef_23_15_8((MultLoop_acc_616_nl)))
      + 15'b000001000110111;
  assign MultLoop_625_MultLoop_acc_3_nl = nl_MultLoop_625_MultLoop_acc_3_nl[14:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_199_itm_1 
      = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4204_nl))) + conv_s2s_15_16(MultLoop_625_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_4674_nl = conv_s2u_18_19(data_rsci_idat[773:756]) + conv_s2u_14_19(MultLoop_acc_2520_cse_1[19:6]);
  assign MultLoop_acc_4674_nl = nl_MultLoop_acc_4674_nl[18:0];
  assign nl_MultLoop_acc_4207_nl = conv_s2u_17_18(readslicef_19_17_2((MultLoop_acc_4674_nl)))
      + (~ (data_rsci_idat[773:756]));
  assign MultLoop_acc_4207_nl = nl_MultLoop_acc_4207_nl[17:0];
  assign nl_MultLoop_acc_2523_nl = conv_s2s_20_21({(data_rsci_idat[737:720]) , 2'b00})
      + conv_s2s_19_21(MultLoop_acc_2522_cse_1);
  assign MultLoop_acc_2523_nl = nl_MultLoop_acc_2523_nl[20:0];
  assign nl_MultLoop_acc_1300_nl = conv_s2u_21_23(MultLoop_acc_2523_nl) + conv_s2u_22_23({(data_rsci_idat[737:720])
      , 4'b0000});
  assign MultLoop_acc_1300_nl = nl_MultLoop_acc_1300_nl[22:0];
  assign nl_MultLoop_acc_2526_nl = ({(~ (data_rsci_idat[629:612])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2525_cse_1);
  assign MultLoop_acc_2526_nl = nl_MultLoop_acc_2526_nl[19:0];
  assign nl_MultLoop_acc_2527_nl = ({(data_rsci_idat[629:612]) , 4'b0100}) + conv_s2s_20_22(MultLoop_acc_2526_nl);
  assign MultLoop_acc_2527_nl = nl_MultLoop_acc_2527_nl[21:0];
  assign nl_MultLoop_acc_4209_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2527_nl)))
      + (~ (data_rsci_idat[629:612]));
  assign MultLoop_acc_4209_nl = nl_MultLoop_acc_4209_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_215_itm_1 
      = conv_s2s_16_17(readslicef_23_16_7((MultLoop_acc_1300_nl))) + conv_s2s_16_17(readslicef_18_16_2((MultLoop_acc_4209_nl)));
  assign nl_MultLoop_acc_2537_nl = conv_s2s_18_19(data_rsci_idat[449:432]) + conv_s2s_16_19(data_rsci_idat[449:434]);
  assign MultLoop_acc_2537_nl = nl_MultLoop_acc_2537_nl[18:0];
  assign nl_MultLoop_acc_1297_nl = conv_s2u_19_22(MultLoop_acc_2537_nl) + conv_s2u_21_22({(data_rsci_idat[449:432])
      , 3'b000});
  assign MultLoop_acc_1297_nl = nl_MultLoop_acc_1297_nl[21:0];
  assign nl_MultLoop_acc_641_nl = conv_s2u_12_18(data_rsci_idat[467:456]) - (data_rsci_idat[467:450]);
  assign MultLoop_acc_641_nl = nl_MultLoop_acc_641_nl[17:0];
  assign nl_MultLoop_acc_651_nl = conv_s2s_23_24({(~ (data_rsci_idat[647:630])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[647:630])) , 3'b001}) + conv_s2s_19_24({MultLoop_MultLoop_conc_834_18_5
      , (~ (data_rsci_idat[634:630]))});
  assign MultLoop_acc_651_nl = nl_MultLoop_acc_651_nl[23:0];
  assign nl_MultLoop_acc_4211_nl =  -conv_s2s_13_14(data_rsci_idat[557:545]);
  assign MultLoop_acc_4211_nl = nl_MultLoop_acc_4211_nl[13:0];
  assign nl_MultLoop_acc_646_nl = conv_s2s_23_24({(~ (data_rsci_idat[557:540])) ,
      5'b01000}) + conv_s2s_21_24({(~ (data_rsci_idat[557:540])) , 3'b001}) + conv_s2s_19_24({(MultLoop_acc_4211_nl)
      , (~ (data_rsci_idat[544:540]))});
  assign MultLoop_acc_646_nl = nl_MultLoop_acc_646_nl[23:0];
  assign nl_MultLoop_acc_2533_nl = (~ (data_rsci_idat[575:558])) + conv_s2s_16_18({MultLoop_acc_4212_cse_1
      , (data_rsci_idat[565:561])});
  assign MultLoop_acc_2533_nl = nl_MultLoop_acc_2533_nl[17:0];
  assign nl_MultLoop_acc_2534_nl = ({(data_rsci_idat[575:558]) , 3'b001}) + conv_s2s_18_21(MultLoop_acc_2533_nl);
  assign MultLoop_acc_2534_nl = nl_MultLoop_acc_2534_nl[20:0];
  assign nl_MultLoop_acc_647_nl = conv_s2u_21_23(MultLoop_acc_2534_nl) + ({(~ (data_rsci_idat[575:558]))
      , 5'b00000});
  assign MultLoop_acc_647_nl = nl_MultLoop_acc_647_nl[22:0];
  assign nl_MultLoop_acc_2536_nl = conv_s2s_21_22({(~ (data_rsci_idat[485:468]))
      , 3'b001}) + conv_s2s_18_22(MultLoop_acc_2535_cse_1);
  assign MultLoop_acc_2536_nl = nl_MultLoop_acc_2536_nl[21:0];
  assign nl_MultLoop_acc_1298_nl = conv_s2u_22_23(MultLoop_acc_2536_nl) + ({(data_rsci_idat[485:468])
      , 5'b01000});
  assign MultLoop_acc_1298_nl = nl_MultLoop_acc_1298_nl[22:0];
  assign nl_MultLoop_acc_2540_nl = ({(data_rsci_idat[323:306]) , 6'b000100}) + conv_s2s_20_24({(~
      (data_rsci_idat[323:306])) , 2'b01}) + conv_s2s_19_24({MultLoop_MultLoop_conc_836_18_8
      , (~ (data_rsci_idat[313:306]))});
  assign MultLoop_acc_2540_nl = nl_MultLoop_acc_2540_nl[23:0];
  assign nl_MultLoop_acc_4214_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_2540_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_4214_nl = nl_MultLoop_acc_4214_nl[17:0];
  assign nl_MultLoop_acc_629_nl = conv_s2u_14_18(data_rsci_idat[251:238]) - (data_rsci_idat[251:234]);
  assign MultLoop_acc_629_nl = nl_MultLoop_acc_629_nl[17:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_232_itm_1 
      = conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1297_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_641_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_651_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_646_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_647_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1298_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4214_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_629_nl)));
  assign nl_MultLoop_acc_2542_nl = ({(~ (data_rsci_idat[161:144])) , 3'b000}) + conv_s2s_18_21(data_rsci_idat[161:144])
      + conv_s2s_15_21(data_rsci_idat[161:147]);
  assign MultLoop_acc_2542_nl = nl_MultLoop_acc_2542_nl[20:0];
  assign nl_MultLoop_acc_1290_nl = conv_s2u_21_23(MultLoop_acc_2542_nl) + ({(data_rsci_idat[161:144])
      , 5'b01000});
  assign MultLoop_acc_1290_nl = nl_MultLoop_acc_1290_nl[22:0];
  assign nl_MultLoop_acc_2544_nl = ({(data_rsci_idat[179:162]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_826_18_5
      , (~ (data_rsci_idat[166:162]))});
  assign MultLoop_acc_2544_nl = nl_MultLoop_acc_2544_nl[19:0];
  assign nl_MultLoop_acc_625_nl = conv_s2s_20_23(MultLoop_acc_2544_nl) + ({(~ (data_rsci_idat[179:162]))
      , 5'b00000});
  assign MultLoop_acc_625_nl = nl_MultLoop_acc_625_nl[22:0];
  assign nl_MultLoop_acc_4624_nl = conv_s2u_19_24(MultLoop_acc_1485_cse_1[20:2])
      + ({(data_rsci_idat[89:72]) , 6'b000001});
  assign MultLoop_acc_4624_nl = nl_MultLoop_acc_4624_nl[23:0];
  assign nl_MultLoop_acc_631_nl = conv_s2u_14_18(data_rsci_idat[287:274]) - (data_rsci_idat[287:270]);
  assign MultLoop_acc_631_nl = nl_MultLoop_acc_631_nl[17:0];
  assign nl_MultLoop_acc_4216_nl = conv_s2s_14_15(data_rsci_idat[233:220]) + 15'b000000000000001;
  assign MultLoop_acc_4216_nl = nl_MultLoop_acc_4216_nl[14:0];
  assign nl_MultLoop_acc_2478_nl = conv_s2s_18_19(data_rsci_idat[233:216]) + conv_s2s_17_19({(MultLoop_acc_4216_nl)
      , (data_rsci_idat[219:218])});
  assign MultLoop_acc_2478_nl = nl_MultLoop_acc_2478_nl[18:0];
  assign nl_MultLoop_acc_628_nl = conv_s2u_19_20(MultLoop_acc_2478_nl) + ({(~ (data_rsci_idat[233:216]))
      , 2'b00});
  assign MultLoop_acc_628_nl = nl_MultLoop_acc_628_nl[19:0];
  assign nl_MultLoop_acc_627_nl = conv_s2u_16_18(data_rsci_idat[215:200]) - (data_rsci_idat[215:198]);
  assign MultLoop_acc_627_nl = nl_MultLoop_acc_627_nl[17:0];
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl = ~((data_rsci_idat[816:810]!=7'b0000000));
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl = conv_s2s_11_12(~
      (data_rsci_idat[827:817])) + conv_s2s_11_12(readslicef_18_11_7((MultLoop_acc_627_nl)))
      + conv_u2s_1_12(nnet_product_input_t_config2_weight_t_config2_accum_t_nor_4_nl);
  assign nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl = nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl[11:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_224_itm_1 
      = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1290_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_625_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_4624_nl))) + conv_s2s_13_18(readslicef_18_13_5((MultLoop_acc_631_nl)))
      + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_628_nl))) + conv_s2s_13_18(MultLoop_acc_1741_cse_1[18:6])
      + conv_s2s_12_18(nnet_product_input_t_config2_weight_t_config2_accum_t_acc_191_nl);
  assign nl_MultLoop_acc_2547_nl = (~ (data_rsci_idat[863:846])) + conv_s2s_17_18({MultLoop_acc_4011_cse_1
      , (data_rsci_idat[853:848])});
  assign MultLoop_acc_2547_nl = nl_MultLoop_acc_2547_nl[17:0];
  assign nl_MultLoop_acc_1302_nl = conv_s2u_18_25(MultLoop_acc_2547_nl) + conv_s2u_24_25({(~
      (data_rsci_idat[863:846])) , 6'b000001});
  assign MultLoop_acc_1302_nl = nl_MultLoop_acc_1302_nl[24:0];
  assign nl_MultLoop_acc_4218_nl = conv_s2u_13_19(MultLoop_acc_1743_cse_1[20:8])
      + conv_s2u_18_19(data_rsci_idat[665:648]);
  assign MultLoop_acc_4218_nl = nl_MultLoop_acc_4218_nl[18:0];
  assign nl_nnet_product_input_t_config2_weight_t_config2_accum_t_acc_223_itm_1 
      = conv_s2s_17_18(readslicef_25_17_8((MultLoop_acc_1302_nl))) + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4218_nl)));
  assign nl_MultLoop_acc_2849_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_16_18({MultLoop_acc_4076_cse_1
      , (data_rsci_idat[743:741])});
  assign MultLoop_acc_2849_nl = nl_MultLoop_acc_2849_nl[17:0];
  assign nl_MultLoop_acc_1251_nl = conv_s2u_18_22(MultLoop_acc_2849_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[755:738])) , 3'b001});
  assign MultLoop_acc_1251_nl = nl_MultLoop_acc_1251_nl[21:0];
  assign nl_MultLoop_acc_2843_nl = conv_s2s_18_19(data_rsci_idat[107:90]) + conv_s2s_16_19({MultLoop_MultLoop_conc_694_15_3
      , (data_rsci_idat[95:93])});
  assign MultLoop_acc_2843_nl = nl_MultLoop_acc_2843_nl[18:0];
  assign nl_MultLoop_acc_482_nl = conv_s2u_19_21(MultLoop_acc_2843_nl) + ({(~ (data_rsci_idat[107:90]))
      , 3'b000});
  assign MultLoop_acc_482_nl = nl_MultLoop_acc_482_nl[20:0];
  assign nl_MultLoop_acc_1239_nl = conv_s2u_16_19(data_rsci_idat[35:20]) + conv_s2u_18_19(data_rsci_idat[35:18]);
  assign MultLoop_acc_1239_nl = nl_MultLoop_acc_1239_nl[18:0];
  assign nl_MultLoop_acc_2847_nl = (readslicef_19_14_5((MultLoop_acc_1239_nl))) +
      14'b00001000110001;
  assign MultLoop_acc_2847_nl = nl_MultLoop_acc_2847_nl[13:0];
  assign nl_MultLoop_acc_2846_nl = conv_s2s_21_22({(data_rsci_idat[17:0]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[17:0]) + conv_s2s_16_22({MultLoop_acc_4015_cse_1
      , (data_rsci_idat[7:3])});
  assign MultLoop_acc_2846_nl = nl_MultLoop_acc_2846_nl[21:0];
  assign nl_MultLoop_acc_477_nl = conv_s2u_22_23(MultLoop_acc_2846_nl) + ({(~ (data_rsci_idat[17:0]))
      , 5'b00000});
  assign MultLoop_acc_477_nl = nl_MultLoop_acc_477_nl[22:0];
  assign nl_MultLoop_482_MultLoop_acc_3_nl = conv_s2s_14_16(MultLoop_acc_2847_nl)
      + (readslicef_23_16_7((MultLoop_acc_477_nl)));
  assign MultLoop_482_MultLoop_acc_3_nl = nl_MultLoop_482_MultLoop_acc_3_nl[15:0];
  assign nl_MultLoop_acc_2888_itm_1  = conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1251_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_482_nl))) + conv_s2s_16_18(MultLoop_482_MultLoop_acc_3_nl);
  assign nl_MultLoop_acc_2851_nl = ({(data_rsci_idat[521:504]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_726_18_7
      , (~ (data_rsci_idat[510:504]))});
  assign MultLoop_acc_2851_nl = nl_MultLoop_acc_2851_nl[20:0];
  assign nl_MultLoop_acc_2852_nl = ({(~ (data_rsci_idat[521:504])) , 5'b00000}) +
      conv_s2s_21_23(MultLoop_acc_2851_nl);
  assign MultLoop_acc_2852_nl = nl_MultLoop_acc_2852_nl[22:0];
  assign nl_MultLoop_acc_505_nl = conv_s2s_23_26(MultLoop_acc_2852_nl) + conv_s2s_25_26({(~
      (data_rsci_idat[521:504])) , 7'b0100000});
  assign MultLoop_acc_505_nl = nl_MultLoop_acc_505_nl[25:0];
  assign nl_MultLoop_acc_4280_nl =  -conv_s2s_13_14(data_rsci_idat[503:491]);
  assign MultLoop_acc_4280_nl = nl_MultLoop_acc_4280_nl[13:0];
  assign nl_MultLoop_acc_504_nl = conv_s2s_23_24({(~ (data_rsci_idat[503:486])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[503:486])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4280_nl)
      , (~ (data_rsci_idat[490:486]))});
  assign MultLoop_acc_504_nl = nl_MultLoop_acc_504_nl[23:0];
  assign nl_MultLoop_acc_2887_itm_1  = conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_505_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_504_nl)));
  assign nl_MultLoop_acc_4281_nl = conv_s2s_10_11(data_rsci_idat[359:350]) + 11'b00000000001;
  assign MultLoop_acc_4281_nl = nl_MultLoop_acc_4281_nl[10:0];
  assign nl_MultLoop_acc_2856_nl = (~ (data_rsci_idat[359:342])) + conv_s2s_13_18({(MultLoop_acc_4281_nl)
      , (data_rsci_idat[349:348])});
  assign MultLoop_acc_2856_nl = nl_MultLoop_acc_2856_nl[17:0];
  assign nl_MultLoop_acc_1245_nl = conv_s2u_18_21(MultLoop_acc_2856_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[359:342])) , 2'b01});
  assign MultLoop_acc_1245_nl = nl_MultLoop_acc_1245_nl[20:0];
  assign nl_MultLoop_acc_4282_nl = conv_s2s_14_15(data_rsci_idat[125:112]) + 15'b000000000000001;
  assign MultLoop_acc_4282_nl = nl_MultLoop_acc_4282_nl[14:0];
  assign nl_MultLoop_acc_2858_nl = conv_s2s_18_19(data_rsci_idat[125:108]) + conv_s2s_17_19({(MultLoop_acc_4282_nl)
      , (data_rsci_idat[111:110])});
  assign MultLoop_acc_2858_nl = nl_MultLoop_acc_2858_nl[18:0];
  assign nl_MultLoop_acc_483_nl = conv_s2u_19_20(MultLoop_acc_2858_nl) + ({(~ (data_rsci_idat[125:108]))
      , 2'b00});
  assign MultLoop_acc_483_nl = nl_MultLoop_acc_483_nl[19:0];
  assign nl_MultLoop_acc_2886_itm_1  = conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1245_nl)))
      + conv_s2s_17_18(readslicef_20_17_3((MultLoop_acc_483_nl)));
  assign nl_MultLoop_acc_4285_nl = conv_s2s_12_13(data_rsci_idat[431:420]) + 13'b0000000000001;
  assign MultLoop_acc_4285_nl = nl_MultLoop_acc_4285_nl[12:0];
  assign nl_MultLoop_acc_2786_nl = (~ (data_rsci_idat[431:414])) + conv_s2s_17_18({(MultLoop_acc_4285_nl)
      , (data_rsci_idat[419:416])});
  assign MultLoop_acc_2786_nl = nl_MultLoop_acc_2786_nl[17:0];
  assign nl_MultLoop_acc_2787_nl = ({(data_rsci_idat[431:414]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2786_nl);
  assign MultLoop_acc_2787_nl = nl_MultLoop_acc_2787_nl[19:0];
  assign nl_MultLoop_acc_500_nl = conv_s2u_20_22(MultLoop_acc_2787_nl) + ({(~ (data_rsci_idat[431:414]))
      , 4'b0000});
  assign MultLoop_acc_500_nl = nl_MultLoop_acc_500_nl[21:0];
  assign nl_MultLoop_acc_2789_nl = ({(data_rsci_idat[143:126]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_824_18_6
      , (~ (data_rsci_idat[131:126]))});
  assign MultLoop_acc_2789_nl = nl_MultLoop_acc_2789_nl[19:0];
  assign nl_MultLoop_acc_4287_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_2789_nl)))
      + (~ (data_rsci_idat[143:126]));
  assign MultLoop_acc_4287_nl = nl_MultLoop_acc_4287_nl[17:0];
  assign nl_MultLoop_acc_4283_nl =  -conv_s2s_16_17(data_rsci_idat[197:182]);
  assign MultLoop_acc_4283_nl = nl_MultLoop_acc_4283_nl[16:0];
  assign nl_MultLoop_acc_487_nl = conv_s2s_19_21({(MultLoop_acc_4283_nl) , (~ (data_rsci_idat[181:180]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[197:180])) , 2'b01});
  assign MultLoop_acc_487_nl = nl_MultLoop_acc_487_nl[20:0];
  assign nl_MultLoop_acc_4284_nl =  -conv_s2s_16_17(data_rsci_idat[341:326]);
  assign MultLoop_acc_4284_nl = nl_MultLoop_acc_4284_nl[16:0];
  assign nl_MultLoop_acc_495_nl = conv_s2s_19_21({(MultLoop_acc_4284_nl) , (~ (data_rsci_idat[325:324]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[341:324])) , 2'b01});
  assign MultLoop_acc_495_nl = nl_MultLoop_acc_495_nl[20:0];
  assign nl_MultLoop_acc_2860_nl = (readslicef_21_12_9((MultLoop_acc_495_nl))) +
      conv_s2s_10_12(MultLoop_acc_506_itm_17_5[12:3]) + conv_s2s_9_12(data_rsci_idat[665:657]);
  assign MultLoop_acc_2860_nl = nl_MultLoop_acc_2860_nl[11:0];
  assign nl_MultLoop_acc_2871_itm_1  = conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_500_nl)))
      + conv_s2s_14_16(MultLoop_acc_1243_itm_19_6) + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4287_nl)))
      + conv_s2s_13_16(readslicef_21_13_8((MultLoop_acc_487_nl))) + conv_s2s_12_16(MultLoop_acc_2860_nl);
  assign nl_MultLoop_acc_518_nl = conv_s2s_23_24({(~ (data_rsci_idat[773:756])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[773:756])) , 2'b01}) + conv_s2s_19_24({MultLoop_MultLoop_conc_760_18_5
      , (~ (data_rsci_idat[760:756]))});
  assign MultLoop_acc_518_nl = nl_MultLoop_acc_518_nl[23:0];
  assign nl_MultLoop_acc_2793_nl = (~ (data_rsci_idat[791:774])) + conv_s2s_16_18({MultLoop_acc_4083_cse_1
      , (data_rsci_idat[780:777])});
  assign MultLoop_acc_2793_nl = nl_MultLoop_acc_2793_nl[17:0];
  assign nl_MultLoop_acc_2794_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2793_nl);
  assign MultLoop_acc_2794_nl = nl_MultLoop_acc_2794_nl[19:0];
  assign nl_MultLoop_acc_519_nl = conv_s2u_20_22(MultLoop_acc_2794_nl) + ({(~ (data_rsci_idat[791:774]))
      , 4'b0000});
  assign MultLoop_acc_519_nl = nl_MultLoop_acc_519_nl[21:0];
  assign nl_MultLoop_acc_2870_itm_1  = conv_s2s_15_16(readslicef_24_15_9((MultLoop_acc_518_nl)))
      + conv_s2s_15_16(readslicef_22_15_7((MultLoop_acc_519_nl)));
  assign nl_MultLoop_acc_2795_nl = conv_s2s_18_19(data_rsci_idat[575:558]) + conv_s2s_14_19(data_rsci_idat[575:562]);
  assign MultLoop_acc_2795_nl = nl_MultLoop_acc_2795_nl[18:0];
  assign nl_MultLoop_acc_1247_nl = conv_s2u_19_21(MultLoop_acc_2795_nl) + conv_s2u_20_21({(data_rsci_idat[575:558])
      , 2'b00});
  assign MultLoop_acc_1247_nl = nl_MultLoop_acc_1247_nl[20:0];
  assign nl_MultLoop_acc_2797_nl = ({(data_rsci_idat[485:468]) , 3'b001}) + conv_s2s_19_21({MultLoop_MultLoop_conc_724_18_6
      , (~ (data_rsci_idat[473:468]))});
  assign MultLoop_acc_2797_nl = nl_MultLoop_acc_2797_nl[20:0];
  assign nl_MultLoop_acc_4291_nl = conv_s2u_15_18(readslicef_21_15_6((MultLoop_acc_2797_nl)))
      + (~ (data_rsci_idat[485:468]));
  assign MultLoop_acc_4291_nl = nl_MultLoop_acc_4291_nl[17:0];
  assign nl_MultLoop_acc_2799_nl = ({(~ (data_rsci_idat[449:432])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_4692);
  assign MultLoop_acc_2799_nl = nl_MultLoop_acc_2799_nl[21:0];
  assign nl_MultLoop_acc_501_nl = conv_s2s_22_24(MultLoop_acc_2799_nl) + ({(data_rsci_idat[449:432])
      , 6'b010000});
  assign MultLoop_acc_501_nl = nl_MultLoop_acc_501_nl[23:0];
  assign nl_MultLoop_acc_2801_nl = (~ (data_rsci_idat[413:396])) + conv_s2s_17_18({MultLoop_acc_4032_cse_1
      , (data_rsci_idat[400:398])});
  assign MultLoop_acc_2801_nl = nl_MultLoop_acc_2801_nl[17:0];
  assign nl_MultLoop_acc_1246_nl = conv_s2u_18_22(MultLoop_acc_2801_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[413:396])) , 3'b001});
  assign MultLoop_acc_1246_nl = nl_MultLoop_acc_1246_nl[21:0];
  assign nl_MultLoop_acc_2884_itm_1  = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1247_nl)))
      + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4291_nl))) + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_501_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1246_nl)));
  assign nl_MultLoop_acc_497_nl = conv_s2u_12_18(data_rsci_idat[377:366]) - (data_rsci_idat[377:360]);
  assign MultLoop_acc_497_nl = nl_MultLoop_acc_497_nl[17:0];
  assign nl_MultLoop_acc_4631_nl = conv_s2u_14_19(MultLoop_acc_2802_itm_19_4[15:2])
      + conv_s2u_18_19(data_rsci_idat[251:234]);
  assign MultLoop_acc_4631_nl = nl_MultLoop_acc_4631_nl[18:0];
  assign nl_MultLoop_acc_2805_nl = ({(data_rsci_idat[179:162]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[179:162])) , 2'b01}) + conv_s2s_19_22({MultLoop_MultLoop_conc_850_18_6
      , (~ (data_rsci_idat[167:162]))});
  assign MultLoop_acc_2805_nl = nl_MultLoop_acc_2805_nl[21:0];
  assign nl_MultLoop_acc_4294_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2805_nl)))
      + (~ (data_rsci_idat[179:162]));
  assign MultLoop_acc_4294_nl = nl_MultLoop_acc_4294_nl[17:0];
  assign nl_MultLoop_acc_2806_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_13_18(data_rsci_idat[53:41]);
  assign MultLoop_acc_2806_nl = nl_MultLoop_acc_2806_nl[17:0];
  assign nl_MultLoop_acc_1240_nl = conv_s2u_18_20(MultLoop_acc_2806_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign MultLoop_acc_1240_nl = nl_MultLoop_acc_1240_nl[19:0];
  assign nl_MultLoop_acc_2883_itm_1  = conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_497_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4631_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4294_nl)))
      + conv_s2s_15_17(readslicef_20_15_5((MultLoop_acc_1240_nl)));
  assign nl_MultLoop_acc_2809_nl = (~ (data_rsci_idat[845:828])) + conv_s2s_16_18({Result_acc_216_cse_1
      , (data_rsci_idat[834:831])});
  assign MultLoop_acc_2809_nl = nl_MultLoop_acc_2809_nl[17:0];
  assign nl_MultLoop_acc_2810_nl = ({(data_rsci_idat[845:828]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2809_nl);
  assign MultLoop_acc_2810_nl = nl_MultLoop_acc_2810_nl[19:0];
  assign nl_MultLoop_acc_521_nl = conv_s2u_20_22(MultLoop_acc_2810_nl) + ({(~ (data_rsci_idat[845:828]))
      , 4'b0000});
  assign MultLoop_acc_521_nl = nl_MultLoop_acc_521_nl[21:0];
  assign nl_MultLoop_acc_2813_nl = ({(data_rsci_idat[863:846]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[863:846])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_728_18_8
      , (~ (data_rsci_idat[853:846]))});
  assign MultLoop_acc_2813_nl = nl_MultLoop_acc_2813_nl[22:0];
  assign nl_MultLoop_acc_4298_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_2813_nl)))
      + (~ (data_rsci_idat[863:846]));
  assign MultLoop_acc_4298_nl = nl_MultLoop_acc_4298_nl[17:0];
  assign nl_MultLoop_acc_4632_nl = conv_s2u_17_19(MultLoop_acc_2807_itm_18_2) + conv_s2u_18_19(data_rsci_idat[71:54]);
  assign MultLoop_acc_4632_nl = nl_MultLoop_acc_4632_nl[18:0];
  assign nl_MultLoop_acc_4633_nl = conv_s2u_19_20(MultLoop_acc_2781_cse_1[21:3])
      + ({(data_rsci_idat[395:378]) , 2'b01});
  assign MultLoop_acc_4633_nl = nl_MultLoop_acc_4633_nl[19:0];
  assign nl_MultLoop_acc_4295_nl = conv_s2s_14_15(data_rsci_idat[323:310]) + 15'b000000000000001;
  assign MultLoop_acc_4295_nl = nl_MultLoop_acc_4295_nl[14:0];
  assign nl_MultLoop_acc_2783_nl = conv_s2s_18_19(data_rsci_idat[323:306]) + conv_s2s_17_19({(MultLoop_acc_4295_nl)
      , (data_rsci_idat[309:308])});
  assign MultLoop_acc_2783_nl = nl_MultLoop_acc_2783_nl[18:0];
  assign nl_MultLoop_acc_494_nl = conv_s2u_19_20(MultLoop_acc_2783_nl) + ({(~ (data_rsci_idat[323:306]))
      , 2'b00});
  assign MultLoop_acc_494_nl = nl_MultLoop_acc_494_nl[19:0];
  assign nl_MultLoop_acc_2893_itm_1  = conv_s2s_16_18(MultLoop_acc_3930_itm_17_2)
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_521_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4298_nl)))
      + conv_s2s_15_18(readslicef_19_15_4((MultLoop_acc_4632_nl))) + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_4633_nl)))
      + conv_s2s_13_18(readslicef_20_13_7((MultLoop_acc_494_nl)));
  assign nl_MultLoop_acc_4677_nl = conv_s2u_18_19(data_rsci_idat[629:612]) + conv_s2u_17_19(MultLoop_acc_2525_cse_1[18:2]);
  assign MultLoop_acc_4677_nl = nl_MultLoop_acc_4677_nl[18:0];
  assign nl_MultLoop_acc_4304_nl = conv_s2u_15_18(readslicef_19_15_4((MultLoop_acc_4677_nl)))
      + (~ (data_rsci_idat[629:612]));
  assign MultLoop_acc_4304_nl = nl_MultLoop_acc_4304_nl[17:0];
  assign nl_MultLoop_acc_4299_nl = conv_s2s_10_11(data_rsci_idat[737:728]) + 11'b00000000001;
  assign MultLoop_acc_4299_nl = nl_MultLoop_acc_4299_nl[10:0];
  assign nl_MultLoop_acc_2816_nl = conv_s2s_20_21({(data_rsci_idat[737:720]) , 2'b00})
      + conv_s2s_18_21(data_rsci_idat[737:720]) + conv_s2s_16_21({(MultLoop_acc_4299_nl)
      , (data_rsci_idat[727:723])});
  assign MultLoop_acc_2816_nl = nl_MultLoop_acc_2816_nl[20:0];
  assign nl_MultLoop_acc_516_nl = conv_s2u_21_23(MultLoop_acc_2816_nl) + ({(~ (data_rsci_idat[737:720]))
      , 5'b00000});
  assign MultLoop_acc_516_nl = nl_MultLoop_acc_516_nl[22:0];
  assign nl_MultLoop_acc_4300_nl =  -conv_s2s_16_17(data_rsci_idat[701:686]);
  assign MultLoop_acc_4300_nl = nl_MultLoop_acc_4300_nl[16:0];
  assign nl_MultLoop_acc_514_nl = conv_s2s_19_21({(MultLoop_acc_4300_nl) , (~ (data_rsci_idat[685:684]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[701:684])) , 2'b01});
  assign MultLoop_acc_514_nl = nl_MultLoop_acc_514_nl[20:0];
  assign nl_MultLoop_acc_4301_nl =  -conv_s2s_14_15(data_rsci_idat[719:706]);
  assign MultLoop_acc_4301_nl = nl_MultLoop_acc_4301_nl[14:0];
  assign nl_MultLoop_acc_515_nl = conv_s2s_22_23({(~ (data_rsci_idat[719:702])) ,
      4'b0100}) + conv_s2s_20_23({(~ (data_rsci_idat[719:702])) , 2'b01}) + conv_s2s_19_23({(MultLoop_acc_4301_nl)
      , (~ (data_rsci_idat[705:702]))});
  assign MultLoop_acc_515_nl = nl_MultLoop_acc_515_nl[22:0];
  assign nl_MultLoop_acc_4302_nl = conv_s2s_11_12(data_rsci_idat[683:673]) + 12'b000000000001;
  assign MultLoop_acc_4302_nl = nl_MultLoop_acc_4302_nl[11:0];
  assign nl_MultLoop_acc_2821_nl = (~ (data_rsci_idat[683:666])) + conv_s2s_17_18({(MultLoop_acc_4302_nl)
      , (data_rsci_idat[672:668])});
  assign MultLoop_acc_2821_nl = nl_MultLoop_acc_2821_nl[17:0];
  assign nl_MultLoop_acc_2822_nl = conv_s2s_20_21({(~ (data_rsci_idat[683:666]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2821_nl);
  assign MultLoop_acc_2822_nl = nl_MultLoop_acc_2822_nl[20:0];
  assign nl_MultLoop_acc_1250_nl = conv_s2u_21_24(MultLoop_acc_2822_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[683:666])) , 5'b00100});
  assign MultLoop_acc_1250_nl = nl_MultLoop_acc_1250_nl[23:0];
  assign nl_MultLoop_acc_4678_nl = ({(data_rsci_idat[593:576]) , 2'b01}) + conv_s2u_19_20(MultLoop_acc_1866_itm_20_2_1);
  assign MultLoop_acc_4678_nl = nl_MultLoop_acc_4678_nl[19:0];
  assign nl_MultLoop_acc_4306_nl = conv_s2u_15_18(readslicef_20_15_5((MultLoop_acc_4678_nl)))
      + (~ (data_rsci_idat[593:576]));
  assign MultLoop_acc_4306_nl = nl_MultLoop_acc_4306_nl[17:0];
  assign nl_MultLoop_acc_1248_nl = conv_s2u_12_19(data_rsci_idat[611:600]) + conv_s2u_18_19(data_rsci_idat[611:594]);
  assign MultLoop_acc_1248_nl = nl_MultLoop_acc_1248_nl[18:0];
  assign nl_MultLoop_acc_2898_itm_1  = conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4304_nl)))
      + conv_s2s_16_18(MultLoop_acc_3532_itm_20_5_1) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_516_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_514_nl))) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_515_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1250_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4306_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_1248_nl)));
  assign nl_MultLoop_acc_4310_nl = conv_s2u_13_19(MultLoop_acc_2836_itm_19_6[13:1])
      + conv_s2u_18_19(data_rsci_idat[287:270]);
  assign MultLoop_acc_4310_nl = nl_MultLoop_acc_4310_nl[18:0];
  assign nl_MultLoop_acc_489_nl = conv_s2s_24_25({(~ (data_rsci_idat[233:216])) ,
      6'b010000}) + conv_s2s_22_25({(~ (data_rsci_idat[233:216])) , 4'b0001}) + conv_s2s_19_25({MultLoop_MultLoop_conc_702_18_6
      , (~ (data_rsci_idat[221:216]))});
  assign MultLoop_acc_489_nl = nl_MultLoop_acc_489_nl[24:0];
  assign nl_MultLoop_acc_2831_nl = (~ (data_rsci_idat[557:540])) + conv_s2s_17_18({MultLoop_acc_4146_cse_1
      , (data_rsci_idat[547:542])});
  assign MultLoop_acc_2831_nl = nl_MultLoop_acc_2831_nl[17:0];
  assign nl_MultLoop_acc_2832_nl = ({(data_rsci_idat[557:540]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2831_nl);
  assign MultLoop_acc_2832_nl = nl_MultLoop_acc_2832_nl[19:0];
  assign nl_MultLoop_acc_2833_nl = conv_s2s_22_23({(data_rsci_idat[557:540]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2832_nl);
  assign MultLoop_acc_2833_nl = nl_MultLoop_acc_2833_nl[22:0];
  assign nl_MultLoop_acc_4308_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2833_nl)))
      + (~ (data_rsci_idat[557:540]));
  assign MultLoop_acc_4308_nl = nl_MultLoop_acc_4308_nl[17:0];
  assign nl_MultLoop_acc_4309_nl =  -conv_s2s_14_15(data_rsci_idat[467:454]);
  assign MultLoop_acc_4309_nl = nl_MultLoop_acc_4309_nl[14:0];
  assign nl_MultLoop_acc_502_nl = conv_s2s_19_23({(MultLoop_acc_4309_nl) , (~ (data_rsci_idat[453:450]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[467:450])) , 4'b0001});
  assign MultLoop_acc_502_nl = nl_MultLoop_acc_502_nl[22:0];
  assign nl_MultLoop_acc_2835_nl = conv_s2s_18_19(data_rsci_idat[305:288]) + conv_s2s_16_19(data_rsci_idat[305:290]);
  assign MultLoop_acc_2835_nl = nl_MultLoop_acc_2835_nl[18:0];
  assign nl_MultLoop_acc_1244_nl = conv_s2u_19_21(MultLoop_acc_2835_nl) + conv_s2u_20_21({(data_rsci_idat[305:288])
      , 2'b00});
  assign MultLoop_acc_1244_nl = nl_MultLoop_acc_1244_nl[20:0];
  assign nl_MultLoop_acc_491_nl = conv_s2u_11_18(data_rsci_idat[269:259]) - (data_rsci_idat[269:252]);
  assign MultLoop_acc_491_nl = nl_MultLoop_acc_491_nl[17:0];
  assign nl_MultLoop_acc_2841_nl = ({(~ (data_rsci_idat[161:144])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[161:144])
      + conv_s2s_17_20({MultLoop_acc_4162_cse_1 , (data_rsci_idat[150:146])});
  assign MultLoop_acc_2841_nl = nl_MultLoop_acc_2841_nl[19:0];
  assign nl_MultLoop_acc_1242_nl = conv_s2u_20_24(MultLoop_acc_2841_nl) + conv_s2u_23_24({(~
      (data_rsci_idat[161:144])) , 5'b00100});
  assign MultLoop_acc_1242_nl = nl_MultLoop_acc_1242_nl[23:0];
  assign nl_MultLoop_acc_2897_itm_1  = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4310_nl)))
      + conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_489_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4308_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_502_nl))) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1244_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_491_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1242_nl)))
      + conv_s2s_16_18(MultLoop_acc_149_itm_23_8);
  assign nl_MultLoop_acc_1287_nl = conv_s2u_18_24(MultLoop_acc_2604_cse_1) + conv_s2u_23_24({(~
      (data_rsci_idat[845:828])) , 5'b00001});
  assign MultLoop_acc_1287_nl = nl_MultLoop_acc_1287_nl[23:0];
  assign nl_MultLoop_acc_2602_nl = ({(data_rsci_idat[89:72]) , 5'b01000}) + conv_s2s_21_23({(~
      (data_rsci_idat[89:72])) , 3'b001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_804_18_7
      , (~ (data_rsci_idat[78:72]))});
  assign MultLoop_acc_2602_nl = nl_MultLoop_acc_2602_nl[22:0];
  assign nl_MultLoop_acc_4222_nl = conv_s2u_16_18(readslicef_23_16_7((MultLoop_acc_2602_nl)))
      + (~ (data_rsci_idat[89:72]));
  assign MultLoop_acc_4222_nl = nl_MultLoop_acc_4222_nl[17:0];
  assign nl_MultLoop_acc_1268_nl = (MultLoop_acc_570_itm_21_6[15:2]) + 14'b00000000011111;
  assign MultLoop_acc_1268_nl = nl_MultLoop_acc_1268_nl[13:0];
  assign nl_MultLoop_acc_2594_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_15_18(data_rsci_idat[143:129]);
  assign MultLoop_acc_2594_nl = nl_MultLoop_acc_2594_nl[17:0];
  assign nl_MultLoop_acc_2595_nl = ({(data_rsci_idat[143:126]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2594_nl);
  assign MultLoop_acc_2595_nl = nl_MultLoop_acc_2595_nl[19:0];
  assign nl_MultLoop_acc_1271_nl = conv_s2u_20_23(MultLoop_acc_2595_nl) + conv_s2u_22_23({(data_rsci_idat[143:126])
      , 4'b0000});
  assign MultLoop_acc_1271_nl = nl_MultLoop_acc_1271_nl[22:0];
  assign nl_MultLoop_acc_2596_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_14_18(data_rsci_idat[161:148]);
  assign MultLoop_acc_2596_nl = nl_MultLoop_acc_2596_nl[17:0];
  assign nl_MultLoop_acc_1272_nl = conv_s2u_18_21(MultLoop_acc_2596_nl) + ({(data_rsci_idat[161:144])
      , 3'b001});
  assign MultLoop_acc_1272_nl = nl_MultLoop_acc_1272_nl[20:0];
  assign nl_MultLoop_acc_2598_nl = (~ (data_rsci_idat[107:90])) + conv_s2s_16_18({MultLoop_MultLoop_conc_694_15_3
      , (data_rsci_idat[95:93])});
  assign MultLoop_acc_2598_nl = nl_MultLoop_acc_2598_nl[17:0];
  assign nl_MultLoop_acc_1270_nl = conv_s2u_18_22(MultLoop_acc_2598_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[107:90])) , 3'b001});
  assign MultLoop_acc_1270_nl = nl_MultLoop_acc_1270_nl[21:0];
  assign nl_MultLoop_acc_575_nl = conv_s2s_19_26({MultLoop_MultLoop_conc_832_18_7
      , (~ (data_rsci_idat[114:108]))}) + conv_s2s_25_26({(~ (data_rsci_idat[125:108]))
      , 7'b0000001});
  assign MultLoop_acc_575_nl = nl_MultLoop_acc_575_nl[25:0];
  assign nl_MultLoop_acc_2658_itm_1  = conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_1287_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4222_nl))) + conv_s2s_16_18({(MultLoop_acc_1268_nl)
      , (MultLoop_acc_570_itm_21_6[1:0])}) + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1271_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_1272_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1270_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_575_nl)));
  assign nl_MultLoop_acc_608_nl = conv_s2s_25_26({(~ (data_rsci_idat[737:720])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[737:720])) , 5'b00001}) +
      conv_s2s_19_26({MultLoop_MultLoop_conc_856_18_7 , (~ (data_rsci_idat[726:720]))});
  assign MultLoop_acc_608_nl = nl_MultLoop_acc_608_nl[25:0];
  assign nl_MultLoop_acc_2608_nl = (~ (data_rsci_idat[629:612])) + conv_s2s_15_18({MultLoop_acc_4084_cse_1
      , (data_rsci_idat[619:616])});
  assign MultLoop_acc_2608_nl = nl_MultLoop_acc_2608_nl[17:0];
  assign nl_MultLoop_acc_2609_nl = conv_s2s_20_21({(~ (data_rsci_idat[629:612]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2608_nl);
  assign MultLoop_acc_2609_nl = nl_MultLoop_acc_2609_nl[20:0];
  assign nl_MultLoop_acc_1281_nl = conv_s2u_21_23(MultLoop_acc_2609_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[629:612])) , 4'b0100});
  assign MultLoop_acc_1281_nl = nl_MultLoop_acc_1281_nl[22:0];
  assign nl_MultLoop_acc_2610_nl = ({(data_rsci_idat[467:450]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[467:450]));
  assign MultLoop_acc_2610_nl = nl_MultLoop_acc_2610_nl[19:0];
  assign nl_MultLoop_acc_4226_nl = conv_s2u_13_19(readslicef_20_13_7((MultLoop_acc_2610_nl)))
      + conv_s2u_18_19(data_rsci_idat[467:450]);
  assign MultLoop_acc_4226_nl = nl_MultLoop_acc_4226_nl[18:0];
  assign nl_MultLoop_acc_2657_itm_1  = conv_s2s_17_18(MultLoop_acc_1227_itm_21_5)
      + conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_608_nl))) + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1281_nl)))
      + conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4226_nl)));
  assign nl_MultLoop_acc_4227_nl =  -conv_s2s_11_12(data_rsci_idat[449:439]);
  assign MultLoop_acc_4227_nl = nl_MultLoop_acc_4227_nl[11:0];
  assign nl_MultLoop_acc_593_nl = conv_s2s_25_26({(~ (data_rsci_idat[449:432])) ,
      7'b0100000}) + conv_s2s_23_26({(~ (data_rsci_idat[449:432])) , 5'b00001}) +
      conv_s2s_19_26({(MultLoop_acc_4227_nl) , (~ (data_rsci_idat[438:432]))});
  assign MultLoop_acc_593_nl = nl_MultLoop_acc_593_nl[25:0];
  assign nl_MultLoop_acc_2614_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_17_18({MultLoop_MultLoop_conc_790_16_4
      , (data_rsci_idat[383:380])});
  assign MultLoop_acc_2614_nl = nl_MultLoop_acc_2614_nl[17:0];
  assign nl_MultLoop_acc_1278_nl = conv_s2u_18_23(MultLoop_acc_2614_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[395:378])) , 4'b0001});
  assign MultLoop_acc_1278_nl = nl_MultLoop_acc_1278_nl[22:0];
  assign nl_MultLoop_acc_2616_nl = (~ (data_rsci_idat[377:360])) + conv_s2s_14_18({MultLoop_acc_4229_cse_1
      , (data_rsci_idat[367:365])});
  assign MultLoop_acc_2616_nl = nl_MultLoop_acc_2616_nl[17:0];
  assign nl_MultLoop_acc_1277_nl = conv_s2u_18_22(MultLoop_acc_2616_nl) + conv_s2u_21_22({(~
      (data_rsci_idat[377:360])) , 3'b001});
  assign MultLoop_acc_1277_nl = nl_MultLoop_acc_1277_nl[21:0];
  assign nl_MultLoop_acc_2619_nl = ({(~ (data_rsci_idat[71:54])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[71:54])
      + conv_s2s_16_20({MultLoop_acc_3955_cse_1 , (data_rsci_idat[60:57])});
  assign MultLoop_acc_2619_nl = nl_MultLoop_acc_2619_nl[19:0];
  assign nl_MultLoop_acc_1269_nl = conv_s2u_20_23(MultLoop_acc_2619_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[71:54])) , 4'b0100});
  assign MultLoop_acc_1269_nl = nl_MultLoop_acc_1269_nl[22:0];
  assign nl_MultLoop_acc_2656_itm_1  = conv_s2s_17_18(readslicef_26_17_9((MultLoop_acc_593_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1278_nl))) + conv_s2s_17_18(readslicef_22_17_5((MultLoop_acc_1277_nl)))
      + conv_s2s_17_18(readslicef_23_17_6((MultLoop_acc_1269_nl)));
  assign nl_MultLoop_acc_2559_nl = (~ (data_rsci_idat[827:810])) + conv_s2s_14_18(data_rsci_idat[827:814]);
  assign MultLoop_acc_2559_nl = nl_MultLoop_acc_2559_nl[17:0];
  assign nl_MultLoop_acc_1286_nl = conv_s2u_18_20(MultLoop_acc_2559_nl) + ({(data_rsci_idat[827:810])
      , 2'b01});
  assign MultLoop_acc_1286_nl = nl_MultLoop_acc_1286_nl[19:0];
  assign nl_MultLoop_acc_2561_nl = conv_s2s_18_19(data_rsci_idat[539:522]) + conv_s2s_15_19({MultLoop_MultLoop_conc_732_14_2
      , (data_rsci_idat[527:526])});
  assign MultLoop_acc_2561_nl = nl_MultLoop_acc_2561_nl[18:0];
  assign nl_MultLoop_acc_598_nl = conv_s2u_19_20(MultLoop_acc_2561_nl) + ({(~ (data_rsci_idat[539:522]))
      , 2'b00});
  assign MultLoop_acc_598_nl = nl_MultLoop_acc_598_nl[19:0];
  assign nl_MultLoop_acc_571_nl = conv_s2u_12_18(data_rsci_idat[53:42]) - (data_rsci_idat[53:36]);
  assign MultLoop_acc_571_nl = nl_MultLoop_acc_571_nl[17:0];
  assign nl_MultLoop_acc_2631_itm_1  = conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_1286_nl)))
      + conv_s2s_14_16(data_rsci_idat[701:688]) + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_598_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_571_nl)));
  assign nl_MultLoop_acc_4232_nl =  -conv_s2s_14_15(data_rsci_idat[863:850]);
  assign MultLoop_acc_4232_nl = nl_MultLoop_acc_4232_nl[14:0];
  assign nl_MultLoop_acc_615_nl = conv_s2s_19_23({(MultLoop_acc_4232_nl) , (~ (data_rsci_idat[849:846]))})
      + conv_s2s_22_23({(~ (data_rsci_idat[863:846])) , 4'b0001});
  assign MultLoop_acc_615_nl = nl_MultLoop_acc_615_nl[22:0];
  assign nl_MultLoop_acc_2563_nl = (~ (data_rsci_idat[755:738])) + conv_s2s_16_18(data_rsci_idat[755:740]);
  assign MultLoop_acc_2563_nl = nl_MultLoop_acc_2563_nl[17:0];
  assign nl_MultLoop_acc_1284_nl = conv_s2u_18_23(MultLoop_acc_2563_nl) + ({(data_rsci_idat[755:738])
      , 5'b00001});
  assign MultLoop_acc_1284_nl = nl_MultLoop_acc_1284_nl[22:0];
  assign nl_MultLoop_acc_2630_itm_1  = conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_615_nl)))
      + conv_s2s_15_16(readslicef_23_15_8((MultLoop_acc_1284_nl)));
  assign nl_MultLoop_acc_2565_nl = conv_s2s_18_19(data_rsci_idat[773:756]) + conv_s2s_15_19({MultLoop_acc_4233_cse_1
      , (data_rsci_idat[762:760])});
  assign MultLoop_acc_2565_nl = nl_MultLoop_acc_2565_nl[18:0];
  assign nl_MultLoop_acc_610_nl = conv_s2u_19_21(MultLoop_acc_2565_nl) + ({(~ (data_rsci_idat[773:756]))
      , 3'b000});
  assign MultLoop_acc_610_nl = nl_MultLoop_acc_610_nl[20:0];
  assign nl_MultLoop_acc_4625_nl = conv_s2u_17_19(MultLoop_acc_2566_cse_1[18:2])
      + conv_s2u_18_19(data_rsci_idat[719:702]);
  assign MultLoop_acc_4625_nl = nl_MultLoop_acc_4625_nl[18:0];
  assign nl_MultLoop_acc_4626_nl = conv_s2u_19_23(MultLoop_acc_2385_cse_1[20:2])
      + ({(data_rsci_idat[683:666]) , 5'b00001});
  assign MultLoop_acc_4626_nl = nl_MultLoop_acc_4626_nl[22:0];
  assign nl_MultLoop_acc_2569_nl = conv_s2s_21_22({(~ (data_rsci_idat[647:630]))
      , 3'b001}) + conv_s2s_18_22(MultLoop_acc_2568_cse_1);
  assign MultLoop_acc_2569_nl = nl_MultLoop_acc_2569_nl[21:0];
  assign nl_MultLoop_acc_1282_nl = conv_s2u_22_23(MultLoop_acc_2569_nl) + ({(data_rsci_idat[647:630])
      , 5'b01000});
  assign MultLoop_acc_1282_nl = nl_MultLoop_acc_1282_nl[22:0];
  assign nl_MultLoop_acc_2643_itm_1  = conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_610_nl)))
      + conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4625_nl))) + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_4626_nl)))
      + conv_s2s_15_17(readslicef_23_15_8((MultLoop_acc_1282_nl)));
  assign nl_MultLoop_acc_4627_nl = conv_s2u_15_19(Result_acc_127_cse_1[18:4]) + conv_s2u_18_19(data_rsci_idat[575:558]);
  assign MultLoop_acc_4627_nl = nl_MultLoop_acc_4627_nl[18:0];
  assign nl_MultLoop_acc_4234_nl =  -conv_s2s_16_17(data_rsci_idat[593:578]);
  assign MultLoop_acc_4234_nl = nl_MultLoop_acc_4234_nl[16:0];
  assign nl_MultLoop_acc_601_nl = conv_s2s_19_21({(MultLoop_acc_4234_nl) , (~ (data_rsci_idat[577:576]))})
      + conv_s2s_20_21({(~ (data_rsci_idat[593:576])) , 2'b01});
  assign MultLoop_acc_601_nl = nl_MultLoop_acc_601_nl[20:0];
  assign nl_MultLoop_acc_2573_nl = ({(data_rsci_idat[485:468]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_692_18_7
      , (~ (data_rsci_idat[474:468]))});
  assign MultLoop_acc_2573_nl = nl_MultLoop_acc_2573_nl[21:0];
  assign nl_MultLoop_acc_4236_nl = conv_s2u_15_18(readslicef_22_15_7((MultLoop_acc_2573_nl)))
      + (~ (data_rsci_idat[485:468]));
  assign MultLoop_acc_4236_nl = nl_MultLoop_acc_4236_nl[17:0];
  assign nl_MultLoop_acc_2642_itm_1  = conv_s2s_15_17(readslicef_19_15_4((MultLoop_acc_4627_nl)))
      + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_601_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4236_nl)))
      + conv_s2s_15_17(MultLoop_acc_307_itm_21_7);
  assign nl_MultLoop_acc_2575_nl = conv_s2s_20_21({(~ (data_rsci_idat[341:324]))
      , 2'b01}) + conv_s2s_18_21(MultLoop_acc_2574_cse_1);
  assign MultLoop_acc_2575_nl = nl_MultLoop_acc_2575_nl[20:0];
  assign nl_MultLoop_acc_1276_nl = conv_s2u_21_22(MultLoop_acc_2575_nl) + ({(data_rsci_idat[341:324])
      , 4'b0100});
  assign MultLoop_acc_1276_nl = nl_MultLoop_acc_1276_nl[21:0];
  assign nl_MultLoop_acc_4237_nl =  -conv_s2s_13_14(data_rsci_idat[215:203]);
  assign MultLoop_acc_4237_nl = nl_MultLoop_acc_4237_nl[13:0];
  assign nl_MultLoop_acc_580_nl = conv_s2s_23_24({(~ (data_rsci_idat[215:198])) ,
      5'b00100}) + conv_s2s_20_24({(~ (data_rsci_idat[215:198])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4237_nl)
      , (~ (data_rsci_idat[202:198]))});
  assign MultLoop_acc_580_nl = nl_MultLoop_acc_580_nl[23:0];
  assign nl_MultLoop_acc_2578_nl = (~ (data_rsci_idat[179:162])) + conv_s2s_16_18(data_rsci_idat[179:164]);
  assign MultLoop_acc_2578_nl = nl_MultLoop_acc_2578_nl[17:0];
  assign nl_MultLoop_acc_1273_nl = conv_s2u_18_22(MultLoop_acc_2578_nl) + ({(data_rsci_idat[179:162])
      , 4'b0001});
  assign MultLoop_acc_1273_nl = nl_MultLoop_acc_1273_nl[21:0];
  assign nl_MultLoop_acc_591_nl = conv_s2s_18_21(~ (data_rsci_idat[413:396])) + ({(data_rsci_idat[413:396])
      , 3'b001});
  assign MultLoop_acc_591_nl = nl_MultLoop_acc_591_nl[20:0];
  assign nl_MultLoop_acc_4238_nl =  -conv_s2s_15_16(data_rsci_idat[791:777]);
  assign MultLoop_acc_4238_nl = nl_MultLoop_acc_4238_nl[15:0];
  assign nl_MultLoop_acc_611_nl = conv_s2s_19_22({(MultLoop_acc_4238_nl) , (~ (data_rsci_idat[776:774]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[791:774])) , 3'b001});
  assign MultLoop_acc_611_nl = nl_MultLoop_acc_611_nl[21:0];
  assign nl_MultLoop_acc_585_nl = conv_s2s_18_20(~ (data_rsci_idat[305:288])) + ({(data_rsci_idat[305:288])
      , 2'b01});
  assign MultLoop_acc_585_nl = nl_MultLoop_acc_585_nl[19:0];
  assign nl_MultLoop_acc_2620_nl = (readslicef_22_12_10((MultLoop_acc_611_nl))) +
      conv_s2s_10_12(readslicef_20_10_10((MultLoop_acc_585_nl)));
  assign MultLoop_acc_2620_nl = nl_MultLoop_acc_2620_nl[11:0];
  assign nl_MultLoop_acc_2641_itm_1  = conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1276_nl)))
      + conv_s2s_15_17(readslicef_24_15_9((MultLoop_acc_580_nl))) + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1273_nl)))
      + conv_s2s_13_17(readslicef_21_13_8((MultLoop_acc_591_nl))) + conv_s2s_12_17(MultLoop_acc_2620_nl);
  assign nl_MultLoop_acc_2579_nl = conv_s2s_20_21({(~ (data_rsci_idat[665:648]))
      , 2'b01}) + conv_s2s_18_21(~ (data_rsci_idat[665:648]));
  assign MultLoop_acc_2579_nl = nl_MultLoop_acc_2579_nl[20:0];
  assign nl_MultLoop_acc_605_nl = conv_s2s_21_25(MultLoop_acc_2579_nl) + ({(data_rsci_idat[665:648])
      , 7'b0000100});
  assign MultLoop_acc_605_nl = nl_MultLoop_acc_605_nl[24:0];
  assign nl_MultLoop_acc_2581_nl = ({(data_rsci_idat[611:594]) , 5'b00100}) + conv_s2s_20_23({(~
      (data_rsci_idat[611:594])) , 2'b01}) + conv_s2s_18_23(~ (data_rsci_idat[611:594]));
  assign MultLoop_acc_2581_nl = nl_MultLoop_acc_2581_nl[22:0];
  assign nl_MultLoop_acc_4239_nl = conv_s2u_16_19(readslicef_23_16_7((MultLoop_acc_2581_nl)))
      + conv_s2u_18_19(data_rsci_idat[611:594]);
  assign MultLoop_acc_4239_nl = nl_MultLoop_acc_4239_nl[18:0];
  assign nl_MultLoop_acc_596_nl = conv_s2u_12_18(data_rsci_idat[503:492]) - (data_rsci_idat[503:486]);
  assign MultLoop_acc_596_nl = nl_MultLoop_acc_596_nl[17:0];
  assign nl_MultLoop_acc_2653_itm_1  = conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_605_nl)))
      + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4239_nl))) + conv_s2s_16_18(MultLoop_acc_1152_itm_18_3)
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_596_nl)));
  assign nl_MultLoop_acc_4629_nl = conv_s2u_14_19(MultLoop_acc_2591_cse_1[18:5])
      + conv_s2u_18_19(data_rsci_idat[251:234]);
  assign MultLoop_acc_4629_nl = nl_MultLoop_acc_4629_nl[18:0];
  assign nl_MultLoop_acc_4628_nl = conv_s2u_19_21(MultLoop_acc_1603_cse_1[21:3])
      + ({(data_rsci_idat[521:504]) , 3'b001});
  assign MultLoop_acc_4628_nl = nl_MultLoop_acc_4628_nl[20:0];
  assign nl_MultLoop_acc_4675_nl = conv_s2u_14_18(MultLoop_acc_2584_cse_1[18:5])
      + (~ (data_rsci_idat[431:414]));
  assign MultLoop_acc_4675_nl = nl_MultLoop_acc_4675_nl[17:0];
  assign nl_MultLoop_acc_2586_nl = (~ (data_rsci_idat[323:306])) + conv_s2s_17_18({MultLoop_MultLoop_conc_778_16_6
      , (data_rsci_idat[313:308])});
  assign MultLoop_acc_2586_nl = nl_MultLoop_acc_2586_nl[17:0];
  assign nl_MultLoop_acc_2587_nl = ({(data_rsci_idat[323:306]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2586_nl);
  assign MultLoop_acc_2587_nl = nl_MultLoop_acc_2587_nl[19:0];
  assign nl_MultLoop_acc_4242_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_2587_nl)))
      + (~ (data_rsci_idat[323:306]));
  assign MultLoop_acc_4242_nl = nl_MultLoop_acc_4242_nl[17:0];
  assign nl_MultLoop_acc_2590_nl = ({(data_rsci_idat[287:270]) , 6'b000100}) + conv_s2s_20_24({(~
      (data_rsci_idat[287:270])) , 2'b01}) + conv_s2s_19_24({MultLoop_MultLoop_conc_814_18_8
      , (~ (data_rsci_idat[277:270]))});
  assign MultLoop_acc_2590_nl = nl_MultLoop_acc_2590_nl[23:0];
  assign nl_MultLoop_acc_4244_nl = conv_s2u_16_18(readslicef_24_16_8((MultLoop_acc_2590_nl)))
      + (~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_4244_nl = nl_MultLoop_acc_4244_nl[17:0];
  assign nl_MultLoop_acc_2593_nl = conv_s2s_24_25({(~ (data_rsci_idat[233:216]))
      , 6'b001000}) + conv_s2s_22_25(MultLoop_acc_2592_cse_1);
  assign MultLoop_acc_2593_nl = nl_MultLoop_acc_2593_nl[24:0];
  assign nl_MultLoop_acc_581_nl = conv_s2s_25_26(MultLoop_acc_2593_nl) + ({(data_rsci_idat[233:216])
      , 8'b01000000});
  assign MultLoop_acc_581_nl = nl_MultLoop_acc_581_nl[25:0];
  assign nl_MultLoop_acc_2659_itm_1  = conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4629_nl)))
      + conv_s2s_16_18(MultLoop_acc_1275_itm_20_5) + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_4628_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4675_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4242_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4244_nl))) + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_581_nl)))
      + conv_s2s_16_18(MultLoop_acc_579_itm_19_4);
  assign nl_MultLoop_acc_2723_nl = conv_s2s_18_19(data_rsci_idat[755:738]) + conv_s2s_14_19(data_rsci_idat[755:742]);
  assign MultLoop_acc_2723_nl = nl_MultLoop_acc_2723_nl[18:0];
  assign nl_MultLoop_acc_1266_nl = conv_s2u_19_21(MultLoop_acc_2723_nl) + conv_s2u_20_21({(data_rsci_idat[755:738])
      , 2'b00});
  assign MultLoop_acc_1266_nl = nl_MultLoop_acc_1266_nl[20:0];
  assign nl_MultLoop_acc_2725_nl = ({(data_rsci_idat[701:684]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_782_18_8
      , (~ (data_rsci_idat[691:684]))});
  assign MultLoop_acc_2725_nl = nl_MultLoop_acc_2725_nl[19:0];
  assign nl_MultLoop_acc_4246_nl = (~ (data_rsci_idat[701:684])) + conv_s2s_14_18(readslicef_20_14_6((MultLoop_acc_2725_nl)));
  assign MultLoop_acc_4246_nl = nl_MultLoop_acc_4246_nl[17:0];
  assign nl_MultLoop_acc_4247_nl = conv_s2u_18_21(MultLoop_acc_4246_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[701:684])) , 2'b01});
  assign MultLoop_acc_4247_nl = nl_MultLoop_acc_4247_nl[20:0];
  assign nl_MultLoop_acc_4248_nl =  -conv_s2s_10_11(data_rsci_idat[395:386]);
  assign MultLoop_acc_4248_nl = nl_MultLoop_acc_4248_nl[10:0];
  assign nl_MultLoop_acc_2729_nl = ({(data_rsci_idat[395:378]) , 4'b0100}) + conv_s2s_20_22({(~
      (data_rsci_idat[395:378])) , 2'b01}) + conv_s2s_19_22({(MultLoop_acc_4248_nl)
      , (~ (data_rsci_idat[385:378]))});
  assign MultLoop_acc_2729_nl = nl_MultLoop_acc_2729_nl[21:0];
  assign nl_MultLoop_acc_4249_nl = (~ (data_rsci_idat[395:378])) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_2729_nl)));
  assign MultLoop_acc_4249_nl = nl_MultLoop_acc_4249_nl[17:0];
  assign nl_MultLoop_acc_4250_nl = conv_s2u_18_21(MultLoop_acc_4249_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[395:378])) , 2'b01});
  assign MultLoop_acc_4250_nl = nl_MultLoop_acc_4250_nl[20:0];
  assign nl_MultLoop_acc_4251_nl =  -conv_s2s_13_14(data_rsci_idat[17:5]);
  assign MultLoop_acc_4251_nl = nl_MultLoop_acc_4251_nl[13:0];
  assign nl_MultLoop_acc_523_nl = conv_s2s_23_24({(~ (data_rsci_idat[17:0])) , 5'b00100})
      + conv_s2s_20_24({(~ (data_rsci_idat[17:0])) , 2'b01}) + conv_s2s_19_24({(MultLoop_acc_4251_nl)
      , (~ (data_rsci_idat[4:0]))});
  assign MultLoop_acc_523_nl = nl_MultLoop_acc_523_nl[23:0];
  assign nl_MultLoop_acc_2773_itm_1  = conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_1266_nl)))
      + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_4247_nl))) + conv_s2s_17_18(readslicef_21_17_4((MultLoop_acc_4250_nl)))
      + conv_s2s_17_18(readslicef_24_17_7((MultLoop_acc_523_nl)));
  assign nl_MultLoop_acc_2667_nl = (~ (data_rsci_idat[863:846])) + conv_s2s_15_18(data_rsci_idat[863:849]);
  assign MultLoop_acc_2667_nl = nl_MultLoop_acc_2667_nl[17:0];
  assign nl_MultLoop_acc_1267_nl = conv_s2u_18_21(MultLoop_acc_2667_nl) + ({(data_rsci_idat[863:846])
      , 3'b001});
  assign MultLoop_acc_1267_nl = nl_MultLoop_acc_1267_nl[20:0];
  assign nl_MultLoop_acc_567_nl = conv_s2s_18_24(~ (data_rsci_idat[827:810])) + ({(data_rsci_idat[827:810])
      , 6'b000001});
  assign MultLoop_acc_567_nl = nl_MultLoop_acc_567_nl[23:0];
  assign nl_MultLoop_acc_559_nl = conv_s2s_19_23({MultLoop_MultLoop_conc_838_18_4
      , (~ (data_rsci_idat[669:666]))}) + conv_s2s_22_23({(~ (data_rsci_idat[683:666]))
      , 4'b0001});
  assign MultLoop_acc_559_nl = nl_MultLoop_acc_559_nl[22:0];
  assign nl_MultLoop_acc_4630_nl = conv_s2u_19_20(MultLoop_acc_2669_itm_20_2_1) +
      ({(data_rsci_idat[557:540]) , 2'b01});
  assign MultLoop_acc_4630_nl = nl_MultLoop_acc_4630_nl[19:0];
  assign nl_MultLoop_acc_2750_itm_1  = conv_s2s_14_16(readslicef_21_14_7((MultLoop_acc_1267_nl)))
      + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_567_nl))) + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_559_nl)))
      + conv_s2s_14_16(readslicef_20_14_6((MultLoop_acc_4630_nl)));
  assign nl_MultLoop_acc_2671_nl = ({(data_rsci_idat[503:486]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_742_18_6
      , (~ (data_rsci_idat[491:486]))});
  assign MultLoop_acc_2671_nl = nl_MultLoop_acc_2671_nl[19:0];
  assign nl_MultLoop_acc_2672_nl = conv_s2s_22_23({(data_rsci_idat[503:486]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2671_nl);
  assign MultLoop_acc_2672_nl = nl_MultLoop_acc_2672_nl[22:0];
  assign nl_MultLoop_acc_4254_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2672_nl)))
      + (~ (data_rsci_idat[503:486]));
  assign MultLoop_acc_4254_nl = nl_MultLoop_acc_4254_nl[17:0];
  assign nl_MultLoop_acc_2673_nl = ({(data_rsci_idat[449:432]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[449:432]));
  assign MultLoop_acc_2673_nl = nl_MultLoop_acc_2673_nl[20:0];
  assign nl_MultLoop_acc_546_nl = conv_s2s_21_24(MultLoop_acc_2673_nl) + conv_s2s_23_24({(data_rsci_idat[449:432])
      , 5'b00000});
  assign MultLoop_acc_546_nl = nl_MultLoop_acc_546_nl[23:0];
  assign nl_MultLoop_acc_540_nl = conv_s2s_18_23(~ (data_rsci_idat[341:324])) + ({(data_rsci_idat[341:324])
      , 5'b00001});
  assign MultLoop_acc_540_nl = nl_MultLoop_acc_540_nl[22:0];
  assign nl_MultLoop_acc_2749_itm_1  = conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4254_nl)))
      + conv_s2s_14_16(readslicef_24_14_10((MultLoop_acc_546_nl))) + conv_s2s_14_16(readslicef_23_14_9((MultLoop_acc_540_nl)))
      + conv_s2s_14_16(MultLoop_acc_541_itm_23_8[15:2]);
  assign nl_MultLoop_acc_4255_nl =  -conv_s2s_15_16(data_rsci_idat[305:291]);
  assign MultLoop_acc_4255_nl = nl_MultLoop_acc_4255_nl[15:0];
  assign nl_MultLoop_acc_538_nl = conv_s2s_19_22({(MultLoop_acc_4255_nl) , (~ (data_rsci_idat[290:288]))})
      + conv_s2s_21_22({(~ (data_rsci_idat[305:288])) , 3'b001});
  assign MultLoop_acc_538_nl = nl_MultLoop_acc_538_nl[21:0];
  assign nl_MultLoop_acc_2676_nl = ({(data_rsci_idat[287:270]) , 4'b0001}) + conv_s2s_19_22({MultLoop_MultLoop_conc_752_18_6
      , (~ (data_rsci_idat[275:270]))});
  assign MultLoop_acc_2676_nl = nl_MultLoop_acc_2676_nl[21:0];
  assign nl_MultLoop_acc_4257_nl = conv_s2u_16_18(readslicef_22_16_6((MultLoop_acc_2676_nl)))
      + (~ (data_rsci_idat[287:270]));
  assign MultLoop_acc_4257_nl = nl_MultLoop_acc_4257_nl[17:0];
  assign nl_MultLoop_acc_1255_nl = conv_s2u_13_19(data_rsci_idat[233:221]) + conv_s2u_18_19(data_rsci_idat[233:216]);
  assign MultLoop_acc_1255_nl = nl_MultLoop_acc_1255_nl[18:0];
  assign nl_MultLoop_acc_535_nl = conv_s2u_13_18(data_rsci_idat[251:239]) - (data_rsci_idat[251:234]);
  assign MultLoop_acc_535_nl = nl_MultLoop_acc_535_nl[17:0];
  assign nl_MultLoop_acc_2748_itm_1  = conv_s2s_14_16(readslicef_22_14_8((MultLoop_acc_538_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_4257_nl))) + conv_s2s_14_16(readslicef_19_14_5((MultLoop_acc_1255_nl)))
      + conv_s2s_14_16(readslicef_18_14_4((MultLoop_acc_535_nl)));
  assign nl_MultLoop_acc_2678_nl = ({(data_rsci_idat[791:774]) , 2'b01}) + conv_s2s_19_20({MultLoop_MultLoop_conc_676_18_6
      , (~ (data_rsci_idat[779:774]))});
  assign MultLoop_acc_2678_nl = nl_MultLoop_acc_2678_nl[19:0];
  assign nl_MultLoop_acc_2679_nl = conv_s2s_22_23({(data_rsci_idat[791:774]) , 4'b0000})
      + conv_s2s_20_23(MultLoop_acc_2678_nl);
  assign MultLoop_acc_2679_nl = nl_MultLoop_acc_2679_nl[22:0];
  assign nl_MultLoop_acc_4259_nl = conv_s2u_17_18(readslicef_23_17_6((MultLoop_acc_2679_nl)))
      + (~ (data_rsci_idat[791:774]));
  assign MultLoop_acc_4259_nl = nl_MultLoop_acc_4259_nl[17:0];
  assign nl_MultLoop_acc_1261_nl = conv_s2u_14_19(data_rsci_idat[539:526]) + conv_s2u_18_19(data_rsci_idat[539:522]);
  assign MultLoop_acc_1261_nl = nl_MultLoop_acc_1261_nl[18:0];
  assign nl_MultLoop_acc_2747_itm_1  = conv_s2s_15_16(readslicef_18_15_3((MultLoop_acc_4259_nl)))
      + conv_s2s_15_16(readslicef_19_15_4((MultLoop_acc_1261_nl)));
  assign nl_MultLoop_acc_544_nl = conv_s2u_13_18(data_rsci_idat[413:401]) - (data_rsci_idat[413:396]);
  assign MultLoop_acc_544_nl = nl_MultLoop_acc_544_nl[17:0];
  assign nl_MultLoop_acc_2681_nl = ({(~ (data_rsci_idat[377:360])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2500_cse_1);
  assign MultLoop_acc_2681_nl = nl_MultLoop_acc_2681_nl[19:0];
  assign nl_MultLoop_acc_1257_nl = conv_s2u_20_22(MultLoop_acc_2681_nl) + ({(data_rsci_idat[377:360])
      , 4'b0100});
  assign MultLoop_acc_1257_nl = nl_MultLoop_acc_1257_nl[21:0];
  assign nl_MultLoop_acc_4260_nl =  -conv_s2s_11_12(data_rsci_idat[269:259]);
  assign MultLoop_acc_4260_nl = nl_MultLoop_acc_4260_nl[11:0];
  assign nl_MultLoop_acc_2683_nl = ({(data_rsci_idat[269:252]) , 3'b001}) + conv_s2s_19_21({(MultLoop_acc_4260_nl)
      , (~ (data_rsci_idat[258:252]))});
  assign MultLoop_acc_2683_nl = nl_MultLoop_acc_2683_nl[20:0];
  assign nl_MultLoop_acc_4261_nl = conv_s2u_14_18(readslicef_21_14_7((MultLoop_acc_2683_nl)))
      + (~ (data_rsci_idat[269:252]));
  assign MultLoop_acc_4261_nl = nl_MultLoop_acc_4261_nl[17:0];
  assign nl_MultLoop_acc_2684_nl = conv_s2s_18_19(data_rsci_idat[215:198]) + conv_s2s_16_19(data_rsci_idat[215:200]);
  assign MultLoop_acc_2684_nl = nl_MultLoop_acc_2684_nl[18:0];
  assign nl_MultLoop_acc_1254_nl = conv_s2u_19_22(MultLoop_acc_2684_nl) + conv_s2u_21_22({(data_rsci_idat[215:198])
      , 3'b000});
  assign MultLoop_acc_1254_nl = nl_MultLoop_acc_1254_nl[21:0];
  assign nl_MultLoop_acc_2761_itm_1  = conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_544_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1257_nl))) + conv_s2s_15_17(readslicef_18_15_3((MultLoop_acc_4261_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_1254_nl)));
  assign nl_MultLoop_acc_4263_nl = conv_s2s_14_15(data_rsci_idat[467:454]) + 15'b000000000000001;
  assign MultLoop_acc_4263_nl = nl_MultLoop_acc_4263_nl[14:0];
  assign nl_MultLoop_acc_2666_nl = (~ (data_rsci_idat[467:450])) + conv_s2s_17_18({(MultLoop_acc_4263_nl)
      , (data_rsci_idat[453:452])});
  assign MultLoop_acc_2666_nl = nl_MultLoop_acc_2666_nl[17:0];
  assign nl_MultLoop_acc_1259_nl = conv_s2u_18_21(MultLoop_acc_2666_nl) + conv_s2u_20_21({(~
      (data_rsci_idat[467:450])) , 2'b01});
  assign MultLoop_acc_1259_nl = nl_MultLoop_acc_1259_nl[20:0];
  assign nl_MultLoop_acc_2733_nl = conv_s2s_9_10(data_rsci_idat[179:171]) + 10'b0001101001;
  assign MultLoop_acc_2733_nl = nl_MultLoop_acc_2733_nl[9:0];
  assign nl_MultLoop_acc_2743_nl = MultLoop_acc_528_itm_24_10 + conv_s2s_13_15(readslicef_21_13_8((MultLoop_acc_1259_nl)))
      + conv_s2s_12_15(MultLoop_acc_1476_itm_18_2[16:5]) + conv_s2s_11_15(MultLoop_acc_340_itm_17_3[14:4])
      + conv_s2s_10_15(MultLoop_acc_2733_nl);
  assign MultLoop_acc_2743_nl = nl_MultLoop_acc_2743_nl[14:0];
  assign nl_MultLoop_acc_1253_nl = conv_s2u_18_21(MultLoop_acc_2685_cse_1) + ({(data_rsci_idat[125:108])
      , 3'b001});
  assign MultLoop_acc_1253_nl = nl_MultLoop_acc_1253_nl[20:0];
  assign nl_MultLoop_acc_2687_nl = (~ (data_rsci_idat[143:126])) + conv_s2s_17_18({MultLoop_acc_4021_cse_1
      , (data_rsci_idat[131:128])});
  assign MultLoop_acc_2687_nl = nl_MultLoop_acc_2687_nl[17:0];
  assign nl_MultLoop_acc_2688_nl = ({(data_rsci_idat[143:126]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2687_nl);
  assign MultLoop_acc_2688_nl = nl_MultLoop_acc_2688_nl[19:0];
  assign nl_MultLoop_acc_530_nl = conv_s2u_20_22(MultLoop_acc_2688_nl) + ({(~ (data_rsci_idat[143:126]))
      , 4'b0000});
  assign MultLoop_acc_530_nl = nl_MultLoop_acc_530_nl[21:0];
  assign nl_MultLoop_acc_2760_itm_1  = conv_s2s_15_17(MultLoop_acc_2743_nl) + conv_s2s_15_17(readslicef_21_15_6((MultLoop_acc_1253_nl)))
      + conv_s2s_15_17(readslicef_22_15_7((MultLoop_acc_530_nl)));
  assign nl_MultLoop_acc_2689_nl = ({(data_rsci_idat[845:828]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[845:828]));
  assign MultLoop_acc_2689_nl = nl_MultLoop_acc_2689_nl[19:0];
  assign nl_MultLoop_acc_568_nl = conv_s2s_20_25(MultLoop_acc_2689_nl) + conv_s2s_24_25({(data_rsci_idat[845:828])
      , 6'b000000});
  assign MultLoop_acc_568_nl = nl_MultLoop_acc_568_nl[24:0];
  assign nl_MultLoop_acc_4264_nl = conv_s2s_10_11(data_rsci_idat[773:764]) + 11'b00000000001;
  assign MultLoop_acc_4264_nl = nl_MultLoop_acc_4264_nl[10:0];
  assign nl_MultLoop_acc_2691_nl = conv_s2s_18_19(data_rsci_idat[773:756]) + conv_s2s_14_19({(MultLoop_acc_4264_nl)
      , (data_rsci_idat[763:761])});
  assign MultLoop_acc_2691_nl = nl_MultLoop_acc_2691_nl[18:0];
  assign nl_MultLoop_acc_564_nl = conv_s2u_19_21(MultLoop_acc_2691_nl) + ({(~ (data_rsci_idat[773:756]))
      , 3'b000});
  assign MultLoop_acc_564_nl = nl_MultLoop_acc_564_nl[20:0];
  assign nl_MultLoop_acc_2692_nl = ({(data_rsci_idat[737:720]) , 3'b001}) + conv_s2s_18_21(~
      (data_rsci_idat[737:720]));
  assign MultLoop_acc_2692_nl = nl_MultLoop_acc_2692_nl[20:0];
  assign nl_MultLoop_acc_562_nl = conv_s2s_21_24(MultLoop_acc_2692_nl) + conv_s2s_23_24({(data_rsci_idat[737:720])
      , 5'b00000});
  assign MultLoop_acc_562_nl = nl_MultLoop_acc_562_nl[23:0];
  assign nl_MultLoop_acc_2694_nl = ({(~ (data_rsci_idat[719:702])) , 2'b00}) + conv_s2s_19_20(MultLoop_acc_2566_cse_1);
  assign MultLoop_acc_2694_nl = nl_MultLoop_acc_2694_nl[19:0];
  assign nl_MultLoop_acc_1265_nl = conv_s2u_20_24(MultLoop_acc_2694_nl) + ({(data_rsci_idat[719:702])
      , 6'b000100});
  assign MultLoop_acc_1265_nl = nl_MultLoop_acc_1265_nl[23:0];
  assign nl_MultLoop_acc_2770_itm_1  = conv_s2s_16_18(readslicef_25_16_9((MultLoop_acc_568_nl)))
      + conv_s2s_16_18(readslicef_21_16_5((MultLoop_acc_564_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_562_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1265_nl)));
  assign nl_MultLoop_acc_2703_nl = (~ (data_rsci_idat[611:594])) + conv_s2s_17_18({MultLoop_MultLoop_conc_774_16_4
      , (data_rsci_idat[599:596])});
  assign MultLoop_acc_2703_nl = nl_MultLoop_acc_2703_nl[17:0];
  assign nl_MultLoop_acc_1262_nl = conv_s2u_18_23(MultLoop_acc_2703_nl) + conv_s2u_22_23({(~
      (data_rsci_idat[611:594])) , 4'b0001});
  assign MultLoop_acc_1262_nl = nl_MultLoop_acc_1262_nl[22:0];
  assign nl_MultLoop_acc_2704_nl = ({(data_rsci_idat[575:558]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[575:558]));
  assign MultLoop_acc_2704_nl = nl_MultLoop_acc_2704_nl[19:0];
  assign nl_MultLoop_acc_2705_nl = ({(~ (data_rsci_idat[575:558])) , 4'b0000}) +
      conv_s2s_20_22(MultLoop_acc_2704_nl);
  assign MultLoop_acc_2705_nl = nl_MultLoop_acc_2705_nl[21:0];
  assign nl_MultLoop_acc_553_nl = conv_s2s_22_26(MultLoop_acc_2705_nl) + ({(data_rsci_idat[575:558])
      , 8'b00010000});
  assign MultLoop_acc_553_nl = nl_MultLoop_acc_553_nl[25:0];
  assign nl_MultLoop_acc_2696_nl = ({(~ (data_rsci_idat[665:648])) , 4'b0000}) +
      conv_s2s_19_22(MultLoop_acc_2073_cse_1);
  assign MultLoop_acc_2696_nl = nl_MultLoop_acc_2696_nl[21:0];
  assign nl_MultLoop_acc_1264_nl = conv_s2u_22_24(MultLoop_acc_2696_nl) + ({(data_rsci_idat[665:648])
      , 6'b010000});
  assign MultLoop_acc_1264_nl = nl_MultLoop_acc_1264_nl[23:0];
  assign nl_MultLoop_acc_2697_nl = (~ (data_rsci_idat[629:612])) + conv_s2s_14_18(data_rsci_idat[629:616]);
  assign MultLoop_acc_2697_nl = nl_MultLoop_acc_2697_nl[17:0];
  assign nl_MultLoop_acc_1263_nl = conv_s2u_18_22(MultLoop_acc_2697_nl) + ({(data_rsci_idat[629:612])
      , 4'b0001});
  assign MultLoop_acc_1263_nl = nl_MultLoop_acc_1263_nl[21:0];
  assign nl_MultLoop_acc_2698_nl = ({(data_rsci_idat[647:630]) , 4'b0001}) + conv_s2s_18_22(~
      (data_rsci_idat[647:630]));
  assign MultLoop_acc_2698_nl = nl_MultLoop_acc_2698_nl[21:0];
  assign nl_MultLoop_acc_4265_nl = conv_s2u_15_19(readslicef_22_15_7((MultLoop_acc_2698_nl)))
      + conv_s2u_18_19(data_rsci_idat[647:630]);
  assign MultLoop_acc_4265_nl = nl_MultLoop_acc_4265_nl[18:0];
  assign nl_MultLoop_acc_4266_nl = conv_s2s_10_11(data_rsci_idat[593:584]) + 11'b00000000001;
  assign MultLoop_acc_4266_nl = nl_MultLoop_acc_4266_nl[10:0];
  assign nl_MultLoop_acc_2700_nl = (~ (data_rsci_idat[593:576])) + conv_s2s_16_18({(MultLoop_acc_4266_nl)
      , (data_rsci_idat[583:579])});
  assign MultLoop_acc_2700_nl = nl_MultLoop_acc_2700_nl[17:0];
  assign nl_MultLoop_acc_2701_nl = ({(data_rsci_idat[593:576]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2700_nl);
  assign MultLoop_acc_2701_nl = nl_MultLoop_acc_2701_nl[19:0];
  assign nl_MultLoop_acc_554_nl = conv_s2u_20_23(MultLoop_acc_2701_nl) + ({(~ (data_rsci_idat[593:576]))
      , 5'b00000});
  assign MultLoop_acc_554_nl = nl_MultLoop_acc_554_nl[22:0];
  assign nl_MultLoop_acc_2707_nl = ({(~ (data_rsci_idat[521:504])) , 2'b00}) + conv_s2s_18_20(data_rsci_idat[521:504])
      + conv_s2s_14_20(data_rsci_idat[521:508]);
  assign MultLoop_acc_2707_nl = nl_MultLoop_acc_2707_nl[19:0];
  assign nl_MultLoop_acc_1260_nl = conv_s2u_20_22(MultLoop_acc_2707_nl) + ({(data_rsci_idat[521:504])
      , 4'b0100});
  assign MultLoop_acc_1260_nl = nl_MultLoop_acc_1260_nl[21:0];
  assign nl_MultLoop_acc_2709_nl = ({(data_rsci_idat[485:468]) , 5'b00001}) + conv_s2s_19_23({MultLoop_MultLoop_conc_796_18_8
      , (~ (data_rsci_idat[475:468]))});
  assign MultLoop_acc_2709_nl = nl_MultLoop_acc_2709_nl[22:0];
  assign nl_MultLoop_acc_4269_nl = conv_s2u_15_18(readslicef_23_15_8((MultLoop_acc_2709_nl)))
      + (~ (data_rsci_idat[485:468]));
  assign MultLoop_acc_4269_nl = nl_MultLoop_acc_4269_nl[17:0];
  assign nl_MultLoop_acc_2775_itm_1  = conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_1262_nl)))
      + conv_s2s_16_18(readslicef_26_16_10((MultLoop_acc_553_nl))) + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1264_nl)))
      + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1263_nl))) + conv_s2s_16_18(readslicef_19_16_3((MultLoop_acc_4265_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_554_nl))) + conv_s2s_16_18(readslicef_22_16_6((MultLoop_acc_1260_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4269_nl)));
  assign nl_MultLoop_acc_2722_nl = ({(data_rsci_idat[809:792]) , 2'b01}) + conv_s2s_18_20(~
      (data_rsci_idat[809:792]));
  assign MultLoop_acc_2722_nl = nl_MultLoop_acc_2722_nl[19:0];
  assign nl_MultLoop_acc_4275_nl = conv_s2u_12_19(readslicef_20_12_8((MultLoop_acc_2722_nl)))
      + conv_s2u_18_19(data_rsci_idat[809:792]);
  assign MultLoop_acc_4275_nl = nl_MultLoop_acc_4275_nl[18:0];
  assign nl_MultLoop_acc_526_nl = conv_s2u_12_18(data_rsci_idat[71:60]) - (data_rsci_idat[71:54]);
  assign MultLoop_acc_526_nl = nl_MultLoop_acc_526_nl[17:0];
  assign nl_MultLoop_acc_4676_nl = conv_s2u_18_19(data_rsci_idat[35:18]) + conv_s2u_16_19(MultLoop_acc_2340_itm_19_4);
  assign MultLoop_acc_4676_nl = nl_MultLoop_acc_4676_nl[18:0];
  assign nl_MultLoop_acc_4274_nl = conv_s2u_15_18(readslicef_19_15_4((MultLoop_acc_4676_nl)))
      + (~ (data_rsci_idat[35:18]));
  assign MultLoop_acc_4274_nl = nl_MultLoop_acc_4274_nl[17:0];
  assign nl_MultLoop_acc_2711_nl = conv_s2s_21_22({(data_rsci_idat[323:306]) , 3'b000})
      + conv_s2s_18_22(data_rsci_idat[323:306]) + conv_s2s_16_22(data_rsci_idat[323:308]);
  assign MultLoop_acc_2711_nl = nl_MultLoop_acc_2711_nl[21:0];
  assign nl_MultLoop_acc_1256_nl = conv_s2u_22_24(MultLoop_acc_2711_nl) + conv_s2u_23_24({(data_rsci_idat[323:306])
      , 5'b00000});
  assign MultLoop_acc_1256_nl = nl_MultLoop_acc_1256_nl[23:0];
  assign nl_MultLoop_acc_2713_nl = (~ (data_rsci_idat[197:180])) + conv_s2s_17_18({MultLoop_acc_4191_cse_1
      , (data_rsci_idat[187:182])});
  assign MultLoop_acc_2713_nl = nl_MultLoop_acc_2713_nl[17:0];
  assign nl_MultLoop_acc_2714_nl = ({(data_rsci_idat[197:180]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2713_nl);
  assign MultLoop_acc_2714_nl = nl_MultLoop_acc_2714_nl[19:0];
  assign nl_MultLoop_acc_4271_nl = conv_s2u_14_18(readslicef_20_14_6((MultLoop_acc_2714_nl)))
      + (~ (data_rsci_idat[197:180]));
  assign MultLoop_acc_4271_nl = nl_MultLoop_acc_4271_nl[17:0];
  assign nl_MultLoop_acc_2716_nl = (~ (data_rsci_idat[161:144])) + conv_s2s_16_18({MultLoop_acc_4153_cse_1
      , (data_rsci_idat[151:147])});
  assign MultLoop_acc_2716_nl = nl_MultLoop_acc_2716_nl[17:0];
  assign nl_MultLoop_acc_2717_nl = ({(data_rsci_idat[161:144]) , 2'b01}) + conv_s2s_18_20(MultLoop_acc_2716_nl);
  assign MultLoop_acc_2717_nl = nl_MultLoop_acc_2717_nl[19:0];
  assign nl_MultLoop_acc_531_nl = conv_s2u_20_23(MultLoop_acc_2717_nl) + ({(~ (data_rsci_idat[161:144]))
      , 5'b00000});
  assign MultLoop_acc_531_nl = nl_MultLoop_acc_531_nl[22:0];
  assign nl_MultLoop_acc_2718_nl = (~ (data_rsci_idat[53:36])) + conv_s2s_12_18(data_rsci_idat[53:42]);
  assign MultLoop_acc_2718_nl = nl_MultLoop_acc_2718_nl[17:0];
  assign nl_MultLoop_acc_1252_nl = conv_s2u_18_20(MultLoop_acc_2718_nl) + ({(data_rsci_idat[53:36])
      , 2'b01});
  assign MultLoop_acc_1252_nl = nl_MultLoop_acc_1252_nl[19:0];
  assign nl_MultLoop_acc_2774_itm_1  = conv_s2s_17_18(readslicef_19_17_2((MultLoop_acc_4275_nl)))
      + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_526_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4274_nl)))
      + conv_s2s_16_18(readslicef_24_16_8((MultLoop_acc_1256_nl))) + conv_s2s_16_18(readslicef_18_16_2((MultLoop_acc_4271_nl)))
      + conv_s2s_16_18(readslicef_23_16_7((MultLoop_acc_531_nl))) + conv_s2s_16_18(readslicef_20_16_4((MultLoop_acc_1252_nl)));

  function automatic [9:0] readslicef_18_10_8;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_18_10_8 = tmp[9:0];
  end
  endfunction


  function automatic [10:0] readslicef_18_11_7;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_18_11_7 = tmp[10:0];
  end
  endfunction


  function automatic [11:0] readslicef_18_12_6;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_18_12_6 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_18_13_5;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_18_13_5 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_18_14_4;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_18_14_4 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_18_15_3;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_18_15_3 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_18_16_2;
    input [17:0] vector;
    reg [17:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_18_16_2 = tmp[15:0];
  end
  endfunction


  function automatic [12:0] readslicef_19_13_6;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_19_13_6 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_19_14_5;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_19_14_5 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_19_15_4;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_19_15_4 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_19_16_3;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_19_16_3 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_19_17_2;
    input [18:0] vector;
    reg [18:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_19_17_2 = tmp[16:0];
  end
  endfunction


  function automatic [9:0] readslicef_20_10_10;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_20_10_10 = tmp[9:0];
  end
  endfunction


  function automatic [11:0] readslicef_20_12_8;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_20_12_8 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_20_13_7;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_20_13_7 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_20_14_6;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_20_14_6 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_20_15_5;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_20_15_5 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_20_16_4;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_20_16_4 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_20_17_3;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_20_17_3 = tmp[16:0];
  end
  endfunction


  function automatic [17:0] readslicef_20_18_2;
    input [19:0] vector;
    reg [19:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_20_18_2 = tmp[17:0];
  end
  endfunction


  function automatic [11:0] readslicef_21_12_9;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_21_12_9 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_21_13_8;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_21_13_8 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_21_14_7;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_21_14_7 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_21_15_6;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_21_15_6 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_21_16_5;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_21_16_5 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_21_17_4;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_21_17_4 = tmp[16:0];
  end
  endfunction


  function automatic [18:0] readslicef_21_19_2;
    input [20:0] vector;
    reg [20:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_21_19_2 = tmp[18:0];
  end
  endfunction


  function automatic [11:0] readslicef_22_12_10;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_22_12_10 = tmp[11:0];
  end
  endfunction


  function automatic [12:0] readslicef_22_13_9;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_22_13_9 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_22_14_8;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_22_14_8 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_22_15_7;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_22_15_7 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_22_16_6;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_22_16_6 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_22_17_5;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_22_17_5 = tmp[16:0];
  end
  endfunction


  function automatic [18:0] readslicef_22_19_3;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_22_19_3 = tmp[18:0];
  end
  endfunction


  function automatic [12:0] readslicef_23_13_10;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_23_13_10 = tmp[12:0];
  end
  endfunction


  function automatic [13:0] readslicef_23_14_9;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_23_14_9 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_23_15_8;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_23_15_8 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_23_16_7;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_23_16_7 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_23_17_6;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_23_17_6 = tmp[16:0];
  end
  endfunction


  function automatic [18:0] readslicef_23_19_4;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_23_19_4 = tmp[18:0];
  end
  endfunction


  function automatic [13:0] readslicef_24_14_10;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_24_14_10 = tmp[13:0];
  end
  endfunction


  function automatic [14:0] readslicef_24_15_9;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_24_15_9 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_24_16_8;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_24_16_8 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_24_17_7;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_24_17_7 = tmp[16:0];
  end
  endfunction


  function automatic [14:0] readslicef_25_15_10;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_25_15_10 = tmp[14:0];
  end
  endfunction


  function automatic [15:0] readslicef_25_16_9;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_25_16_9 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_25_17_8;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_25_17_8 = tmp[16:0];
  end
  endfunction


  function automatic [15:0] readslicef_26_16_10;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_26_16_10 = tmp[15:0];
  end
  endfunction


  function automatic [16:0] readslicef_26_17_9;
    input [25:0] vector;
    reg [25:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_26_17_9 = tmp[16:0];
  end
  endfunction


  function automatic [16:0] readslicef_27_17_10;
    input [26:0] vector;
    reg [26:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_27_17_10 = tmp[16:0];
  end
  endfunction


  function automatic [16:0] conv_s2s_8_17 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_17 = {{9{vector[7]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_9_10 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_10 = {vector[8], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_9_12 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_12 = {{3{vector[8]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_9_13 ;
    input [8:0]  vector ;
  begin
    conv_s2s_9_13 = {{4{vector[8]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_10_12 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_12 = {{2{vector[9]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_10_15 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_15 = {{5{vector[9]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_10_16 ;
    input [9:0]  vector ;
  begin
    conv_s2s_10_16 = {{6{vector[9]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_11_15 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_15 = {{4{vector[10]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_11_16 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_16 = {{5{vector[10]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_11_17 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_17 = {{6{vector[10]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2s_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_12_14 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_14 = {{2{vector[11]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_12_15 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_15 = {{3{vector[11]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_12_16 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_16 = {{4{vector[11]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_12_17 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_17 = {{5{vector[11]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_12_19 ;
    input [11:0]  vector ;
  begin
    conv_s2s_12_19 = {{7{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2s_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_13_15 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_15 = {{2{vector[12]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_13_16 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_16 = {{3{vector[12]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_13_17 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_17 = {{4{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_13_19 ;
    input [12:0]  vector ;
  begin
    conv_s2s_13_19 = {{6{vector[12]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2s_14_15 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_15 = {vector[13], vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_14_16 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_16 = {{2{vector[13]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_14_17 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_17 = {{3{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_14_20 ;
    input [13:0]  vector ;
  begin
    conv_s2s_14_20 = {{6{vector[13]}}, vector};
  end
  endfunction


  function automatic [15:0] conv_s2s_15_16 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_16 = {vector[14], vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_15_17 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_17 = {{2{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_15_20 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_20 = {{5{vector[14]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_15_21 ;
    input [14:0]  vector ;
  begin
    conv_s2s_15_21 = {{6{vector[14]}}, vector};
  end
  endfunction


  function automatic [16:0] conv_s2s_16_17 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_17 = {vector[15], vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_16_20 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_20 = {{4{vector[15]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_16_21 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_21 = {{5{vector[15]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_16_22 ;
    input [15:0]  vector ;
  begin
    conv_s2s_16_22 = {{6{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_17_20 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_20 = {{3{vector[16]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_17_21 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_21 = {{4{vector[16]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_17_22 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_22 = {{5{vector[16]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_17_23 ;
    input [16:0]  vector ;
  begin
    conv_s2s_17_23 = {{6{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2s_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_18_26 ;
    input [17:0]  vector ;
  begin
    conv_s2s_18_26 = {{8{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2s_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_19_25 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_25 = {{6{vector[18]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_19_26 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_26 = {{7{vector[18]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_19_27 ;
    input [18:0]  vector ;
  begin
    conv_s2s_19_27 = {{8{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_20_26 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_26 = {{6{vector[19]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_20_27 ;
    input [19:0]  vector ;
  begin
    conv_s2s_20_27 = {{7{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_21_25 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_25 = {{4{vector[20]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_21_26 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_26 = {{5{vector[20]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_21_27 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_27 = {{6{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_22_26 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_26 = {{4{vector[21]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_22_27 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_27 = {{5{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2s_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_23_26 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_26 = {{3{vector[22]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_23_27 ;
    input [22:0]  vector ;
  begin
    conv_s2s_23_27 = {{4{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2s_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_24_26 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_26 = {{2{vector[23]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_24_27 ;
    input [23:0]  vector ;
  begin
    conv_s2s_24_27 = {{3{vector[23]}}, vector};
  end
  endfunction


  function automatic [25:0] conv_s2s_25_26 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_26 = {vector[24], vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_25_27 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_27 = {{2{vector[24]}}, vector};
  end
  endfunction


  function automatic [26:0] conv_s2s_26_27 ;
    input [25:0]  vector ;
  begin
    conv_s2s_26_27 = {vector[25], vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_10_18 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_18 = {{8{vector[9]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_10_19 ;
    input [9:0]  vector ;
  begin
    conv_s2u_10_19 = {{9{vector[9]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_11_18 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_18 = {{7{vector[10]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_11_19 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_19 = {{8{vector[10]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_12_18 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_18 = {{6{vector[11]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_12_19 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_19 = {{7{vector[11]}}, vector};
  end
  endfunction


  function automatic [13:0] conv_s2u_13_14 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_14 = {vector[12], vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_13_18 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_18 = {{5{vector[12]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_13_19 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_19 = {{6{vector[12]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_14_18 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_18 = {{4{vector[13]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_14_19 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_19 = {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_15_18 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_18 = {{3{vector[14]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_15_19 ;
    input [14:0]  vector ;
  begin
    conv_s2u_15_19 = {{4{vector[14]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_16_18 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_18 = {{2{vector[15]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_16_19 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_19 = {{3{vector[15]}}, vector};
  end
  endfunction


  function automatic [17:0] conv_s2u_17_18 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_18 = {vector[16], vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_17_19 ;
    input [16:0]  vector ;
  begin
    conv_s2u_17_19 = {{2{vector[16]}}, vector};
  end
  endfunction


  function automatic [18:0] conv_s2u_18_19 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_19 = {vector[17], vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_18_21 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_21 = {{3{vector[17]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_18_22 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_22 = {{4{vector[17]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_18_23 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_23 = {{5{vector[17]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_18_24 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_24 = {{6{vector[17]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_18_25 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_25 = {{7{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_19_21 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_21 = {{2{vector[18]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_19_22 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_22 = {{3{vector[18]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_19_23 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_23 = {{4{vector[18]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_19_24 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_24 = {{5{vector[18]}}, vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_20_23 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_23 = {{3{vector[19]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_20_24 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_24 = {{4{vector[19]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_20_25 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_25 = {{5{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_21_23 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_23 = {{2{vector[20]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_21_24 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_24 = {{3{vector[20]}}, vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_22_24 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_24 = {{2{vector[21]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_22_25 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_25 = {{3{vector[21]}}, vector};
  end
  endfunction


  function automatic [23:0] conv_s2u_23_24 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_24 = {vector[22], vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_23_25 ;
    input [22:0]  vector ;
  begin
    conv_s2u_23_25 = {{2{vector[22]}}, vector};
  end
  endfunction


  function automatic [24:0] conv_s2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_s2u_24_25 = {vector[23], vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_1_12 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_12 = {{11{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_1_13 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_13 = {{12{1'b0}}, vector};
  end
  endfunction


  function automatic [13:0] conv_u2s_1_14 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_14 = {{13{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_9_11 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_11 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2s_9_13 ;
    input [8:0]  vector ;
  begin
    conv_u2s_9_13 = {{4{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    nnet_dense_large_input_t_layer2_t_config2
// ------------------------------------------------------------------


module nnet_dense_large_input_t_layer2_t_config2 (
  data_rsc_dat, res_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk, ccs_ccore_srst,
      ccs_ccore_en
);
  input [863:0] data_rsc_dat;
  output [431:0] res_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  nnet_dense_large_input_t_layer2_t_config2_core nnet_dense_large_input_t_layer2_t_config2_core_inst
      (
      .data_rsc_dat(data_rsc_dat),
      .res_rsc_z(res_rsc_z),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@fastml02
//  Generated date: Sat Feb  8 11:24:03 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    econV0_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module econV0_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [11:0] fsm_output;
  reg [11:0] fsm_output;


  // FSM State Type Declaration for econV0_core_core_fsm_1
  parameter
    core_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8,
    main_C_8 = 4'd9,
    main_C_9 = 4'd10,
    main_C_10 = 4'd11;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : econV0_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 12'b000000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 12'b000000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 12'b000000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 12'b000000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 12'b000000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 12'b000001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 12'b000010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 12'b000100000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 12'b001000000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 12'b010000000000;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 12'b100000000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 12'b000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_staller
// ------------------------------------------------------------------


module econV0_core_staller (
  clk, rst, core_wen, core_wten, input_48_rsci_wen_comp, layer7_out_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_48_rsci_wen_comp;
  input layer7_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_48_rsci_wen_comp & layer7_out_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_out_1_rsc_triosy_obj_iswt0, const_size_out_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;
  output const_size_out_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsc_triosy_obj_ld_core_sct = const_size_out_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_in_1_rsc_triosy_obj_iswt0, const_size_in_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;
  output const_size_in_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsc_triosy_obj_ld_core_sct = const_size_in_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl (
  core_wten, layer7_out_rsc_triosy_obj_iswt0, layer7_out_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input layer7_out_rsc_triosy_obj_iswt0;
  output layer7_out_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsc_triosy_obj_ld_core_sct = layer7_out_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl (
  core_wten, input_48_rsc_triosy_obj_iswt0, input_48_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input input_48_rsc_triosy_obj_iswt0;
  output input_48_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsc_triosy_obj_ld_core_sct = input_48_rsc_triosy_obj_iswt0 & (~
      core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wten, const_size_out_1_rsci_iswt0, const_size_out_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_out_1_rsci_iswt0;
  output const_size_out_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wten, const_size_in_1_rsci_iswt0, const_size_in_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_in_1_rsci_iswt0;
  output const_size_in_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp (
  clk, rst, layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_biwt,
      layer7_out_rsci_bdwt, layer7_out_rsci_bcwt
);
  input clk;
  input rst;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input layer7_out_rsci_biwt;
  input layer7_out_rsci_bdwt;
  output layer7_out_rsci_bcwt;
  reg layer7_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_wen_comp = (~ layer7_out_rsci_oswt) | layer7_out_rsci_biwt
      | layer7_out_rsci_bcwt;
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_bcwt <= 1'b0;
    end
    else begin
      layer7_out_rsci_bcwt <= ~((~(layer7_out_rsci_bcwt | layer7_out_rsci_biwt))
          | layer7_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl (
  core_wen, layer7_out_rsci_oswt, layer7_out_rsci_irdy, layer7_out_rsci_biwt, layer7_out_rsci_bdwt,
      layer7_out_rsci_bcwt, layer7_out_rsci_ivld_core_sct
);
  input core_wen;
  input layer7_out_rsci_oswt;
  input layer7_out_rsci_irdy;
  output layer7_out_rsci_biwt;
  output layer7_out_rsci_bdwt;
  input layer7_out_rsci_bcwt;
  output layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire layer7_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign layer7_out_rsci_bdwt = layer7_out_rsci_oswt & core_wen;
  assign layer7_out_rsci_biwt = layer7_out_rsci_ogwt & layer7_out_rsci_irdy;
  assign layer7_out_rsci_ogwt = layer7_out_rsci_oswt & (~ layer7_out_rsci_bcwt);
  assign layer7_out_rsci_ivld_core_sct = layer7_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci_input_48_rsc_wait_dp
// ------------------------------------------------------------------


module econV0_core_input_48_rsci_input_48_rsc_wait_dp (
  clk, rst, input_48_rsci_oswt, input_48_rsci_wen_comp, input_48_rsci_idat_mxwt,
      input_48_rsci_biwt, input_48_rsci_bdwt, input_48_rsci_bcwt, input_48_rsci_idat
);
  input clk;
  input rst;
  input input_48_rsci_oswt;
  output input_48_rsci_wen_comp;
  output [863:0] input_48_rsci_idat_mxwt;
  input input_48_rsci_biwt;
  input input_48_rsci_bdwt;
  output input_48_rsci_bcwt;
  reg input_48_rsci_bcwt;
  input [863:0] input_48_rsci_idat;


  // Interconnect Declarations
  reg [863:0] input_48_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsci_wen_comp = (~ input_48_rsci_oswt) | input_48_rsci_biwt | input_48_rsci_bcwt;
  assign input_48_rsci_idat_mxwt = MUX_v_864_2_2(input_48_rsci_idat, input_48_rsci_idat_bfwt,
      input_48_rsci_bcwt);
  always @(posedge clk) begin
    if ( rst ) begin
      input_48_rsci_bcwt <= 1'b0;
      input_48_rsci_idat_bfwt <= 864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else begin
      input_48_rsci_bcwt <= ~((~(input_48_rsci_bcwt | input_48_rsci_biwt)) | input_48_rsci_bdwt);
      input_48_rsci_idat_bfwt <= input_48_rsci_idat_mxwt;
    end
  end

  function automatic [863:0] MUX_v_864_2_2;
    input [863:0] input_0;
    input [863:0] input_1;
    input [0:0] sel;
    reg [863:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_864_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci_input_48_rsc_wait_ctrl
// ------------------------------------------------------------------


module econV0_core_input_48_rsci_input_48_rsc_wait_ctrl (
  core_wen, input_48_rsci_oswt, input_48_rsci_biwt, input_48_rsci_bdwt, input_48_rsci_bcwt,
      input_48_rsci_irdy_core_sct, input_48_rsci_ivld
);
  input core_wen;
  input input_48_rsci_oswt;
  output input_48_rsci_biwt;
  output input_48_rsci_bdwt;
  input input_48_rsci_bcwt;
  output input_48_rsci_irdy_core_sct;
  input input_48_rsci_ivld;


  // Interconnect Declarations
  wire input_48_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign input_48_rsci_bdwt = input_48_rsci_oswt & core_wen;
  assign input_48_rsci_biwt = input_48_rsci_ogwt & input_48_rsci_ivld;
  assign input_48_rsci_ogwt = input_48_rsci_oswt & (~ input_48_rsci_bcwt);
  assign input_48_rsci_irdy_core_sct = input_48_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsc_triosy_obj (
  const_size_out_1_rsc_triosy_lz, core_wten, const_size_out_1_rsc_triosy_obj_iswt0
);
  output const_size_out_1_rsc_triosy_lz;
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_out_1_rsc_triosy_obj (
      .ld(const_size_out_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_out_1_rsc_triosy_lz)
    );
  econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
      econV0_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(const_size_out_1_rsc_triosy_obj_iswt0),
      .const_size_out_1_rsc_triosy_obj_ld_core_sct(const_size_out_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsc_triosy_obj (
  const_size_in_1_rsc_triosy_lz, core_wten, const_size_in_1_rsc_triosy_obj_iswt0
);
  output const_size_in_1_rsc_triosy_lz;
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_in_1_rsc_triosy_obj (
      .ld(const_size_in_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_in_1_rsc_triosy_lz)
    );
  econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
      econV0_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(const_size_in_1_rsc_triosy_obj_iswt0),
      .const_size_in_1_rsc_triosy_obj_ld_core_sct(const_size_in_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsc_triosy_obj (
  layer7_out_rsc_triosy_lz, core_wten, layer7_out_rsc_triosy_obj_iswt0
);
  output layer7_out_rsc_triosy_lz;
  input core_wten;
  input layer7_out_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire layer7_out_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) layer7_out_rsc_triosy_obj (
      .ld(layer7_out_rsc_triosy_obj_ld_core_sct),
      .lz(layer7_out_rsc_triosy_lz)
    );
  econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl econV0_core_layer7_out_rsc_triosy_obj_layer7_out_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer7_out_rsc_triosy_obj_iswt0(layer7_out_rsc_triosy_obj_iswt0),
      .layer7_out_rsc_triosy_obj_ld_core_sct(layer7_out_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsc_triosy_obj
// ------------------------------------------------------------------


module econV0_core_input_48_rsc_triosy_obj (
  input_48_rsc_triosy_lz, core_wten, input_48_rsc_triosy_obj_iswt0
);
  output input_48_rsc_triosy_lz;
  input core_wten;
  input input_48_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire input_48_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) input_48_rsc_triosy_obj (
      .ld(input_48_rsc_triosy_obj_ld_core_sct),
      .lz(input_48_rsc_triosy_lz)
    );
  econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl econV0_core_input_48_rsc_triosy_obj_input_48_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .input_48_rsc_triosy_obj_iswt0(input_48_rsc_triosy_obj_iswt0),
      .input_48_rsc_triosy_obj_ld_core_sct(input_48_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module econV0_core_const_size_out_1_rsci (
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, core_wten, const_size_out_1_rsci_iswt0
);
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input core_wten;
  input const_size_out_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd25),
  .width(32'sd16)) const_size_out_1_rsci (
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000000011),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl econV0_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(const_size_out_1_rsci_iswt0),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module econV0_core_const_size_in_1_rsci (
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, core_wten, const_size_in_1_rsci_iswt0
);
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input core_wten;
  input const_size_in_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd24),
  .width(32'sd16)) const_size_in_1_rsci (
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000110000),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl econV0_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(const_size_in_1_rsci_iswt0),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_layer7_out_rsci
// ------------------------------------------------------------------


module econV0_core_layer7_out_rsci (
  clk, rst, layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, core_wen,
      layer7_out_rsci_oswt, layer7_out_rsci_wen_comp, layer7_out_rsci_idat
);
  input clk;
  input rst;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  input core_wen;
  input layer7_out_rsci_oswt;
  output layer7_out_rsci_wen_comp;
  input [53:0] layer7_out_rsci_idat;


  // Interconnect Declarations
  wire layer7_out_rsci_irdy;
  wire layer7_out_rsci_biwt;
  wire layer7_out_rsci_bdwt;
  wire layer7_out_rsci_bcwt;
  wire layer7_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd23),
  .width(32'sd54)) layer7_out_rsci (
      .irdy(layer7_out_rsci_irdy),
      .ivld(layer7_out_rsci_ivld_core_sct),
      .idat(layer7_out_rsci_idat),
      .rdy(layer7_out_rsc_rdy),
      .vld(layer7_out_rsc_vld),
      .dat(layer7_out_rsc_dat)
    );
  econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl econV0_core_layer7_out_rsci_layer7_out_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_irdy(layer7_out_rsci_irdy),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt),
      .layer7_out_rsci_ivld_core_sct(layer7_out_rsci_ivld_core_sct)
    );
  econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp econV0_core_layer7_out_rsci_layer7_out_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsci_oswt(layer7_out_rsci_oswt),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_biwt(layer7_out_rsci_biwt),
      .layer7_out_rsci_bdwt(layer7_out_rsci_bdwt),
      .layer7_out_rsci_bcwt(layer7_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core_input_48_rsci
// ------------------------------------------------------------------


module econV0_core_input_48_rsci (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, core_wen, input_48_rsci_oswt,
      input_48_rsci_wen_comp, input_48_rsci_idat_mxwt
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  input core_wen;
  input input_48_rsci_oswt;
  output input_48_rsci_wen_comp;
  output [863:0] input_48_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_48_rsci_biwt;
  wire input_48_rsci_bdwt;
  wire input_48_rsci_bcwt;
  wire input_48_rsci_irdy_core_sct;
  wire input_48_rsci_ivld;
  wire [863:0] input_48_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd22),
  .width(32'sd864)) input_48_rsci (
      .rdy(input_48_rsc_rdy),
      .vld(input_48_rsc_vld),
      .dat(input_48_rsc_dat),
      .irdy(input_48_rsci_irdy_core_sct),
      .ivld(input_48_rsci_ivld),
      .idat(input_48_rsci_idat)
    );
  econV0_core_input_48_rsci_input_48_rsc_wait_ctrl econV0_core_input_48_rsci_input_48_rsc_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .input_48_rsci_oswt(input_48_rsci_oswt),
      .input_48_rsci_biwt(input_48_rsci_biwt),
      .input_48_rsci_bdwt(input_48_rsci_bdwt),
      .input_48_rsci_bcwt(input_48_rsci_bcwt),
      .input_48_rsci_irdy_core_sct(input_48_rsci_irdy_core_sct),
      .input_48_rsci_ivld(input_48_rsci_ivld)
    );
  econV0_core_input_48_rsci_input_48_rsc_wait_dp econV0_core_input_48_rsci_input_48_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .input_48_rsci_oswt(input_48_rsci_oswt),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .input_48_rsci_idat_mxwt(input_48_rsci_idat_mxwt),
      .input_48_rsci_biwt(input_48_rsci_biwt),
      .input_48_rsci_bdwt(input_48_rsci_bdwt),
      .input_48_rsci_bcwt(input_48_rsci_bcwt),
      .input_48_rsci_idat(input_48_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0_core
// ------------------------------------------------------------------


module econV0_core (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, input_48_rsc_triosy_lz,
      layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, layer7_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_triosy_lz,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  output input_48_rsc_triosy_lz;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output layer7_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_48_rsci_wen_comp;
  wire [863:0] input_48_rsci_idat_mxwt;
  wire layer7_out_rsci_wen_comp;
  reg [53:0] layer7_out_rsci_idat;
  wire [53:0] nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z;
  wire [53:0] nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z;
  wire [107:0] nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z;
  wire [107:0] nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z;
  wire [431:0] nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z;
  wire [431:0] nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z;
  wire [11:0] fsm_output;
  reg reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse;
  reg [107:0] nnet_dense_large_layer5_t_layer6_t_config6_layer5_out_sva;
  reg [431:0] nnet_dense_large_layer3_t_layer4_t_config4_layer3_out_sva;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[9];
  wire [107:0] nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_data_rsc_dat;
  assign nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_data_rsc_dat = nnet_dense_large_layer5_t_layer6_t_config6_layer5_out_sva;
  wire [0:0] nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[8];
  wire [0:0] nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[6];
  wire [431:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_data_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_data_rsc_dat = nnet_dense_large_layer3_t_layer4_t_config4_layer3_out_sva;
  wire [0:0] nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[5];
  wire [0:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[3];
  wire [0:0] nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat;
  assign nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat
      = fsm_output[1];
  nnet_relu_layer6_t_result_t_relu_config7  nnet_relu_layer6_t_result_t_relu_config7_cmp
      (
      .data_rsc_dat(nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer6_t_result_t_relu_config7_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_layer5_t_layer6_t_config6  nnet_dense_large_layer5_t_layer6_t_config6_cmp
      (
      .data_rsc_dat(nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_data_rsc_dat[107:0]),
      .res_rsc_z(nnet_dense_large_layer5_t_layer6_t_config6_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_layer5_t_layer6_t_config6_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_relu_layer4_t_layer5_t_relu_config5  nnet_relu_layer4_t_layer5_t_relu_config5_cmp
      (
      .data_rsc_dat(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer4_t_layer5_t_relu_config5_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_layer3_t_layer4_t_config4  nnet_dense_large_layer3_t_layer4_t_config4_cmp
      (
      .data_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_data_rsc_dat[431:0]),
      .res_rsc_z(nnet_dense_large_layer3_t_layer4_t_config4_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_layer3_t_layer4_t_config4_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_relu_layer2_t_layer3_t_relu_config3  nnet_relu_layer2_t_layer3_t_relu_config3_cmp
      (
      .data_rsc_dat(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .res_rsc_z(nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_relu_layer2_t_layer3_t_relu_config3_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  nnet_dense_large_input_t_layer2_t_config2  nnet_dense_large_input_t_layer2_t_config2_cmp
      (
      .data_rsc_dat(input_48_rsci_idat_mxwt),
      .res_rsc_z(nnet_dense_large_input_t_layer2_t_config2_cmp_res_rsc_z),
      .ccs_ccore_clk(clk),
      .ccs_ccore_en(core_wen),
      .ccs_ccore_srst(rst),
      .ccs_ccore_start_rsc_dat(nl_nnet_dense_large_input_t_layer2_t_config2_cmp_ccs_ccore_start_rsc_dat[0:0])
    );
  econV0_core_input_48_rsci econV0_core_input_48_rsci_inst (
      .clk(clk),
      .rst(rst),
      .input_48_rsc_dat(input_48_rsc_dat),
      .input_48_rsc_vld(input_48_rsc_vld),
      .input_48_rsc_rdy(input_48_rsc_rdy),
      .core_wen(core_wen),
      .input_48_rsci_oswt(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .input_48_rsci_idat_mxwt(input_48_rsci_idat_mxwt)
    );
  econV0_core_layer7_out_rsci econV0_core_layer7_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .core_wen(core_wen),
      .layer7_out_rsci_oswt(reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp),
      .layer7_out_rsci_idat(layer7_out_rsci_idat)
    );
  econV0_core_const_size_in_1_rsci econV0_core_const_size_in_1_rsci_inst (
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_out_1_rsci econV0_core_const_size_out_1_rsci_inst (
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_input_48_rsc_triosy_obj econV0_core_input_48_rsc_triosy_obj_inst (
      .input_48_rsc_triosy_lz(input_48_rsc_triosy_lz),
      .core_wten(core_wten),
      .input_48_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_layer7_out_rsc_triosy_obj econV0_core_layer7_out_rsc_triosy_obj_inst
      (
      .layer7_out_rsc_triosy_lz(layer7_out_rsc_triosy_lz),
      .core_wten(core_wten),
      .layer7_out_rsc_triosy_obj_iswt0(reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_in_1_rsc_triosy_obj econV0_core_const_size_in_1_rsc_triosy_obj_inst
      (
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_const_size_out_1_rsc_triosy_obj econV0_core_const_size_out_1_rsc_triosy_obj_inst
      (
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse)
    );
  econV0_core_staller econV0_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_48_rsci_wen_comp(input_48_rsci_wen_comp),
      .layer7_out_rsci_wen_comp(layer7_out_rsci_wen_comp)
    );
  econV0_core_core_fsm econV0_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  always @(posedge clk) begin
    if ( rst ) begin
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      nnet_dense_large_layer3_t_layer4_t_config4_layer3_out_sva <= 432'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nnet_dense_large_layer5_t_layer6_t_config6_layer5_out_sva <= 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen ) begin
      reg_const_size_out_1_rsc_triosy_obj_ld_core_psct_cse <= (fsm_output[11]) |
          (fsm_output[0]);
      reg_layer7_out_rsc_triosy_obj_ld_core_psct_cse <= fsm_output[10];
      nnet_dense_large_layer3_t_layer4_t_config4_layer3_out_sva <= nnet_relu_layer2_t_layer3_t_relu_config3_cmp_res_rsc_z;
      nnet_dense_large_layer5_t_layer6_t_config6_layer5_out_sva <= nnet_relu_layer4_t_layer5_t_relu_config5_cmp_res_rsc_z;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      layer7_out_rsci_idat <= 54'b000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (fsm_output[10]) ) begin
      layer7_out_rsci_idat <= nnet_relu_layer6_t_result_t_relu_config7_cmp_res_rsc_z;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econV0
// ------------------------------------------------------------------


module econV0 (
  clk, rst, input_48_rsc_dat, input_48_rsc_vld, input_48_rsc_rdy, input_48_rsc_triosy_lz,
      layer7_out_rsc_dat, layer7_out_rsc_vld, layer7_out_rsc_rdy, layer7_out_rsc_triosy_lz,
      const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, const_size_in_1_rsc_triosy_lz,
      const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, const_size_out_1_rsc_triosy_lz
);
  input clk;
  input rst;
  input [863:0] input_48_rsc_dat;
  input input_48_rsc_vld;
  output input_48_rsc_rdy;
  output input_48_rsc_triosy_lz;
  output [53:0] layer7_out_rsc_dat;
  output layer7_out_rsc_vld;
  input layer7_out_rsc_rdy;
  output layer7_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  econV0_core econV0_core_inst (
      .clk(clk),
      .rst(rst),
      .input_48_rsc_dat(input_48_rsc_dat),
      .input_48_rsc_vld(input_48_rsc_vld),
      .input_48_rsc_rdy(input_48_rsc_rdy),
      .input_48_rsc_triosy_lz(input_48_rsc_triosy_lz),
      .layer7_out_rsc_dat(layer7_out_rsc_dat),
      .layer7_out_rsc_vld(layer7_out_rsc_vld),
      .layer7_out_rsc_rdy(layer7_out_rsc_rdy),
      .layer7_out_rsc_triosy_lz(layer7_out_rsc_triosy_lz),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz)
    );
endmodule



