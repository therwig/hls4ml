
//------> /opt/cad/catapult/pkgs/siflibs/ccs_in_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This doocument may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_vld_v1 (idat, ivld, dat, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             ivld;
  input  [width-1:0] dat;
  input              vld;

  wire   [width-1:0] idat;
  wire               ivld;

  assign idat = dat;
  assign ivld = vld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/ccs_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_vld_v1 (dat, vld, idat, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             vld;
  input  [width-1:0] idat;
  input              ivld;

  wire   [width-1:0] dat;
  wire               vld;

  assign dat = idat;
  assign vld = ivld;

endmodule


//------> /opt/cad/catapult/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4c/853139 Production Release
//  HLS Date:       Thu Jan 16 19:19:57 PST 2020
// 
//  Generated by:   giuseppe@gandalf
//  Generated date: Tue Mar  3 18:40:33 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module econ_4x4_d10_core_core_fsm (
  clk, rst, core_wen, fsm_output
);
  input clk;
  input rst;
  input core_wen;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;


  // FSM State Type Declaration for econ_4x4_d10_core_core_fsm_1
  parameter
    core_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    main_C_5 = 4'd6,
    main_C_6 = 4'd7,
    main_C_7 = 4'd8,
    main_C_8 = 4'd9;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : econ_4x4_d10_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 10'b0000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_staller
// ------------------------------------------------------------------


module econ_4x4_d10_core_staller (
  clk, rst, core_wen, core_wten, input_1_rsci_wen_comp, w2_rsci_wen_comp, b2_rsci_wen_comp,
      w4_rsci_wen_comp, b4_rsci_wen_comp
);
  input clk;
  input rst;
  output core_wen;
  output core_wten;
  reg core_wten;
  input input_1_rsci_wen_comp;
  input w2_rsci_wen_comp;
  input b2_rsci_wen_comp;
  input w4_rsci_wen_comp;
  input b4_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = input_1_rsci_wen_comp & w2_rsci_wen_comp & b2_rsci_wen_comp &
      w4_rsci_wen_comp & b4_rsci_wen_comp;
  always @(posedge clk) begin
    if ( rst ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl (
  core_wten, b4_rsc_triosy_obj_iswt0, b4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;
  output b4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b4_rsc_triosy_obj_ld_core_sct = b4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl (
  core_wten, w4_rsc_triosy_obj_iswt0, w4_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;
  output w4_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w4_rsc_triosy_obj_ld_core_sct = w4_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl (
  core_wten, b2_rsc_triosy_obj_iswt0, b2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;
  output b2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign b2_rsc_triosy_obj_ld_core_sct = b2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl (
  core_wten, w2_rsc_triosy_obj_iswt0, w2_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;
  output w2_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign w2_rsc_triosy_obj_ld_core_sct = w2_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_out_1_rsc_triosy_obj_iswt0, const_size_out_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;
  output const_size_out_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsc_triosy_obj_ld_core_sct = const_size_out_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
    (
  core_wten, const_size_in_1_rsc_triosy_obj_iswt0, const_size_in_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;
  output const_size_in_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsc_triosy_obj_ld_core_sct = const_size_in_1_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl
    (
  core_wten, layer5_out_rsc_triosy_obj_iswt0, layer5_out_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;
  output layer5_out_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsc_triosy_obj_ld_core_sct = layer5_out_rsc_triosy_obj_iswt0
      & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl (
  core_wten, input_1_rsc_triosy_obj_iswt0, input_1_rsc_triosy_obj_ld_core_sct
);
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;
  output input_1_rsc_triosy_obj_ld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign input_1_rsc_triosy_obj_ld_core_sct = input_1_rsc_triosy_obj_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsci (
  b4_rsc_dat, b4_rsc_vld, b4_rsci_oswt, b4_rsci_wen_comp, b4_rsci_idat_mxwt
);
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  input b4_rsci_oswt;
  output b4_rsci_wen_comp;
  output [79:0] b4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b4_rsci_ivld;
  wire [79:0] b4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd8),
  .width(32'sd80)) b4_rsci (
      .vld(b4_rsc_vld),
      .dat(b4_rsc_dat),
      .ivld(b4_rsci_ivld),
      .idat(b4_rsci_idat)
    );
  assign b4_rsci_idat_mxwt = b4_rsci_idat;
  assign b4_rsci_wen_comp = (~ b4_rsci_oswt) | b4_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsci (
  w4_rsc_dat, w4_rsc_vld, w4_rsci_oswt, w4_rsci_wen_comp, w4_rsci_idat_mxwt
);
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  input w4_rsci_oswt;
  output w4_rsci_wen_comp;
  output [10239:0] w4_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w4_rsci_ivld;
  wire [10239:0] w4_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd7),
  .width(32'sd10240)) w4_rsci (
      .vld(w4_rsc_vld),
      .dat(w4_rsc_dat),
      .ivld(w4_rsci_ivld),
      .idat(w4_rsci_idat)
    );
  assign w4_rsci_idat_mxwt = w4_rsci_idat;
  assign w4_rsci_wen_comp = (~ w4_rsci_oswt) | w4_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsci (
  b2_rsc_dat, b2_rsc_vld, b2_rsci_oswt, b2_rsci_wen_comp, b2_rsci_idat_mxwt
);
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  input b2_rsci_oswt;
  output b2_rsci_wen_comp;
  output [63:0] b2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b2_rsci_ivld;
  wire [63:0] b2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd6),
  .width(32'sd64)) b2_rsci (
      .vld(b2_rsc_vld),
      .dat(b2_rsc_dat),
      .ivld(b2_rsci_ivld),
      .idat(b2_rsci_idat)
    );
  assign b2_rsci_idat_mxwt = b2_rsci_idat;
  assign b2_rsci_wen_comp = (~ b2_rsci_oswt) | b2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsci (
  w2_rsc_dat, w2_rsc_vld, w2_rsci_oswt, w2_rsci_wen_comp, w2_rsci_idat_mxwt
);
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  input w2_rsci_oswt;
  output w2_rsci_wen_comp;
  output [1727:0] w2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire w2_rsci_ivld;
  wire [1727:0] w2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd5),
  .width(32'sd1728)) w2_rsci (
      .vld(w2_rsc_vld),
      .dat(w2_rsc_dat),
      .ivld(w2_rsci_ivld),
      .idat(w2_rsci_idat)
    );
  assign w2_rsci_idat_mxwt = w2_rsci_idat;
  assign w2_rsci_wen_comp = (~ w2_rsci_oswt) | w2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl (
  core_wten, const_size_out_1_rsci_iswt0, const_size_out_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_out_1_rsci_iswt0;
  output const_size_out_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_out_1_rsci_ivld_core_sct = const_size_out_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl (
  core_wten, const_size_in_1_rsci_iswt0, const_size_in_1_rsci_ivld_core_sct
);
  input core_wten;
  input const_size_in_1_rsci_iswt0;
  output const_size_in_1_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign const_size_in_1_rsci_ivld_core_sct = const_size_in_1_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl (
  core_wten, layer5_out_rsci_iswt0, layer5_out_rsci_ivld_core_sct
);
  input core_wten;
  input layer5_out_rsci_iswt0;
  output layer5_out_rsci_ivld_core_sct;



  // Interconnect Declarations for Component Instantiations 
  assign layer5_out_rsci_ivld_core_sct = layer5_out_rsci_iswt0 & (~ core_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsci (
  input_1_rsc_dat, input_1_rsc_vld, input_1_rsci_oswt, input_1_rsci_wen_comp, input_1_rsci_idat_mxwt
);
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  input input_1_rsci_oswt;
  output input_1_rsci_wen_comp;
  output [1055:0] input_1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire input_1_rsci_ivld;
  wire [1055:0] input_1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_vld_v1 #(.rscid(32'sd1),
  .width(32'sd1056)) input_1_rsci (
      .vld(input_1_rsc_vld),
      .dat(input_1_rsc_dat),
      .ivld(input_1_rsci_ivld),
      .idat(input_1_rsci_idat)
    );
  assign input_1_rsci_idat_mxwt = input_1_rsci_idat;
  assign input_1_rsci_wen_comp = (~ input_1_rsci_oswt) | input_1_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b4_rsc_triosy_obj (
  b4_rsc_triosy_lz, core_wten, b4_rsc_triosy_obj_iswt0
);
  output b4_rsc_triosy_lz;
  input core_wten;
  input b4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b4_rsc_triosy_obj (
      .ld(b4_rsc_triosy_obj_ld_core_sct),
      .lz(b4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl econ_4x4_d10_core_b4_rsc_triosy_obj_b4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(b4_rsc_triosy_obj_iswt0),
      .b4_rsc_triosy_obj_ld_core_sct(b4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w4_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w4_rsc_triosy_obj (
  w4_rsc_triosy_lz, core_wten, w4_rsc_triosy_obj_iswt0
);
  output w4_rsc_triosy_lz;
  input core_wten;
  input w4_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w4_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w4_rsc_triosy_obj (
      .ld(w4_rsc_triosy_obj_ld_core_sct),
      .lz(w4_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl econ_4x4_d10_core_w4_rsc_triosy_obj_w4_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(w4_rsc_triosy_obj_iswt0),
      .w4_rsc_triosy_obj_ld_core_sct(w4_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_b2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_b2_rsc_triosy_obj (
  b2_rsc_triosy_lz, core_wten, b2_rsc_triosy_obj_iswt0
);
  output b2_rsc_triosy_lz;
  input core_wten;
  input b2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire b2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) b2_rsc_triosy_obj (
      .ld(b2_rsc_triosy_obj_ld_core_sct),
      .lz(b2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl econ_4x4_d10_core_b2_rsc_triosy_obj_b2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(b2_rsc_triosy_obj_iswt0),
      .b2_rsc_triosy_obj_ld_core_sct(b2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_w2_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_w2_rsc_triosy_obj (
  w2_rsc_triosy_lz, core_wten, w2_rsc_triosy_obj_iswt0
);
  output w2_rsc_triosy_lz;
  input core_wten;
  input w2_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire w2_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) w2_rsc_triosy_obj (
      .ld(w2_rsc_triosy_obj_ld_core_sct),
      .lz(w2_rsc_triosy_lz)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl econ_4x4_d10_core_w2_rsc_triosy_obj_w2_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(w2_rsc_triosy_obj_iswt0),
      .w2_rsc_triosy_obj_ld_core_sct(w2_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj (
  const_size_out_1_rsc_triosy_lz, core_wten, const_size_out_1_rsc_triosy_obj_iswt0
);
  output const_size_out_1_rsc_triosy_lz;
  input core_wten;
  input const_size_out_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_out_1_rsc_triosy_obj (
      .ld(const_size_out_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_out_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_const_size_out_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(const_size_out_1_rsc_triosy_obj_iswt0),
      .const_size_out_1_rsc_triosy_obj_ld_core_sct(const_size_out_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj (
  const_size_in_1_rsc_triosy_lz, core_wten, const_size_in_1_rsc_triosy_obj_iswt0
);
  output const_size_in_1_rsc_triosy_lz;
  input core_wten;
  input const_size_in_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) const_size_in_1_rsc_triosy_obj (
      .ld(const_size_in_1_rsc_triosy_obj_ld_core_sct),
      .lz(const_size_in_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl
      econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_const_size_in_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(const_size_in_1_rsc_triosy_obj_iswt0),
      .const_size_in_1_rsc_triosy_obj_ld_core_sct(const_size_in_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsc_triosy_obj (
  layer5_out_rsc_triosy_lz, core_wten, layer5_out_rsc_triosy_obj_iswt0
);
  output layer5_out_rsc_triosy_lz;
  input core_wten;
  input layer5_out_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire layer5_out_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) layer5_out_rsc_triosy_obj (
      .ld(layer5_out_rsc_triosy_obj_ld_core_sct),
      .lz(layer5_out_rsc_triosy_lz)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl econ_4x4_d10_core_layer5_out_rsc_triosy_obj_layer5_out_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(layer5_out_rsc_triosy_obj_iswt0),
      .layer5_out_rsc_triosy_obj_ld_core_sct(layer5_out_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_input_1_rsc_triosy_obj
// ------------------------------------------------------------------


module econ_4x4_d10_core_input_1_rsc_triosy_obj (
  input_1_rsc_triosy_lz, core_wten, input_1_rsc_triosy_obj_iswt0
);
  output input_1_rsc_triosy_lz;
  input core_wten;
  input input_1_rsc_triosy_obj_iswt0;


  // Interconnect Declarations
  wire input_1_rsc_triosy_obj_ld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  mgc_io_sync_v2 #(.valid(32'sd0)) input_1_rsc_triosy_obj (
      .ld(input_1_rsc_triosy_obj_ld_core_sct),
      .lz(input_1_rsc_triosy_lz)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl econ_4x4_d10_core_input_1_rsc_triosy_obj_input_1_rsc_triosy_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(input_1_rsc_triosy_obj_iswt0),
      .input_1_rsc_triosy_obj_ld_core_sct(input_1_rsc_triosy_obj_ld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_out_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_out_1_rsci (
  const_size_out_1_rsc_dat, const_size_out_1_rsc_vld, core_wten, const_size_out_1_rsci_iswt0
);
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  input core_wten;
  input const_size_out_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_out_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd4),
  .width(32'sd16)) const_size_out_1_rsci (
      .ivld(const_size_out_1_rsci_ivld_core_sct),
      .idat(16'b0000000000001010),
      .vld(const_size_out_1_rsc_vld),
      .dat(const_size_out_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_out_1_rsci_const_size_out_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(const_size_out_1_rsci_iswt0),
      .const_size_out_1_rsci_ivld_core_sct(const_size_out_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_const_size_in_1_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_const_size_in_1_rsci (
  const_size_in_1_rsc_dat, const_size_in_1_rsc_vld, core_wten, const_size_in_1_rsci_iswt0
);
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  input core_wten;
  input const_size_in_1_rsci_iswt0;


  // Interconnect Declarations
  wire const_size_in_1_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_vld_v1 #(.rscid(32'sd3),
  .width(32'sd16)) const_size_in_1_rsci (
      .ivld(const_size_in_1_rsci_ivld_core_sct),
      .idat(16'b0000000000110000),
      .vld(const_size_in_1_rsc_vld),
      .dat(const_size_in_1_rsc_dat)
    );
  econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl econ_4x4_d10_core_const_size_in_1_rsci_const_size_in_1_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(const_size_in_1_rsci_iswt0),
      .const_size_in_1_rsci_ivld_core_sct(const_size_in_1_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core_layer5_out_rsci
// ------------------------------------------------------------------


module econ_4x4_d10_core_layer5_out_rsci (
  layer5_out_rsc_dat, layer5_out_rsc_vld, core_wten, layer5_out_rsci_iswt0, layer5_out_rsci_idat
);
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  input core_wten;
  input layer5_out_rsci_iswt0;
  input [219:0] layer5_out_rsci_idat;


  // Interconnect Declarations
  wire layer5_out_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [219:0] nl_layer5_out_rsci_idat;
  assign nl_layer5_out_rsci_idat = {1'b0 , (layer5_out_rsci_idat[218:198]) , 1'b0
      , (layer5_out_rsci_idat[196:176]) , 1'b0 , (layer5_out_rsci_idat[174:154])
      , 1'b0 , (layer5_out_rsci_idat[152:132]) , 1'b0 , (layer5_out_rsci_idat[130:110])
      , 1'b0 , (layer5_out_rsci_idat[108:88]) , 1'b0 , (layer5_out_rsci_idat[86:66])
      , 1'b0 , (layer5_out_rsci_idat[64:44]) , 1'b0 , (layer5_out_rsci_idat[42:22])
      , 1'b0 , (layer5_out_rsci_idat[20:0])};
  ccs_out_vld_v1 #(.rscid(32'sd2),
  .width(32'sd220)) layer5_out_rsci (
      .ivld(layer5_out_rsci_ivld_core_sct),
      .idat(nl_layer5_out_rsci_idat[219:0]),
      .vld(layer5_out_rsc_vld),
      .dat(layer5_out_rsc_dat)
    );
  econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl econ_4x4_d10_core_layer5_out_rsci_layer5_out_rsc_wait_ctrl_inst
      (
      .core_wten(core_wten),
      .layer5_out_rsci_iswt0(layer5_out_rsci_iswt0),
      .layer5_out_rsci_ivld_core_sct(layer5_out_rsci_ivld_core_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10_core
// ------------------------------------------------------------------


module econ_4x4_d10_core (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_triosy_lz, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_triosy_lz, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld, w2_rsc_triosy_lz, b2_rsc_dat,
      b2_rsc_vld, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_triosy_lz, b4_rsc_dat,
      b4_rsc_vld, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_triosy_lz;
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_triosy_lz;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire input_1_rsci_wen_comp;
  wire [1055:0] input_1_rsci_idat_mxwt;
  wire w2_rsci_wen_comp;
  wire [1727:0] w2_rsci_idat_mxwt;
  wire b2_rsci_wen_comp;
  wire [63:0] b2_rsci_idat_mxwt;
  wire w4_rsci_wen_comp;
  wire [10239:0] w4_rsci_idat_mxwt;
  wire b4_rsci_wen_comp;
  wire [79:0] b4_rsci_idat_mxwt;
  reg [20:0] layer5_out_rsci_idat_196_176;
  reg [20:0] layer5_out_rsci_idat_174_154;
  reg [20:0] layer5_out_rsci_idat_152_132;
  reg [20:0] layer5_out_rsci_idat_130_110;
  reg [20:0] layer5_out_rsci_idat_108_88;
  reg [20:0] layer5_out_rsci_idat_86_66;
  reg [20:0] layer5_out_rsci_idat_64_44;
  reg [20:0] layer5_out_rsci_idat_42_22;
  reg [20:0] layer5_out_rsci_idat_20_0;
  reg [20:0] layer5_out_rsci_idat_218_198;
  wire [9:0] fsm_output;
  wire [21:0] AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [22:0] nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [22:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1;
  wire [21:0] nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire [22:0] nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1;
  wire layer5_out_and_cse;
  reg reg_b4_rsc_triosy_obj_ld_core_psct_cse;
  reg reg_layer5_out_rsc_triosy_obj_ld_core_psct_cse;
  wire InitAccum_and_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_1_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_cse;
  wire AccumDotWidth_and_5_cse;
  wire AccumDotWidth_and_7_cse;
  wire AccumDotWidth_and_3_cse;
  wire AccumDotWidth_and_10_cse;
  wire MultLoop_and_2_cse;
  wire AccumDotWidth_and_8_cse;
  wire MultLoop_and_4_cse;
  wire MultLoop_and_11_cse;
  wire MultLoop_and_1_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_10_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_29_cse;
  wire AccumDotWidth_and_25_cse;
  wire MultLoop_and_35_cse;
  wire AccumDotWidth_and_26_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_11_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_32_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_34_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_31_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_47_cse;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_59_cse;
  wire [9:0] z_out_25;
  wire [10:0] nl_z_out_25;
  wire [9:0] z_out_27;
  wire [10:0] nl_z_out_27;
  wire [9:0] z_out_28;
  wire [10:0] nl_z_out_28;
  wire [9:0] z_out_30;
  wire [10:0] nl_z_out_30;
  wire [9:0] z_out_31;
  wire [10:0] nl_z_out_31;
  wire [9:0] z_out_32;
  wire [10:0] nl_z_out_32;
  wire [9:0] z_out_33;
  wire [10:0] nl_z_out_33;
  wire [21:0] z_out_194;
  wire [22:0] nl_z_out_194;
  wire [21:0] z_out_195;
  wire [22:0] nl_z_out_195;
  wire [21:0] z_out_196;
  wire [22:0] nl_z_out_196;
  wire [21:0] z_out_197;
  wire [22:0] nl_z_out_197;
  wire [21:0] z_out_198;
  wire [22:0] nl_z_out_198;
  wire [21:0] z_out_199;
  wire [22:0] nl_z_out_199;
  wire [21:0] z_out_200;
  wire [22:0] nl_z_out_200;
  wire [21:0] z_out_201;
  wire [22:0] nl_z_out_201;
  wire [21:0] z_out_202;
  wire [22:0] nl_z_out_202;
  wire [21:0] z_out_203;
  wire [22:0] nl_z_out_203;
  wire [21:0] z_out_204;
  wire [22:0] nl_z_out_204;
  wire [21:0] z_out_205;
  wire [22:0] nl_z_out_205;
  wire [21:0] z_out_206;
  wire [22:0] nl_z_out_206;
  wire [21:0] z_out_207;
  wire [22:0] nl_z_out_207;
  wire [21:0] z_out_208;
  wire [22:0] nl_z_out_208;
  wire [21:0] z_out_209;
  wire [22:0] nl_z_out_209;
  wire [21:0] z_out_210;
  wire [22:0] nl_z_out_210;
  wire [21:0] z_out_211;
  wire [22:0] nl_z_out_211;
  wire [21:0] z_out_212;
  wire [22:0] nl_z_out_212;
  wire [21:0] z_out_213;
  wire [22:0] nl_z_out_213;
  wire [21:0] z_out_214;
  wire [22:0] nl_z_out_214;
  wire [21:0] z_out_215;
  wire [22:0] nl_z_out_215;
  wire [21:0] z_out_216;
  wire [22:0] nl_z_out_216;
  wire [21:0] z_out_217;
  wire [22:0] nl_z_out_217;
  wire [21:0] z_out_218;
  wire [22:0] nl_z_out_218;
  wire [21:0] z_out_219;
  wire [22:0] nl_z_out_219;
  wire [21:0] z_out_220;
  wire [22:0] nl_z_out_220;
  wire [21:0] z_out_221;
  wire [22:0] nl_z_out_221;
  wire [21:0] z_out_222;
  wire [22:0] nl_z_out_222;
  wire [21:0] z_out_223;
  wire [22:0] nl_z_out_223;
  wire [21:0] z_out_224;
  wire [22:0] nl_z_out_224;
  wire [21:0] z_out_225;
  wire [22:0] nl_z_out_225;
  wire [21:0] z_out_226;
  wire [22:0] nl_z_out_226;
  wire [21:0] z_out_227;
  wire [22:0] nl_z_out_227;
  wire [21:0] z_out_228;
  wire [22:0] nl_z_out_228;
  wire [21:0] z_out_229;
  wire [22:0] nl_z_out_229;
  wire [21:0] z_out_230;
  wire [22:0] nl_z_out_230;
  wire [21:0] z_out_231;
  wire [22:0] nl_z_out_231;
  wire [21:0] z_out_232;
  wire [22:0] nl_z_out_232;
  wire [21:0] z_out_233;
  wire [22:0] nl_z_out_233;
  wire [21:0] z_out_234;
  wire [22:0] nl_z_out_234;
  wire [21:0] z_out_235;
  wire [22:0] nl_z_out_235;
  wire [21:0] z_out_236;
  wire [22:0] nl_z_out_236;
  wire [21:0] z_out_237;
  wire [22:0] nl_z_out_237;
  wire [21:0] z_out_238;
  wire [22:0] nl_z_out_238;
  wire [21:0] z_out_239;
  wire [22:0] nl_z_out_239;
  wire [21:0] z_out_240;
  wire [22:0] nl_z_out_240;
  wire [21:0] z_out_241;
  wire [22:0] nl_z_out_241;
  wire [21:0] z_out_242;
  wire [22:0] nl_z_out_242;
  wire [21:0] z_out_243;
  wire [22:0] nl_z_out_243;
  wire [21:0] z_out_244;
  wire [22:0] nl_z_out_244;
  wire [21:0] z_out_245;
  wire [22:0] nl_z_out_245;
  wire [21:0] z_out_246;
  wire [22:0] nl_z_out_246;
  wire [21:0] z_out_247;
  wire [22:0] nl_z_out_247;
  wire [21:0] z_out_248;
  wire [22:0] nl_z_out_248;
  wire [21:0] z_out_249;
  wire [22:0] nl_z_out_249;
  wire [21:0] z_out_250;
  wire [22:0] nl_z_out_250;
  wire [21:0] z_out_251;
  wire [22:0] nl_z_out_251;
  wire [21:0] z_out_252;
  wire [22:0] nl_z_out_252;
  wire [21:0] z_out_253;
  wire [22:0] nl_z_out_253;
  wire [21:0] z_out_254;
  wire [22:0] nl_z_out_254;
  wire [21:0] z_out_255;
  wire [22:0] nl_z_out_255;
  wire [21:0] z_out_256;
  wire [22:0] nl_z_out_256;
  wire [21:0] z_out_257;
  wire [22:0] nl_z_out_257;
  wire [21:0] z_out_258;
  wire [22:0] nl_z_out_258;
  wire [21:0] z_out_259;
  wire [22:0] nl_z_out_259;
  wire [21:0] z_out_260;
  wire [22:0] nl_z_out_260;
  wire [21:0] z_out_261;
  wire [22:0] nl_z_out_261;
  wire [21:0] z_out_262;
  wire [22:0] nl_z_out_262;
  wire [21:0] z_out_263;
  wire [22:0] nl_z_out_263;
  wire [21:0] z_out_264;
  wire [22:0] nl_z_out_264;
  wire [21:0] z_out_265;
  wire [22:0] nl_z_out_265;
  wire [21:0] z_out_266;
  wire [22:0] nl_z_out_266;
  wire [21:0] z_out_267;
  wire [22:0] nl_z_out_267;
  wire [21:0] z_out_268;
  wire [22:0] nl_z_out_268;
  wire [21:0] z_out_269;
  wire [22:0] nl_z_out_269;
  wire [21:0] z_out_270;
  wire [22:0] nl_z_out_270;
  wire [21:0] z_out_271;
  wire [22:0] nl_z_out_271;
  wire [21:0] z_out_272;
  wire [22:0] nl_z_out_272;
  wire [21:0] z_out_273;
  wire [22:0] nl_z_out_273;
  wire [21:0] z_out_274;
  wire [22:0] nl_z_out_274;
  wire [21:0] z_out_275;
  wire [22:0] nl_z_out_275;
  wire [21:0] z_out_276;
  wire [22:0] nl_z_out_276;
  wire [21:0] z_out_277;
  wire [22:0] nl_z_out_277;
  wire [21:0] z_out_278;
  wire [22:0] nl_z_out_278;
  wire [21:0] z_out_279;
  wire [22:0] nl_z_out_279;
  wire [21:0] z_out_280;
  wire [22:0] nl_z_out_280;
  wire [21:0] z_out_281;
  wire [22:0] nl_z_out_281;
  wire [21:0] z_out_282;
  wire [22:0] nl_z_out_282;
  wire [21:0] z_out_283;
  wire [22:0] nl_z_out_283;
  wire [21:0] z_out_284;
  wire [22:0] nl_z_out_284;
  wire [21:0] z_out_285;
  wire [22:0] nl_z_out_285;
  wire [21:0] z_out_286;
  wire [22:0] nl_z_out_286;
  wire [21:0] z_out_287;
  wire [22:0] nl_z_out_287;
  wire [21:0] z_out_288;
  wire [22:0] nl_z_out_288;
  wire [21:0] z_out_289;
  wire [22:0] nl_z_out_289;
  wire [21:0] z_out_290;
  wire [22:0] nl_z_out_290;
  wire [21:0] z_out_291;
  wire [22:0] nl_z_out_291;
  wire [21:0] z_out_292;
  wire [22:0] nl_z_out_292;
  wire [21:0] z_out_293;
  wire [22:0] nl_z_out_293;
  wire [21:0] z_out_294;
  wire [22:0] nl_z_out_294;
  wire [21:0] z_out_295;
  wire [22:0] nl_z_out_295;
  wire [21:0] z_out_296;
  wire [22:0] nl_z_out_296;
  wire [21:0] z_out_297;
  wire [22:0] nl_z_out_297;
  wire [21:0] z_out_298;
  wire [22:0] nl_z_out_298;
  wire [21:0] z_out_299;
  wire [22:0] nl_z_out_299;
  wire [21:0] z_out_300;
  wire [22:0] nl_z_out_300;
  wire [21:0] z_out_301;
  wire [22:0] nl_z_out_301;
  wire [21:0] z_out_302;
  wire [22:0] nl_z_out_302;
  wire [21:0] z_out_303;
  wire [22:0] nl_z_out_303;
  wire [21:0] z_out_304;
  wire [22:0] nl_z_out_304;
  wire [21:0] z_out_305;
  wire [22:0] nl_z_out_305;
  wire [21:0] z_out_306;
  wire [22:0] nl_z_out_306;
  wire [21:0] z_out_307;
  wire [22:0] nl_z_out_307;
  wire [21:0] z_out_308;
  wire [22:0] nl_z_out_308;
  wire [21:0] z_out_309;
  wire [22:0] nl_z_out_309;
  wire [21:0] z_out_310;
  wire [22:0] nl_z_out_310;
  wire [21:0] z_out_311;
  wire [22:0] nl_z_out_311;
  wire [21:0] z_out_312;
  wire [22:0] nl_z_out_312;
  wire [21:0] z_out_313;
  wire [22:0] nl_z_out_313;
  wire [21:0] z_out_314;
  wire [22:0] nl_z_out_314;
  wire [21:0] z_out_315;
  wire [22:0] nl_z_out_315;
  wire [21:0] z_out_316;
  wire [22:0] nl_z_out_316;
  wire [21:0] z_out_317;
  wire [22:0] nl_z_out_317;
  wire [21:0] z_out_318;
  wire [22:0] nl_z_out_318;
  wire [21:0] z_out_319;
  wire [22:0] nl_z_out_319;
  wire [21:0] z_out_320;
  wire [22:0] nl_z_out_320;
  wire [21:0] z_out_321;
  wire [22:0] nl_z_out_321;
  wire [21:0] z_out_322;
  wire [22:0] nl_z_out_322;
  wire [21:0] z_out_323;
  wire [22:0] nl_z_out_323;
  wire [21:0] z_out_324;
  wire [22:0] nl_z_out_324;
  wire [21:0] z_out_325;
  wire [22:0] nl_z_out_325;
  wire [21:0] z_out_326;
  wire [22:0] nl_z_out_326;
  wire [21:0] z_out_327;
  wire [22:0] nl_z_out_327;
  wire [21:0] z_out_328;
  wire [22:0] nl_z_out_328;
  wire [21:0] z_out_329;
  wire [22:0] nl_z_out_329;
  wire [21:0] z_out_330;
  wire [22:0] nl_z_out_330;
  wire [21:0] z_out_331;
  wire [22:0] nl_z_out_331;
  wire [21:0] z_out_332;
  wire [22:0] nl_z_out_332;
  wire [21:0] z_out_333;
  wire [22:0] nl_z_out_333;
  wire [21:0] z_out_334;
  wire [22:0] nl_z_out_334;
  wire [21:0] z_out_335;
  wire [22:0] nl_z_out_335;
  wire [21:0] z_out_336;
  wire [22:0] nl_z_out_336;
  wire [21:0] z_out_337;
  wire [22:0] nl_z_out_337;
  wire [21:0] z_out_338;
  wire [22:0] nl_z_out_338;
  wire [21:0] z_out_339;
  wire [22:0] nl_z_out_339;
  wire [21:0] z_out_340;
  wire [22:0] nl_z_out_340;
  wire [21:0] z_out_341;
  wire [22:0] nl_z_out_341;
  wire [21:0] z_out_342;
  wire [22:0] nl_z_out_342;
  wire [21:0] z_out_343;
  wire [22:0] nl_z_out_343;
  wire [21:0] z_out_344;
  wire [22:0] nl_z_out_344;
  wire [21:0] z_out_345;
  wire [22:0] nl_z_out_345;
  wire [21:0] z_out_346;
  wire [22:0] nl_z_out_346;
  wire [21:0] z_out_347;
  wire [22:0] nl_z_out_347;
  wire [21:0] z_out_348;
  wire [22:0] nl_z_out_348;
  wire [21:0] z_out_349;
  wire [22:0] nl_z_out_349;
  wire [21:0] z_out_350;
  wire [22:0] nl_z_out_350;
  wire [21:0] z_out_351;
  wire [22:0] nl_z_out_351;
  wire [21:0] z_out_352;
  wire [22:0] nl_z_out_352;
  wire [21:0] z_out_353;
  wire [22:0] nl_z_out_353;
  wire [21:0] z_out_354;
  wire [22:0] nl_z_out_354;
  wire [21:0] z_out_355;
  wire [22:0] nl_z_out_355;
  wire [21:0] z_out_356;
  wire [22:0] nl_z_out_356;
  wire [21:0] z_out_357;
  wire [22:0] nl_z_out_357;
  wire [21:0] z_out_358;
  wire [22:0] nl_z_out_358;
  wire [21:0] z_out_359;
  wire [22:0] nl_z_out_359;
  wire [21:0] z_out_360;
  wire [22:0] nl_z_out_360;
  wire [21:0] z_out_361;
  wire [22:0] nl_z_out_361;
  wire [21:0] z_out_362;
  wire [22:0] nl_z_out_362;
  wire [21:0] z_out_363;
  wire [22:0] nl_z_out_363;
  wire [21:0] z_out_364;
  wire [22:0] nl_z_out_364;
  wire [21:0] z_out_365;
  wire [22:0] nl_z_out_365;
  wire [21:0] z_out_366;
  wire [22:0] nl_z_out_366;
  wire [21:0] z_out_367;
  wire [22:0] nl_z_out_367;
  wire [21:0] z_out_368;
  wire [22:0] nl_z_out_368;
  wire [21:0] z_out_369;
  wire [22:0] nl_z_out_369;
  wire [21:0] z_out_370;
  wire [22:0] nl_z_out_370;
  wire [21:0] z_out_371;
  wire [22:0] nl_z_out_371;
  wire [21:0] z_out_372;
  wire [22:0] nl_z_out_372;
  wire [21:0] z_out_373;
  wire [22:0] nl_z_out_373;
  wire [21:0] z_out_374;
  wire [22:0] nl_z_out_374;
  wire [21:0] z_out_375;
  wire [22:0] nl_z_out_375;
  wire [21:0] z_out_376;
  wire [22:0] nl_z_out_376;
  wire [21:0] z_out_377;
  wire [22:0] nl_z_out_377;
  wire [21:0] z_out_378;
  wire [22:0] nl_z_out_378;
  wire [21:0] z_out_379;
  wire [22:0] nl_z_out_379;
  wire [21:0] z_out_380;
  wire [22:0] nl_z_out_380;
  wire [21:0] z_out_381;
  wire [22:0] nl_z_out_381;
  wire [21:0] z_out_382;
  wire [22:0] nl_z_out_382;
  wire [21:0] z_out_383;
  wire [22:0] nl_z_out_383;
  wire [21:0] z_out_384;
  wire [22:0] nl_z_out_384;
  wire [21:0] z_out_385;
  wire [22:0] nl_z_out_385;
  wire [21:0] z_out_386;
  wire [22:0] nl_z_out_386;
  wire [21:0] z_out_387;
  wire [22:0] nl_z_out_387;
  wire [21:0] z_out_388;
  wire [22:0] nl_z_out_388;
  wire [21:0] z_out_389;
  wire [22:0] nl_z_out_389;
  wire [21:0] z_out_390;
  wire [22:0] nl_z_out_390;
  wire [21:0] z_out_391;
  wire [22:0] nl_z_out_391;
  wire [21:0] z_out_392;
  wire [22:0] nl_z_out_392;
  wire [21:0] z_out_393;
  wire [22:0] nl_z_out_393;
  wire [21:0] z_out_394;
  wire [22:0] nl_z_out_394;
  wire [21:0] z_out_395;
  wire [22:0] nl_z_out_395;
  wire [21:0] z_out_396;
  wire [22:0] nl_z_out_396;
  wire [21:0] z_out_397;
  wire [22:0] nl_z_out_397;
  wire [21:0] z_out_398;
  wire [22:0] nl_z_out_398;
  wire [21:0] z_out_399;
  wire [22:0] nl_z_out_399;
  wire [21:0] z_out_400;
  wire [22:0] nl_z_out_400;
  wire [21:0] z_out_401;
  wire [22:0] nl_z_out_401;
  wire [21:0] z_out_402;
  wire [22:0] nl_z_out_402;
  wire [21:0] z_out_403;
  wire [22:0] nl_z_out_403;
  wire [21:0] z_out_404;
  wire [22:0] nl_z_out_404;
  wire [21:0] z_out_405;
  wire [22:0] nl_z_out_405;
  wire [21:0] z_out_406;
  wire [22:0] nl_z_out_406;
  wire [21:0] z_out_407;
  wire [22:0] nl_z_out_407;
  wire [21:0] z_out_408;
  wire [22:0] nl_z_out_408;
  wire [21:0] z_out_409;
  wire [22:0] nl_z_out_409;
  wire [21:0] z_out_410;
  wire [22:0] nl_z_out_410;
  wire [21:0] z_out_411;
  wire [22:0] nl_z_out_411;
  wire [21:0] z_out_412;
  wire [22:0] nl_z_out_412;
  wire [21:0] z_out_413;
  wire [22:0] nl_z_out_413;
  wire [21:0] z_out_414;
  wire [22:0] nl_z_out_414;
  wire [21:0] z_out_415;
  wire [22:0] nl_z_out_415;
  wire [21:0] z_out_416;
  wire [22:0] nl_z_out_416;
  wire [21:0] z_out_417;
  wire [22:0] nl_z_out_417;
  wire [21:0] z_out_418;
  wire [22:0] nl_z_out_418;
  wire [21:0] z_out_419;
  wire [22:0] nl_z_out_419;
  wire [21:0] z_out_420;
  wire [22:0] nl_z_out_420;
  wire [21:0] z_out_421;
  wire [22:0] nl_z_out_421;
  wire [21:0] z_out_422;
  wire [22:0] nl_z_out_422;
  wire [21:0] z_out_423;
  wire [22:0] nl_z_out_423;
  wire [21:0] z_out_424;
  wire [22:0] nl_z_out_424;
  wire [21:0] z_out_425;
  wire [22:0] nl_z_out_425;
  wire [21:0] z_out_426;
  wire [22:0] nl_z_out_426;
  wire [21:0] z_out_427;
  wire [22:0] nl_z_out_427;
  wire [21:0] z_out_428;
  wire [22:0] nl_z_out_428;
  wire [21:0] z_out_429;
  wire [22:0] nl_z_out_429;
  wire [21:0] z_out_430;
  wire [22:0] nl_z_out_430;
  wire [21:0] z_out_431;
  wire [22:0] nl_z_out_431;
  wire [21:0] z_out_432;
  wire [22:0] nl_z_out_432;
  wire [21:0] z_out_433;
  wire [22:0] nl_z_out_433;
  wire [21:0] z_out_434;
  wire [22:0] nl_z_out_434;
  wire [21:0] z_out_435;
  wire [22:0] nl_z_out_435;
  wire [21:0] z_out_436;
  wire [22:0] nl_z_out_436;
  wire [21:0] z_out_437;
  wire [22:0] nl_z_out_437;
  wire [21:0] z_out_438;
  wire [22:0] nl_z_out_438;
  wire [21:0] z_out_439;
  wire [22:0] nl_z_out_439;
  wire [21:0] z_out_440;
  wire [22:0] nl_z_out_440;
  wire [21:0] z_out_441;
  wire [22:0] nl_z_out_441;
  wire [21:0] z_out_442;
  wire [22:0] nl_z_out_442;
  wire [21:0] z_out_443;
  wire [22:0] nl_z_out_443;
  wire [21:0] z_out_444;
  wire [22:0] nl_z_out_444;
  wire [21:0] z_out_445;
  wire [22:0] nl_z_out_445;
  wire [21:0] z_out_446;
  wire [22:0] nl_z_out_446;
  wire [21:0] z_out_447;
  wire [22:0] nl_z_out_447;
  wire [21:0] z_out_448;
  wire [22:0] nl_z_out_448;
  wire [21:0] z_out_449;
  wire [22:0] nl_z_out_449;
  wire [21:0] z_out_450;
  wire [22:0] nl_z_out_450;
  wire [21:0] z_out_451;
  wire [22:0] nl_z_out_451;
  wire [21:0] z_out_452;
  wire [22:0] nl_z_out_452;
  wire [21:0] z_out_453;
  wire [22:0] nl_z_out_453;
  wire [21:0] z_out_454;
  wire [22:0] nl_z_out_454;
  wire [21:0] z_out_455;
  wire [22:0] nl_z_out_455;
  wire [21:0] z_out_456;
  wire [22:0] nl_z_out_456;
  wire [21:0] z_out_457;
  wire [22:0] nl_z_out_457;
  wire [21:0] z_out_458;
  wire [22:0] nl_z_out_458;
  wire [21:0] z_out_459;
  wire [22:0] nl_z_out_459;
  wire [21:0] z_out_460;
  wire [22:0] nl_z_out_460;
  wire [21:0] z_out_461;
  wire [22:0] nl_z_out_461;
  wire [21:0] z_out_462;
  wire [22:0] nl_z_out_462;
  wire [21:0] z_out_463;
  wire [22:0] nl_z_out_463;
  wire [21:0] z_out_464;
  wire [22:0] nl_z_out_464;
  wire [21:0] z_out_465;
  wire [22:0] nl_z_out_465;
  wire [21:0] z_out_466;
  wire [22:0] nl_z_out_466;
  wire [21:0] z_out_467;
  wire [22:0] nl_z_out_467;
  wire [21:0] z_out_468;
  wire [22:0] nl_z_out_468;
  wire [21:0] z_out_469;
  wire [22:0] nl_z_out_469;
  wire [21:0] z_out_470;
  wire [22:0] nl_z_out_470;
  wire [21:0] z_out_471;
  wire [22:0] nl_z_out_471;
  wire [21:0] z_out_472;
  wire [22:0] nl_z_out_472;
  wire [21:0] z_out_473;
  wire [22:0] nl_z_out_473;
  wire [21:0] z_out_474;
  wire [22:0] nl_z_out_474;
  wire [21:0] z_out_475;
  wire [22:0] nl_z_out_475;
  wire [21:0] z_out_476;
  wire [22:0] nl_z_out_476;
  wire [21:0] z_out_477;
  wire [22:0] nl_z_out_477;
  wire [21:0] z_out_478;
  wire [22:0] nl_z_out_478;
  wire [21:0] z_out_479;
  wire [22:0] nl_z_out_479;
  wire [21:0] z_out_480;
  wire [22:0] nl_z_out_480;
  wire [21:0] z_out_481;
  wire [22:0] nl_z_out_481;
  wire [21:0] z_out_482;
  wire [22:0] nl_z_out_482;
  wire [21:0] z_out_483;
  wire [22:0] nl_z_out_483;
  wire [21:0] z_out_484;
  wire [22:0] nl_z_out_484;
  wire [21:0] z_out_485;
  wire [22:0] nl_z_out_485;
  wire [21:0] z_out_486;
  wire [22:0] nl_z_out_486;
  wire [21:0] z_out_487;
  wire [22:0] nl_z_out_487;
  wire [21:0] z_out_488;
  wire [22:0] nl_z_out_488;
  wire [21:0] z_out_489;
  wire [22:0] nl_z_out_489;
  wire [21:0] z_out_490;
  wire [22:0] nl_z_out_490;
  wire [21:0] z_out_491;
  wire [22:0] nl_z_out_491;
  wire [21:0] z_out_492;
  wire [22:0] nl_z_out_492;
  wire [21:0] z_out_493;
  wire [22:0] nl_z_out_493;
  wire [21:0] z_out_494;
  wire [22:0] nl_z_out_494;
  wire [21:0] z_out_495;
  wire [22:0] nl_z_out_495;
  wire [21:0] z_out_496;
  wire [22:0] nl_z_out_496;
  wire [21:0] z_out_497;
  wire [22:0] nl_z_out_497;
  wire [21:0] z_out_498;
  wire [22:0] nl_z_out_498;
  wire [21:0] z_out_499;
  wire [22:0] nl_z_out_499;
  wire [21:0] z_out_500;
  wire [22:0] nl_z_out_500;
  wire [21:0] z_out_501;
  wire [22:0] nl_z_out_501;
  wire [21:0] z_out_502;
  wire [22:0] nl_z_out_502;
  wire [21:0] z_out_503;
  wire [22:0] nl_z_out_503;
  wire [21:0] z_out_504;
  wire [22:0] nl_z_out_504;
  wire [21:0] z_out_505;
  wire [22:0] nl_z_out_505;
  wire [21:0] z_out_506;
  wire [22:0] nl_z_out_506;
  wire [21:0] z_out_507;
  wire [22:0] nl_z_out_507;
  wire [21:0] z_out_508;
  wire [22:0] nl_z_out_508;
  wire [21:0] z_out_509;
  wire [22:0] nl_z_out_509;
  wire [21:0] z_out_510;
  wire [22:0] nl_z_out_510;
  wire [21:0] z_out_511;
  wire [22:0] nl_z_out_511;
  wire [21:0] z_out_512;
  wire [22:0] nl_z_out_512;
  wire [21:0] z_out_513;
  wire [22:0] nl_z_out_513;
  wire [21:0] z_out_514;
  wire [22:0] nl_z_out_514;
  wire [21:0] z_out_515;
  wire [22:0] nl_z_out_515;
  wire [21:0] z_out_516;
  wire [22:0] nl_z_out_516;
  wire [21:0] z_out_517;
  wire [22:0] nl_z_out_517;
  wire [21:0] z_out_518;
  wire [22:0] nl_z_out_518;
  wire [21:0] z_out_519;
  wire [22:0] nl_z_out_519;
  wire [21:0] z_out_520;
  wire [22:0] nl_z_out_520;
  wire [21:0] z_out_521;
  wire [22:0] nl_z_out_521;
  wire [21:0] z_out_522;
  wire [22:0] nl_z_out_522;
  wire [21:0] z_out_523;
  wire [22:0] nl_z_out_523;
  wire [21:0] z_out_524;
  wire [22:0] nl_z_out_524;
  wire [21:0] z_out_525;
  wire [22:0] nl_z_out_525;
  wire [21:0] z_out_526;
  wire [22:0] nl_z_out_526;
  wire [21:0] z_out_527;
  wire [22:0] nl_z_out_527;
  wire [21:0] z_out_528;
  wire [22:0] nl_z_out_528;
  wire [21:0] z_out_529;
  wire [22:0] nl_z_out_529;
  wire [21:0] z_out_530;
  wire [22:0] nl_z_out_530;
  wire [21:0] z_out_531;
  wire [22:0] nl_z_out_531;
  wire [21:0] z_out_532;
  wire [22:0] nl_z_out_532;
  wire [21:0] z_out_533;
  wire [22:0] nl_z_out_533;
  wire [21:0] z_out_534;
  wire [22:0] nl_z_out_534;
  wire [21:0] z_out_535;
  wire [22:0] nl_z_out_535;
  wire [21:0] z_out_536;
  wire [22:0] nl_z_out_536;
  wire [21:0] z_out_537;
  wire [22:0] nl_z_out_537;
  wire [21:0] z_out_538;
  wire [22:0] nl_z_out_538;
  wire [21:0] z_out_539;
  wire [22:0] nl_z_out_539;
  wire [21:0] z_out_540;
  wire [22:0] nl_z_out_540;
  wire [21:0] z_out_541;
  wire [22:0] nl_z_out_541;
  wire [21:0] z_out_542;
  wire [22:0] nl_z_out_542;
  wire [21:0] z_out_543;
  wire [22:0] nl_z_out_543;
  wire [21:0] z_out_544;
  wire [22:0] nl_z_out_544;
  wire [21:0] z_out_545;
  wire [22:0] nl_z_out_545;
  wire [21:0] z_out_546;
  wire [22:0] nl_z_out_546;
  wire [21:0] z_out_547;
  wire [22:0] nl_z_out_547;
  wire [21:0] z_out_548;
  wire [22:0] nl_z_out_548;
  wire [21:0] z_out_549;
  wire [22:0] nl_z_out_549;
  wire [21:0] z_out_550;
  wire [22:0] nl_z_out_550;
  wire [21:0] z_out_551;
  wire [22:0] nl_z_out_551;
  wire [21:0] z_out_552;
  wire [22:0] nl_z_out_552;
  wire [21:0] z_out_553;
  wire [22:0] nl_z_out_553;
  wire [21:0] z_out_554;
  wire [22:0] nl_z_out_554;
  wire [21:0] z_out_555;
  wire [22:0] nl_z_out_555;
  wire [21:0] z_out_556;
  wire [22:0] nl_z_out_556;
  wire [21:0] z_out_557;
  wire [22:0] nl_z_out_557;
  wire [21:0] z_out_558;
  wire [22:0] nl_z_out_558;
  wire [21:0] z_out_559;
  wire [22:0] nl_z_out_559;
  wire [21:0] z_out_560;
  wire [22:0] nl_z_out_560;
  wire [21:0] z_out_561;
  wire [22:0] nl_z_out_561;
  wire [21:0] z_out_562;
  wire [22:0] nl_z_out_562;
  wire [21:0] z_out_563;
  wire [22:0] nl_z_out_563;
  wire [21:0] z_out_564;
  wire [22:0] nl_z_out_564;
  wire [21:0] z_out_565;
  wire [22:0] nl_z_out_565;
  wire [21:0] z_out_566;
  wire [22:0] nl_z_out_566;
  wire [21:0] z_out_567;
  wire [22:0] nl_z_out_567;
  wire [21:0] z_out_680;
  wire [22:0] nl_z_out_680;
  wire [21:0] z_out_681;
  wire [22:0] nl_z_out_681;
  wire [21:0] z_out_682;
  wire [22:0] nl_z_out_682;
  wire [21:0] z_out_683;
  wire [22:0] nl_z_out_683;
  wire [21:0] z_out_684;
  wire [22:0] nl_z_out_684;
  wire [21:0] z_out_685;
  wire [22:0] nl_z_out_685;
  wire [21:0] z_out_686;
  wire [22:0] nl_z_out_686;
  wire [21:0] z_out_687;
  wire [22:0] nl_z_out_687;
  wire [21:0] z_out_688;
  wire [22:0] nl_z_out_688;
  wire [21:0] z_out_689;
  wire [22:0] nl_z_out_689;
  wire [21:0] z_out_690;
  wire [22:0] nl_z_out_690;
  wire [21:0] z_out_691;
  wire [22:0] nl_z_out_691;
  wire [21:0] z_out_692;
  wire [22:0] nl_z_out_692;
  wire [21:0] z_out_693;
  wire [22:0] nl_z_out_693;
  wire [21:0] z_out_694;
  wire [22:0] nl_z_out_694;
  wire [21:0] z_out_695;
  wire [22:0] nl_z_out_695;
  wire [21:0] z_out_696;
  wire [22:0] nl_z_out_696;
  wire [21:0] z_out_697;
  wire [22:0] nl_z_out_697;
  wire [21:0] z_out_698;
  wire [22:0] nl_z_out_698;
  wire [21:0] z_out_699;
  wire [22:0] nl_z_out_699;
  wire [21:0] z_out_700;
  wire [22:0] nl_z_out_700;
  wire [21:0] z_out_701;
  wire [22:0] nl_z_out_701;
  wire [21:0] z_out_702;
  wire [22:0] nl_z_out_702;
  wire [21:0] z_out_703;
  wire [22:0] nl_z_out_703;
  wire [21:0] z_out_704;
  wire [22:0] nl_z_out_704;
  wire [21:0] z_out_705;
  wire [22:0] nl_z_out_705;
  wire [21:0] z_out_706;
  wire [22:0] nl_z_out_706;
  wire [21:0] z_out_707;
  wire [22:0] nl_z_out_707;
  wire [21:0] z_out_708;
  wire [22:0] nl_z_out_708;
  wire [21:0] z_out_709;
  wire [22:0] nl_z_out_709;
  wire [21:0] z_out_710;
  wire [22:0] nl_z_out_710;
  wire [21:0] z_out_711;
  wire [22:0] nl_z_out_711;
  wire [21:0] z_out_712;
  wire [22:0] nl_z_out_712;
  wire [21:0] z_out_713;
  wire [22:0] nl_z_out_713;
  wire [21:0] z_out_714;
  wire [22:0] nl_z_out_714;
  wire [21:0] z_out_715;
  wire [22:0] nl_z_out_715;
  wire [21:0] z_out_716;
  wire [22:0] nl_z_out_716;
  wire [21:0] z_out_717;
  wire [22:0] nl_z_out_717;
  wire [21:0] z_out_718;
  wire [22:0] nl_z_out_718;
  wire [21:0] z_out_719;
  wire [22:0] nl_z_out_719;
  wire [21:0] z_out_720;
  wire [22:0] nl_z_out_720;
  wire [21:0] z_out_721;
  wire [22:0] nl_z_out_721;
  wire [21:0] z_out_722;
  wire [22:0] nl_z_out_722;
  wire [21:0] z_out_723;
  wire [22:0] nl_z_out_723;
  wire [21:0] z_out_724;
  wire [22:0] nl_z_out_724;
  wire [21:0] z_out_725;
  wire [22:0] nl_z_out_725;
  wire [21:0] z_out_726;
  wire [22:0] nl_z_out_726;
  wire [21:0] z_out_727;
  wire [22:0] nl_z_out_727;
  wire [21:0] z_out_728;
  wire [22:0] nl_z_out_728;
  wire [21:0] z_out_729;
  wire [22:0] nl_z_out_729;
  wire [21:0] z_out_730;
  wire [22:0] nl_z_out_730;
  wire [21:0] z_out_731;
  wire [22:0] nl_z_out_731;
  wire [21:0] z_out_732;
  wire [22:0] nl_z_out_732;
  wire [21:0] z_out_733;
  wire [22:0] nl_z_out_733;
  wire [21:0] z_out_734;
  wire [22:0] nl_z_out_734;
  wire [21:0] z_out_735;
  wire [22:0] nl_z_out_735;
  wire [21:0] z_out_736;
  wire [22:0] nl_z_out_736;
  wire [21:0] z_out_737;
  wire [22:0] nl_z_out_737;
  wire [21:0] z_out_738;
  wire [22:0] nl_z_out_738;
  wire [21:0] z_out_739;
  wire [22:0] nl_z_out_739;
  wire [21:0] z_out_740;
  wire [22:0] nl_z_out_740;
  wire [21:0] z_out_741;
  wire [22:0] nl_z_out_741;
  wire [21:0] z_out_742;
  wire [22:0] nl_z_out_742;
  wire [21:0] z_out_743;
  wire [22:0] nl_z_out_743;
  wire [21:0] z_out_744;
  wire [22:0] nl_z_out_744;
  wire [21:0] z_out_745;
  wire [22:0] nl_z_out_745;
  wire [21:0] z_out_746;
  wire [22:0] nl_z_out_746;
  wire [21:0] z_out_747;
  wire [22:0] nl_z_out_747;
  wire [21:0] z_out_748;
  wire [22:0] nl_z_out_748;
  wire [21:0] z_out_749;
  wire [22:0] nl_z_out_749;
  wire [21:0] z_out_750;
  wire [22:0] nl_z_out_750;
  wire [21:0] z_out_751;
  wire [22:0] nl_z_out_751;
  wire [21:0] z_out_752;
  wire [22:0] nl_z_out_752;
  wire [21:0] z_out_753;
  wire [22:0] nl_z_out_753;
  wire [21:0] z_out_754;
  wire [22:0] nl_z_out_754;
  wire [21:0] z_out_755;
  wire [22:0] nl_z_out_755;
  wire [21:0] z_out_756;
  wire [22:0] nl_z_out_756;
  wire [21:0] z_out_757;
  wire [22:0] nl_z_out_757;
  wire [21:0] z_out_758;
  wire [22:0] nl_z_out_758;
  wire [21:0] z_out_759;
  wire [22:0] nl_z_out_759;
  wire [21:0] z_out_760;
  wire [22:0] nl_z_out_760;
  wire [21:0] z_out_761;
  wire [22:0] nl_z_out_761;
  wire [21:0] z_out_762;
  wire [22:0] nl_z_out_762;
  wire [21:0] z_out_763;
  wire [22:0] nl_z_out_763;
  wire [21:0] z_out_764;
  wire [22:0] nl_z_out_764;
  wire [21:0] z_out_765;
  wire [22:0] nl_z_out_765;
  wire [21:0] z_out_766;
  wire [22:0] nl_z_out_766;
  wire [21:0] z_out_767;
  wire [22:0] nl_z_out_767;
  wire [21:0] z_out_768;
  wire [22:0] nl_z_out_768;
  wire [21:0] z_out_769;
  wire [22:0] nl_z_out_769;
  wire [21:0] z_out_770;
  wire [22:0] nl_z_out_770;
  wire [21:0] z_out_771;
  wire [22:0] nl_z_out_771;
  wire [21:0] z_out_772;
  wire [22:0] nl_z_out_772;
  wire [21:0] z_out_773;
  wire [22:0] nl_z_out_773;
  wire [21:0] z_out_774;
  wire [22:0] nl_z_out_774;
  wire [21:0] z_out_775;
  wire [22:0] nl_z_out_775;
  wire [21:0] z_out_776;
  wire [22:0] nl_z_out_776;
  wire [21:0] z_out_777;
  wire [22:0] nl_z_out_777;
  wire [21:0] z_out_778;
  wire [22:0] nl_z_out_778;
  wire or_tmp_4503;
  wire [21:0] z_out_779;
  wire [22:0] nl_z_out_779;
  wire [21:0] z_out_780;
  wire [22:0] nl_z_out_780;
  wire [21:0] z_out_781;
  wire [22:0] nl_z_out_781;
  wire [21:0] z_out_782;
  wire [22:0] nl_z_out_782;
  wire [21:0] z_out_783;
  wire [22:0] nl_z_out_783;
  wire [21:0] z_out_784;
  wire [22:0] nl_z_out_784;
  wire [21:0] z_out_785;
  wire [22:0] nl_z_out_785;
  wire [21:0] z_out_786;
  wire [22:0] nl_z_out_786;
  wire [21:0] z_out_787;
  wire [22:0] nl_z_out_787;
  wire [21:0] z_out_788;
  wire [22:0] nl_z_out_788;
  wire [21:0] z_out_789;
  wire [22:0] nl_z_out_789;
  wire [21:0] z_out_790;
  wire [22:0] nl_z_out_790;
  wire [21:0] z_out_791;
  wire [22:0] nl_z_out_791;
  wire [21:0] z_out_792;
  wire [22:0] nl_z_out_792;
  wire [21:0] z_out_793;
  wire [22:0] nl_z_out_793;
  wire [21:0] z_out_794;
  wire [22:0] nl_z_out_794;
  wire [21:0] z_out_795;
  wire [22:0] nl_z_out_795;
  wire [21:0] z_out_796;
  wire [22:0] nl_z_out_796;
  wire [21:0] z_out_797;
  wire [22:0] nl_z_out_797;
  wire [21:0] z_out_798;
  wire [22:0] nl_z_out_798;
  wire [21:0] z_out_799;
  wire [22:0] nl_z_out_799;
  wire [21:0] z_out_800;
  wire [22:0] nl_z_out_800;
  wire [21:0] z_out_801;
  wire [22:0] nl_z_out_801;
  wire [21:0] z_out_802;
  wire [22:0] nl_z_out_802;
  wire [21:0] z_out_803;
  wire [22:0] nl_z_out_803;
  wire [21:0] z_out_804;
  wire [22:0] nl_z_out_804;
  wire [21:0] z_out_805;
  wire [22:0] nl_z_out_805;
  wire [21:0] z_out_806;
  wire [22:0] nl_z_out_806;
  wire [21:0] z_out_807;
  wire [22:0] nl_z_out_807;
  wire [21:0] z_out_808;
  wire [22:0] nl_z_out_808;
  wire [21:0] z_out_809;
  wire [22:0] nl_z_out_809;
  wire [21:0] z_out_810;
  wire [22:0] nl_z_out_810;
  wire [21:0] z_out_811;
  wire [22:0] nl_z_out_811;
  wire [21:0] z_out_812;
  wire [22:0] nl_z_out_812;
  wire [21:0] z_out_813;
  wire [22:0] nl_z_out_813;
  wire [21:0] z_out_814;
  wire [22:0] nl_z_out_814;
  wire [21:0] z_out_815;
  wire [22:0] nl_z_out_815;
  wire [21:0] z_out_816;
  wire [22:0] nl_z_out_816;
  wire [21:0] z_out_817;
  wire [22:0] nl_z_out_817;
  wire [21:0] z_out_818;
  wire [22:0] nl_z_out_818;
  wire [21:0] z_out_819;
  wire [22:0] nl_z_out_819;
  wire [21:0] z_out_820;
  wire [22:0] nl_z_out_820;
  wire [21:0] z_out_821;
  wire [22:0] nl_z_out_821;
  wire [21:0] z_out_822;
  wire [22:0] nl_z_out_822;
  wire [21:0] z_out_823;
  wire [22:0] nl_z_out_823;
  wire [21:0] z_out_824;
  wire [22:0] nl_z_out_824;
  wire [21:0] z_out_825;
  wire [22:0] nl_z_out_825;
  wire [21:0] z_out_826;
  wire [22:0] nl_z_out_826;
  wire [21:0] z_out_827;
  wire [22:0] nl_z_out_827;
  wire [21:0] z_out_828;
  wire [22:0] nl_z_out_828;
  wire [21:0] z_out_829;
  wire [22:0] nl_z_out_829;
  wire [21:0] z_out_830;
  wire [22:0] nl_z_out_830;
  wire [21:0] z_out_831;
  wire [22:0] nl_z_out_831;
  wire [21:0] z_out_832;
  wire [22:0] nl_z_out_832;
  wire [21:0] z_out_833;
  wire [22:0] nl_z_out_833;
  wire [21:0] z_out_834;
  wire [22:0] nl_z_out_834;
  wire [21:0] z_out_835;
  wire [22:0] nl_z_out_835;
  wire [21:0] z_out_836;
  wire [22:0] nl_z_out_836;
  wire [21:0] z_out_837;
  wire [22:0] nl_z_out_837;
  wire [21:0] z_out_838;
  wire [22:0] nl_z_out_838;
  wire [21:0] z_out_839;
  wire [22:0] nl_z_out_839;
  wire [21:0] z_out_840;
  wire [22:0] nl_z_out_840;
  wire [21:0] z_out_841;
  wire [22:0] nl_z_out_841;
  wire [21:0] z_out_842;
  wire [22:0] nl_z_out_842;
  wire [21:0] z_out_843;
  wire [22:0] nl_z_out_843;
  wire [21:0] z_out_844;
  wire [22:0] nl_z_out_844;
  wire [21:0] z_out_845;
  wire [22:0] nl_z_out_845;
  wire [21:0] z_out_846;
  wire [22:0] nl_z_out_846;
  wire [21:0] z_out_847;
  wire [22:0] nl_z_out_847;
  wire [21:0] z_out_848;
  wire [22:0] nl_z_out_848;
  wire [21:0] z_out_849;
  wire [22:0] nl_z_out_849;
  wire [21:0] z_out_850;
  wire [22:0] nl_z_out_850;
  wire [21:0] z_out_851;
  wire [22:0] nl_z_out_851;
  wire [21:0] z_out_852;
  wire [22:0] nl_z_out_852;
  reg [1055:0] ConvFiltWidth_else_io_read_input_1_rsc_cse_sva;
  reg [1727:0] ConvFiltWidth_else_io_read_w2_rsc_cse_sva;
  reg [63:0] nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm;
  reg [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm;
  reg [79:0] InitAccum_io_read_b4_rsc_cse_sva;
  reg [10239:0] MultLoop_io_read_w4_rsc_cse_sva;
  reg [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [21:0] AccumDotWidth_acc_1133_itm;
  reg [21:0] AccumDotWidth_acc_1135_itm;
  reg [21:0] AccumDotWidth_acc_1164_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [21:0] AccumDotWidth_acc_1167_itm;
  reg [21:0] AccumDotWidth_acc_1169_itm;
  reg [21:0] AccumDotWidth_acc_1181_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [21:0] AccumDotWidth_acc_1184_itm;
  reg [21:0] AccumDotWidth_acc_1186_itm;
  reg [21:0] AccumDotWidth_acc_1198_itm;
  reg [21:0] AccumDotWidth_acc_1201_itm;
  reg [21:0] AccumDotWidth_acc_1203_itm;
  reg [21:0] AccumDotWidth_acc_1218_itm;
  reg [21:0] AccumDotWidth_acc_1220_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [21:0] AccumDotWidth_acc_1235_itm;
  reg [20:0] ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm;
  reg [21:0] AccumDotWidth_acc_1274_itm;
  reg [21:0] AccumDotWidth_acc_1300_itm;
  reg [21:0] AccumDotWidth_acc_1326_itm;
  reg [21:0] AccumDotWidth_acc_1352_itm;
  reg [21:0] AccumDotWidth_acc_1371_itm;
  reg [21:0] AccumDotWidth_acc_1392_itm;
  reg [21:0] AccumDotWidth_acc_1378_itm;
  reg [21:0] AccumDotWidth_acc_1397_itm;
  reg [21:0] AccumDotWidth_acc_1426_itm;
  reg [21:0] AccumDotWidth_acc_1837_itm;
  reg [21:0] AccumDotWidth_acc_1845_itm;
  reg [21:0] AccumDotWidth_acc_1877_itm;
  reg [21:0] AccumDotWidth_acc_1871_itm;
  reg [21:0] AccumDotWidth_acc_1916_itm;
  reg [21:0] AccumDotWidth_acc_1932_itm;
  reg [21:0] AccumDotWidth_acc_1937_itm;
  reg [21:0] AccumDotWidth_acc_1945_itm;
  reg [21:0] MultLoop_acc_105_itm;
  reg [21:0] MultLoop_acc_102_itm;
  reg [21:0] MultLoop_acc_54_itm;
  reg [21:0] MultLoop_acc_128_itm;
  reg [21:0] MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_89_itm;
  reg [21:0] MultLoop_acc_88_itm;
  reg [21:0] MultLoop_acc_36_itm;
  reg [21:0] MultLoop_acc_113_itm;
  reg [21:0] MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_79_itm;
  reg [21:0] MultLoop_acc_123_itm;
  reg [21:0] MultLoop_acc_229_itm;
  reg [21:0] MultLoop_acc_181_itm;
  reg [21:0] MultLoop_acc_243_itm;
  reg [21:0] MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_215_itm;
  reg [21:0] MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_206_itm;
  reg [21:0] MultLoop_acc_250_itm;
  reg [21:0] MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_356_itm;
  reg [21:0] MultLoop_acc_372_itm;
  reg [21:0] MultLoop_acc_308_itm;
  reg [21:0] MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_333_itm;
  reg [21:0] MultLoop_acc_377_itm;
  reg [21:0] MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_502_itm;
  reg [21:0] MultLoop_acc_483_itm;
  reg [21:0] MultLoop_acc_499_itm;
  reg [21:0] MultLoop_acc_435_itm;
  reg [21:0] MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_470_itm;
  reg [21:0] MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_460_itm;
  reg [21:0] MultLoop_acc_504_itm;
  reg [21:0] MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_613_itm;
  reg [21:0] MultLoop_acc_629_itm;
  reg [21:0] MultLoop_acc_628_itm;
  reg [21:0] MultLoop_acc_626_itm;
  reg [21:0] MultLoop_acc_562_itm;
  reg [21:0] MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_597_itm;
  reg [21:0] MultLoop_acc_596_itm;
  reg [21:0] MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_587_itm;
  reg [21:0] MultLoop_acc_631_itm;
  reg [21:0] MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_740_itm;
  reg [21:0] MultLoop_acc_756_itm;
  reg [21:0] MultLoop_acc_689_itm;
  reg [21:0] MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_724_itm;
  wire [22:0] nl_MultLoop_acc_724_itm;
  reg [21:0] MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_714_itm;
  reg [21:0] MultLoop_acc_758_itm;
  reg [21:0] MultLoop_acc_867_itm;
  reg [21:0] MultLoop_acc_883_itm;
  wire [22:0] nl_MultLoop_acc_883_itm;
  reg [21:0] MultLoop_acc_861_itm;
  reg [21:0] MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_841_itm;
  reg [21:0] MultLoop_acc_885_itm;
  reg [21:0] MultLoop_acc_994_itm;
  reg [21:0] MultLoop_acc_1010_itm;
  reg [21:0] MultLoop_acc_1018_itm;
  reg [21:0] MultLoop_acc_1007_itm;
  reg [21:0] MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_1000_itm;
  reg [21:0] MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_968_itm;
  reg [21:0] MultLoop_acc_1012_itm;
  reg [21:0] MultLoop_acc_1089_itm;
  reg [21:0] MultLoop_acc_1121_itm;
  reg [21:0] MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_1095_itm;
  reg [21:0] MultLoop_acc_1139_itm;
  reg [21:0] MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  reg [21:0] MultLoop_acc_1222_itm;
  reg [21:0] MultLoop_acc_1266_itm;
  reg [10:0] MultLoop_acc_1280_psp;
  wire [11:0] nl_MultLoop_acc_1280_psp;
  reg [10:0] MultLoop_acc_1281_psp;
  wire [11:0] nl_MultLoop_acc_1281_psp;
  reg [10:0] MultLoop_acc_1282_psp;
  wire [11:0] nl_MultLoop_acc_1282_psp;
  reg [10:0] MultLoop_acc_1283_psp;
  wire [11:0] nl_MultLoop_acc_1283_psp;
  reg [10:0] MultLoop_acc_1284_psp;
  wire [11:0] nl_MultLoop_acc_1284_psp;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1;
  wire [21:0] MultLoop_acc_162_sdt;
  wire [22:0] nl_MultLoop_acc_162_sdt;
  wire [21:0] MultLoop_acc_27_sdt;
  wire [22:0] nl_MultLoop_acc_27_sdt;
  wire [21:0] MultLoop_acc_1193_sdt;
  wire [22:0] nl_MultLoop_acc_1193_sdt;
  wire [21:0] MultLoop_acc_1201_sdt;
  wire [22:0] nl_MultLoop_acc_1201_sdt;
  wire nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse;
  wire [20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse;
  wire [21:0] MultLoop_acc_1188_sdt;
  wire [22:0] nl_MultLoop_acc_1188_sdt;
  wire [21:0] MultLoop_acc_1185_sdt;
  wire [22:0] nl_MultLoop_acc_1185_sdt;
  wire [21:0] MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7;
  wire AccumDotWidth_or_38_cse;
  wire MultLoop_or_46_cse;
  wire z_out_22;
  wire z_out_1_22;
  wire z_out_2_22;
  wire z_out_3_22;
  wire z_out_4_22;
  wire z_out_5_22;
  wire z_out_6_22;
  wire z_out_7_22;
  wire z_out_8_22;
  wire z_out_9_22;
  wire z_out_10_22;
  wire z_out_11_22;
  wire z_out_12_22;
  wire z_out_13_22;
  wire z_out_14_22;
  wire z_out_15_22;
  wire z_out_16_22;
  wire z_out_17_22;
  wire z_out_18_22;
  wire z_out_19_22;
  wire z_out_20_22;
  wire z_out_21_22;
  wire z_out_22_22;
  wire z_out_23_22;
  wire z_out_24_22;
  wire [21:0] z_out_34_28_7;
  wire [21:0] z_out_35_28_7;
  wire [21:0] z_out_36_28_7;
  wire [21:0] z_out_37_28_7;
  wire [21:0] z_out_38_28_7;
  wire [21:0] z_out_39_28_7;
  wire [21:0] z_out_40_28_7;
  wire [21:0] z_out_41_28_7;
  wire [21:0] z_out_42_28_7;
  wire [21:0] z_out_43_28_7;
  wire [21:0] z_out_44_28_7;
  wire [21:0] z_out_45_28_7;
  wire [21:0] z_out_46_28_7;
  wire [21:0] z_out_47_28_7;
  wire [21:0] z_out_48_28_7;
  wire [21:0] z_out_49_28_7;
  wire [21:0] z_out_50_28_7;
  wire [21:0] z_out_51_28_7;
  wire [21:0] z_out_52_28_7;
  wire [21:0] z_out_53_28_7;
  wire [21:0] z_out_54_28_7;
  wire [21:0] z_out_55_28_7;
  wire [21:0] z_out_56_28_7;
  wire [21:0] z_out_57_28_7;
  wire [21:0] z_out_58_28_7;
  wire [21:0] z_out_59_28_7;
  wire [21:0] z_out_60_28_7;
  wire [21:0] z_out_61_28_7;
  wire [21:0] z_out_62_28_7;
  wire [21:0] z_out_63_28_7;
  wire [21:0] z_out_64_28_7;
  wire [21:0] z_out_65_28_7;
  wire [21:0] z_out_66_28_7;
  wire [21:0] z_out_67_28_7;
  wire [21:0] z_out_68_28_7;
  wire [21:0] z_out_69_28_7;
  wire [21:0] z_out_70_28_7;
  wire [21:0] z_out_71_28_7;
  wire [21:0] z_out_72_28_7;
  wire [21:0] z_out_73_28_7;
  wire [21:0] z_out_74_28_7;
  wire [21:0] z_out_75_28_7;
  wire [21:0] z_out_76_28_7;
  wire [21:0] z_out_77_28_7;
  wire [21:0] z_out_78_28_7;
  wire [21:0] z_out_79_28_7;
  wire [21:0] z_out_80_28_7;
  wire [21:0] z_out_81_28_7;
  wire [21:0] z_out_82_28_7;
  wire [21:0] z_out_83_28_7;
  wire [21:0] z_out_84_28_7;
  wire [21:0] z_out_85_28_7;
  wire [21:0] z_out_86_28_7;
  wire [21:0] z_out_87_28_7;
  wire [21:0] z_out_88_28_7;
  wire [21:0] z_out_89_28_7;
  wire [21:0] z_out_90_28_7;
  wire [21:0] z_out_91_28_7;
  wire [21:0] z_out_92_28_7;
  wire [21:0] z_out_93_28_7;
  wire [21:0] z_out_94_28_7;
  wire [21:0] z_out_95_28_7;
  wire [21:0] z_out_96_28_7;
  wire [21:0] z_out_97_28_7;
  wire [21:0] z_out_98_28_7;
  wire [21:0] z_out_99_28_7;
  wire [21:0] z_out_100_28_7;
  wire [21:0] z_out_101_28_7;
  wire [21:0] z_out_102_28_7;
  wire [21:0] z_out_103_28_7;
  wire [21:0] z_out_104_28_7;
  wire [21:0] z_out_105_28_7;
  wire [21:0] z_out_106_28_7;
  wire [21:0] z_out_107_28_7;
  wire [21:0] z_out_108_28_7;
  wire [21:0] z_out_109_28_7;
  wire [21:0] z_out_110_28_7;
  wire [21:0] z_out_111_28_7;
  wire [21:0] z_out_112_28_7;
  wire [21:0] z_out_113_28_7;
  wire [21:0] z_out_114_28_7;
  wire [21:0] z_out_115_28_7;
  wire [21:0] z_out_116_28_7;
  wire [21:0] z_out_117_28_7;
  wire [21:0] z_out_118_28_7;
  wire [21:0] z_out_119_28_7;
  wire [21:0] z_out_120_28_7;
  wire [21:0] z_out_121_28_7;
  wire [21:0] z_out_122_28_7;
  wire [21:0] z_out_123_28_7;
  wire [21:0] z_out_124_28_7;
  wire [21:0] z_out_125_28_7;
  wire [21:0] z_out_126_28_7;
  wire [21:0] z_out_127_28_7;
  wire [21:0] z_out_128_28_7;
  wire [21:0] z_out_129_28_7;
  wire [21:0] z_out_130_28_7;
  wire [21:0] z_out_131_28_7;
  wire [21:0] z_out_132_28_7;
  wire [21:0] z_out_133_28_7;
  wire [21:0] z_out_134_28_7;
  wire [21:0] z_out_135_28_7;
  wire [21:0] z_out_136_28_7;
  wire [21:0] z_out_137_28_7;
  wire [21:0] z_out_138_28_7;
  wire [21:0] z_out_139_28_7;
  wire [21:0] z_out_140_28_7;
  wire [21:0] z_out_141_28_7;
  wire [21:0] z_out_142_28_7;
  wire [21:0] z_out_143_28_7;
  wire [21:0] z_out_144_28_7;
  wire [21:0] z_out_145_28_7;
  wire [21:0] z_out_146_28_7;
  wire [21:0] z_out_147_28_7;
  wire [21:0] z_out_148_28_7;
  wire [21:0] z_out_149_28_7;
  wire [21:0] z_out_150_28_7;
  wire [21:0] z_out_151_28_7;
  wire [21:0] z_out_152_28_7;
  wire [21:0] z_out_153_28_7;
  wire [21:0] z_out_154_28_7;
  wire [21:0] z_out_155_28_7;
  wire [21:0] z_out_156_28_7;
  wire [21:0] z_out_157_28_7;
  wire [21:0] z_out_158_28_7;
  wire [21:0] z_out_159_28_7;
  wire [21:0] z_out_160_28_7;
  wire [21:0] z_out_161_28_7;
  wire [21:0] z_out_162_28_7;
  wire [21:0] z_out_163_28_7;
  wire [21:0] z_out_164_28_7;
  wire [21:0] z_out_165_28_7;
  wire [21:0] z_out_166_28_7;
  wire [21:0] z_out_167_28_7;
  wire [21:0] z_out_168_28_7;
  wire [21:0] z_out_169_28_7;
  wire [21:0] z_out_170_28_7;
  wire [21:0] z_out_171_28_7;
  wire [21:0] z_out_172_28_7;
  wire [21:0] z_out_173_28_7;
  wire [21:0] z_out_174_28_7;
  wire [21:0] z_out_175_28_7;
  wire [21:0] z_out_176_28_7;
  wire [21:0] z_out_177_28_7;
  wire [21:0] z_out_178_28_7;
  wire [21:0] z_out_179_28_7;
  wire [21:0] z_out_180_28_7;
  wire [21:0] z_out_181_28_7;
  wire [21:0] z_out_182_28_7;
  wire [21:0] z_out_183_28_7;
  wire [21:0] z_out_184_28_7;
  wire [21:0] z_out_185_28_7;
  wire [21:0] z_out_186_28_7;
  wire [21:0] z_out_187_28_7;
  wire [21:0] z_out_188_28_7;
  wire [21:0] z_out_189_28_7;
  wire [21:0] z_out_190_28_7;
  wire [21:0] z_out_191_28_7;
  wire [21:0] z_out_192_28_7;
  wire [21:0] z_out_193_28_7;
  wire [22:0] z_out_568_29_7;
  wire [22:0] z_out_569_29_7;
  wire [22:0] z_out_570_29_7;
  wire [22:0] z_out_571_29_7;
  wire [22:0] z_out_572_29_7;
  wire [22:0] z_out_573_29_7;
  wire [22:0] z_out_574_29_7;
  wire [22:0] z_out_575_29_7;
  wire [22:0] z_out_576_29_7;
  wire [22:0] z_out_577_29_7;
  wire [22:0] z_out_578_29_7;
  wire [22:0] z_out_579_29_7;
  wire [22:0] z_out_580_29_7;
  wire [22:0] z_out_581_29_7;
  wire [22:0] z_out_582_29_7;
  wire [22:0] z_out_583_29_7;
  wire [22:0] z_out_584_29_7;
  wire [22:0] z_out_585_29_7;
  wire [22:0] z_out_586_29_7;
  wire [22:0] z_out_587_29_7;
  wire [22:0] z_out_588_29_7;
  wire [22:0] z_out_589_29_7;
  wire [22:0] z_out_590_29_7;
  wire [22:0] z_out_591_29_7;
  wire [22:0] z_out_592_29_7;
  wire [22:0] z_out_593_29_7;
  wire [22:0] z_out_594_29_7;
  wire [22:0] z_out_595_29_7;
  wire [22:0] z_out_596_29_7;
  wire [22:0] z_out_597_29_7;
  wire [22:0] z_out_598_29_7;
  wire [22:0] z_out_599_29_7;
  wire [22:0] z_out_600_29_7;
  wire [22:0] z_out_601_29_7;
  wire [22:0] z_out_602_29_7;
  wire [22:0] z_out_603_29_7;
  wire [22:0] z_out_604_29_7;
  wire [22:0] z_out_605_29_7;
  wire [22:0] z_out_606_29_7;
  wire [22:0] z_out_607_29_7;
  wire [22:0] z_out_608_29_7;
  wire [22:0] z_out_609_29_7;
  wire [22:0] z_out_610_29_7;
  wire [22:0] z_out_611_29_7;
  wire [22:0] z_out_612_29_7;
  wire [22:0] z_out_613_29_7;
  wire [22:0] z_out_614_29_7;
  wire [22:0] z_out_615_29_7;
  wire [22:0] z_out_616_29_7;
  wire [22:0] z_out_617_29_7;
  wire [22:0] z_out_618_29_7;
  wire [22:0] z_out_619_29_7;
  wire [22:0] z_out_620_29_7;
  wire [22:0] z_out_621_29_7;
  wire [22:0] z_out_622_29_7;
  wire [22:0] z_out_623_29_7;
  wire [22:0] z_out_624_29_7;
  wire [22:0] z_out_625_29_7;
  wire [22:0] z_out_626_29_7;
  wire [22:0] z_out_627_29_7;
  wire [22:0] z_out_628_29_7;
  wire [22:0] z_out_629_29_7;
  wire [22:0] z_out_630_29_7;
  wire [21:0] z_out_631_28_7;
  wire [21:0] z_out_632_28_7;
  wire [21:0] z_out_633_28_7;
  wire [21:0] z_out_634_28_7;
  wire [21:0] z_out_635_28_7;
  wire [21:0] z_out_636_28_7;
  wire [21:0] z_out_637_28_7;
  wire [21:0] z_out_638_28_7;
  wire [21:0] z_out_639_28_7;
  wire [21:0] z_out_640_28_7;
  wire [21:0] z_out_641_28_7;
  wire [21:0] z_out_642_28_7;
  wire [21:0] z_out_643_28_7;
  wire [21:0] z_out_644_28_7;
  wire [21:0] z_out_645_28_7;
  wire [21:0] z_out_646_28_7;
  wire [21:0] z_out_647_28_7;
  wire [21:0] z_out_648_28_7;
  wire [21:0] z_out_649_28_7;
  wire [21:0] z_out_650_28_7;
  wire [21:0] z_out_651_28_7;
  wire [21:0] z_out_652_28_7;
  wire [21:0] z_out_653_28_7;
  wire [21:0] z_out_654_28_7;
  wire [21:0] z_out_655_28_7;
  wire [21:0] z_out_656_28_7;
  wire [21:0] z_out_657_28_7;
  wire [21:0] z_out_658_28_7;
  wire [21:0] z_out_659_28_7;
  wire [21:0] z_out_660_28_7;
  wire [21:0] z_out_661_28_7;
  wire [21:0] z_out_662_28_7;
  wire [21:0] z_out_663_28_7;
  wire [21:0] z_out_664_28_7;
  wire [21:0] z_out_665_28_7;
  wire [21:0] z_out_666_28_7;
  wire [21:0] z_out_667_28_7;
  wire [21:0] z_out_668_28_7;
  wire [21:0] z_out_669_28_7;
  wire [21:0] z_out_670_28_7;
  wire [21:0] z_out_671_28_7;
  wire [21:0] z_out_672_28_7;
  wire [21:0] z_out_673_28_7;
  wire [21:0] z_out_674_28_7;
  wire [21:0] z_out_675_28_7;
  wire [21:0] z_out_676_28_7;
  wire [21:0] z_out_677_28_7;
  wire [21:0] z_out_678_28_7;
  wire [21:0] z_out_679_28_7;
  wire [22:0] z_out_853_29_7;
  wire [22:0] z_out_854_29_7;
  wire [22:0] z_out_855_29_7;
  wire [22:0] z_out_856_29_7;
  wire [22:0] z_out_857_29_7;
  wire [22:0] z_out_858_29_7;
  wire [22:0] z_out_859_29_7;
  wire [22:0] z_out_860_29_7;
  wire [22:0] z_out_861_29_7;
  wire [22:0] z_out_862_29_7;
  wire [22:0] z_out_863_29_7;
  wire [22:0] z_out_864_29_7;
  wire [22:0] z_out_865_29_7;
  wire [22:0] z_out_866_29_7;
  wire [22:0] z_out_867_29_7;
  wire [22:0] z_out_868_29_7;
  wire [22:0] z_out_869_29_7;
  wire [22:0] z_out_870_29_7;
  wire [22:0] z_out_871_29_7;
  wire [22:0] z_out_872_29_7;
  wire [22:0] z_out_873_29_7;
  wire [22:0] z_out_874_29_7;
  wire [22:0] z_out_875_29_7;
  wire [22:0] z_out_876_29_7;
  wire [22:0] z_out_877_29_7;
  wire [22:0] z_out_878_29_7;
  wire [22:0] z_out_879_29_7;
  wire [22:0] z_out_880_29_7;
  wire [22:0] z_out_881_29_7;
  wire [22:0] z_out_882_29_7;
  wire [22:0] z_out_883_29_7;
  wire [22:0] z_out_884_29_7;
  wire [22:0] z_out_885_29_7;
  wire [22:0] z_out_886_29_7;
  wire [22:0] z_out_887_29_7;
  wire [22:0] z_out_888_29_7;
  wire [22:0] z_out_889_29_7;
  wire [22:0] z_out_890_29_7;
  wire [22:0] z_out_891_29_7;
  wire [22:0] z_out_892_29_7;
  wire [22:0] z_out_893_29_7;
  wire [22:0] z_out_894_29_7;
  wire [22:0] z_out_895_29_7;
  wire [22:0] z_out_896_29_7;
  wire [22:0] z_out_897_29_7;
  wire [22:0] z_out_898_29_7;
  wire [22:0] z_out_899_29_7;
  wire [22:0] z_out_900_29_7;
  wire [22:0] z_out_901_29_7;
  wire [22:0] z_out_902_29_7;
  wire [22:0] z_out_903_29_7;
  wire [20:0] z_out_904_29_9;
  wire [22:0] z_out_905_29_7;
  wire [22:0] z_out_906_29_7;
  wire [22:0] z_out_907_29_7;
  wire [22:0] z_out_908_29_7;
  wire [22:0] z_out_909_29_7;
  wire [22:0] z_out_910_29_7;
  wire [22:0] z_out_911_29_7;
  wire [22:0] z_out_912_29_7;
  wire [22:0] z_out_913_29_7;
  wire [22:0] z_out_914_29_7;
  wire [22:0] z_out_915_29_7;
  wire [22:0] z_out_916_29_7;
  wire [22:0] z_out_917_29_7;
  wire [22:0] z_out_918_29_7;
  wire [22:0] z_out_919_29_7;
  wire [22:0] z_out_920_29_7;
  wire [22:0] z_out_921_29_7;
  wire [22:0] z_out_922_29_7;
  wire [22:0] z_out_923_29_7;
  wire [22:0] z_out_924_29_7;
  wire [22:0] z_out_925_29_7;
  wire [22:0] z_out_926_29_7;
  wire [22:0] z_out_927_29_7;
  wire [22:0] z_out_928_29_7;
  wire [22:0] z_out_929_29_7;
  wire [22:0] z_out_930_29_7;
  wire [22:0] z_out_931_29_7;
  wire [22:0] z_out_932_29_7;
  wire [22:0] z_out_933_29_7;
  wire [22:0] z_out_934_29_7;
  wire [22:0] z_out_935_29_7;
  wire [22:0] z_out_936_29_7;
  wire [22:0] z_out_937_29_7;
  wire [22:0] z_out_938_29_7;
  wire [22:0] z_out_939_29_7;
  wire [22:0] z_out_940_29_7;
  wire [22:0] z_out_941_29_7;
  wire [20:0] z_out_942_29_9;
  wire [22:0] z_out_943_29_7;
  wire [22:0] z_out_944_29_7;
  wire [22:0] z_out_945_29_7;
  wire [22:0] z_out_946_29_7;
  wire [22:0] z_out_947_29_7;
  wire [22:0] z_out_948_29_7;
  wire [22:0] z_out_949_29_7;
  wire [22:0] z_out_950_29_7;
  wire [22:0] z_out_951_29_7;
  wire [22:0] z_out_952_29_7;
  wire [22:0] z_out_953_29_7;
  wire [22:0] z_out_954_29_7;
  wire [22:0] z_out_955_29_7;
  wire [22:0] z_out_956_29_7;
  wire [22:0] z_out_957_29_7;
  wire [22:0] z_out_958_29_7;
  wire [22:0] z_out_959_29_7;
  wire [22:0] z_out_960_29_7;
  wire [22:0] z_out_961_29_7;
  wire [20:0] z_out_962_29_9;
  wire [20:0] z_out_963_29_9;
  wire [22:0] z_out_964_29_7;
  wire [20:0] z_out_965_29_9;
  wire [22:0] z_out_966_29_7;
  wire [22:0] z_out_967_29_7;
  wire [22:0] z_out_968_29_7;
  wire [22:0] z_out_969_29_7;
  wire [22:0] z_out_970_29_7;
  wire [22:0] z_out_971_29_7;
  wire [22:0] z_out_972_29_7;
  wire [22:0] z_out_973_29_7;
  wire [22:0] z_out_974_29_7;
  wire [22:0] z_out_975_29_7;
  wire [22:0] z_out_976_29_7;
  wire [22:0] z_out_977_29_7;
  wire [20:0] z_out_978_29_9;
  wire [20:0] z_out_979_29_9;
  wire [22:0] z_out_980_29_7;
  wire [22:0] z_out_981_29_7;
  wire [22:0] z_out_982_29_7;
  wire [22:0] z_out_983_29_7;
  wire [22:0] z_out_984_29_7;
  wire [22:0] z_out_985_29_7;
  wire [22:0] z_out_986_29_7;
  wire [22:0] z_out_987_29_7;
  wire [20:0] z_out_988_29_9;
  wire [20:0] z_out_989_29_9;
  wire [22:0] z_out_990_29_7;
  wire [22:0] z_out_991_29_7;
  wire [20:0] z_out_992_29_9;
  wire [20:0] z_out_993_29_9;
  wire [22:0] z_out_994_29_7;
  wire [22:0] z_out_995_29_7;
  wire [22:0] z_out_996_29_7;
  wire [22:0] z_out_997_29_7;
  wire [22:0] z_out_998_29_7;
  wire [22:0] z_out_999_29_7;
  wire [22:0] z_out_1000_29_7;
  wire [22:0] z_out_1001_29_7;
  wire [22:0] z_out_1002_29_7;
  wire [20:0] z_out_1003_29_9;
  wire [20:0] z_out_1004_29_9;
  wire [22:0] z_out_1005_29_7;
  wire [20:0] z_out_1006_29_9;
  wire [22:0] z_out_1007_29_7;
  wire [22:0] z_out_1008_29_7;
  wire [22:0] z_out_1009_29_7;
  wire [22:0] z_out_1010_29_7;
  wire [22:0] z_out_1011_29_7;
  wire [22:0] z_out_1012_29_7;
  wire [22:0] z_out_1013_29_7;
  wire [22:0] z_out_1014_29_7;
  wire [22:0] z_out_1015_29_7;
  wire [22:0] z_out_1016_29_7;
  wire [20:0] z_out_1017_29_9;
  wire [20:0] z_out_1018_29_9;
  wire [22:0] z_out_1019_29_7;
  wire [20:0] z_out_1020_29_9;
  wire [22:0] z_out_1021_29_7;
  wire [22:0] z_out_1022_29_7;
  wire [22:0] z_out_1023_29_7;
  wire [22:0] z_out_1024_29_7;
  wire [22:0] z_out_1025_29_7;
  wire [22:0] z_out_1026_29_7;
  wire [22:0] z_out_1027_29_7;
  wire [22:0] z_out_1028_29_7;
  wire [22:0] z_out_1029_29_7;
  wire [22:0] z_out_1030_29_7;
  wire [20:0] z_out_1031_29_9;
  wire [20:0] z_out_1032_29_9;
  wire [20:0] z_out_1033_29_9;
  wire [22:0] z_out_1034_29_7;
  wire [22:0] z_out_1035_29_7;
  wire [22:0] z_out_1036_29_7;
  wire [22:0] z_out_1037_29_7;
  wire [22:0] z_out_1038_29_7;
  wire [22:0] z_out_1039_29_7;
  wire [22:0] z_out_1040_29_7;
  wire [22:0] z_out_1041_29_7;
  wire [22:0] z_out_1042_29_7;
  wire [22:0] z_out_1043_29_7;
  wire [22:0] z_out_1044_29_7;
  wire [22:0] z_out_1045_29_7;
  wire [20:0] z_out_1046_29_9;
  wire [20:0] z_out_1047_29_9;
  wire [20:0] z_out_1048_29_9;
  wire [22:0] z_out_1049_29_7;
  wire [22:0] z_out_1050_29_7;
  wire [22:0] z_out_1051_29_7;
  wire [22:0] z_out_1052_29_7;
  wire [22:0] z_out_1053_29_7;
  wire [22:0] z_out_1054_29_7;
  wire [22:0] z_out_1055_29_7;
  wire [22:0] z_out_1056_29_7;
  wire [22:0] z_out_1057_29_7;
  wire [22:0] z_out_1058_29_7;
  wire [20:0] z_out_1059_29_9;
  wire [20:0] z_out_1060_29_9;
  wire [20:0] z_out_1061_29_9;
  wire [20:0] z_out_1062_29_9;
  wire [20:0] z_out_1063_29_9;
  wire [22:0] z_out_1064_29_7;
  wire [20:0] z_out_1065_29_9;
  wire [20:0] z_out_1066_29_9;
  wire [20:0] z_out_1067_29_9;
  wire [22:0] z_out_1068_29_7;
  wire [22:0] z_out_1069_29_7;
  wire [22:0] z_out_1070_29_7;
  wire [22:0] z_out_1071_29_7;
  wire [22:0] z_out_1072_29_7;
  wire [22:0] z_out_1073_29_7;
  wire [22:0] z_out_1074_29_7;
  wire [22:0] z_out_1075_29_7;
  wire [22:0] z_out_1076_29_7;
  wire [22:0] z_out_1077_29_7;
  wire [22:0] z_out_1078_29_7;
  wire [22:0] z_out_1079_29_7;
  wire [22:0] z_out_1080_29_7;
  wire [22:0] z_out_1081_29_7;
  wire [22:0] z_out_1082_29_7;
  wire [22:0] z_out_1083_29_7;
  wire [22:0] z_out_1084_29_7;
  wire [22:0] z_out_1085_29_7;
  wire [22:0] z_out_1086_29_7;
  wire [22:0] z_out_1087_29_7;
  wire [22:0] z_out_1088_29_7;
  wire [22:0] z_out_1089_29_7;
  wire [22:0] z_out_1090_29_7;
  wire [22:0] z_out_1091_29_7;
  wire [22:0] z_out_1092_29_7;
  wire [22:0] z_out_1093_29_7;
  wire [22:0] z_out_1094_29_7;
  wire [22:0] z_out_1095_29_7;
  wire [22:0] z_out_1096_29_7;
  wire [22:0] z_out_1097_29_7;
  wire [22:0] z_out_1098_29_7;
  wire [22:0] z_out_1099_29_7;
  wire [22:0] z_out_1100_29_7;
  wire [22:0] z_out_1101_29_7;
  wire [22:0] z_out_1102_29_7;
  wire [22:0] z_out_1103_29_7;
  wire [22:0] z_out_1104_29_7;
  wire [22:0] z_out_1105_29_7;
  wire [22:0] z_out_1106_29_7;
  wire [22:0] z_out_1107_29_7;
  wire [22:0] z_out_1108_29_7;
  wire [22:0] z_out_1109_29_7;
  wire [22:0] z_out_1110_29_7;
  wire [22:0] z_out_1111_29_7;
  wire [22:0] z_out_1112_29_7;
  wire [22:0] z_out_1113_29_7;
  wire [22:0] z_out_1114_29_7;
  wire [22:0] z_out_1115_29_7;
  wire [22:0] z_out_1116_29_7;
  wire [22:0] z_out_1117_29_7;
  wire [22:0] z_out_1118_29_7;
  wire [22:0] z_out_1119_29_7;
  wire [22:0] z_out_1120_29_7;
  wire [22:0] z_out_1121_29_7;
  wire [22:0] z_out_1122_29_7;
  wire [22:0] z_out_1123_29_7;
  wire [22:0] z_out_1124_29_7;
  wire [22:0] z_out_1125_29_7;
  wire [22:0] z_out_1126_29_7;
  wire [22:0] z_out_1127_29_7;
  wire [22:0] z_out_1128_29_7;
  wire [22:0] z_out_1129_29_7;
  wire [22:0] z_out_1130_29_7;
  wire [22:0] z_out_1131_29_7;
  wire [20:0] z_out_1132_29_9;
  wire [20:0] z_out_1133_29_9;
  wire [20:0] z_out_1134_29_9;
  wire [20:0] z_out_1135_29_9;
  wire [20:0] z_out_1136_29_9;
  wire [20:0] z_out_1137_29_9;
  wire [20:0] z_out_1138_29_9;
  wire [20:0] z_out_1139_29_9;
  wire [20:0] z_out_1140_29_9;
  wire [20:0] z_out_1141_29_9;
  wire [20:0] z_out_1142_29_9;
  wire [20:0] z_out_1143_29_9;
  wire [20:0] z_out_1144_29_9;
  wire [22:0] z_out_1145_29_7;
  wire [22:0] z_out_1146_29_7;
  wire [22:0] z_out_1147_29_7;
  wire [22:0] z_out_1148_29_7;
  wire [22:0] z_out_1149_29_7;
  wire [22:0] z_out_1150_29_7;
  wire [22:0] z_out_1151_29_7;
  wire [22:0] z_out_1152_29_7;
  wire [22:0] z_out_1153_29_7;
  wire [22:0] z_out_1154_29_7;
  wire [22:0] z_out_1155_29_7;
  wire [22:0] z_out_1156_29_7;
  wire [22:0] z_out_1157_29_7;
  wire [22:0] z_out_1158_29_7;
  wire [22:0] z_out_1159_29_7;
  wire [22:0] z_out_1160_29_7;
  wire [22:0] z_out_1161_29_7;
  wire [22:0] z_out_1162_29_7;
  wire [22:0] z_out_1163_29_7;
  wire [22:0] z_out_1164_29_7;
  wire [22:0] z_out_1165_29_7;
  wire [22:0] z_out_1166_29_7;
  wire [22:0] z_out_1167_29_7;
  wire [22:0] z_out_1168_29_7;
  wire [22:0] z_out_1169_29_7;
  wire [22:0] z_out_1170_29_7;
  wire [22:0] z_out_1171_29_7;
  wire [22:0] z_out_1172_29_7;
  wire [22:0] z_out_1173_29_7;
  wire [22:0] z_out_1174_29_7;
  wire [22:0] z_out_1175_29_7;
  wire [22:0] z_out_1176_29_7;
  wire [22:0] z_out_1177_29_7;
  wire [22:0] z_out_1178_29_7;
  wire [22:0] z_out_1179_29_7;
  wire [22:0] z_out_1180_29_7;
  wire [22:0] z_out_1181_29_7;
  wire [22:0] z_out_1182_29_7;
  wire [22:0] z_out_1183_29_7;
  wire [22:0] z_out_1184_29_7;
  wire [22:0] z_out_1185_29_7;
  wire [22:0] z_out_1186_29_7;
  wire [22:0] z_out_1187_29_7;
  wire [20:0] z_out_1188_29_9;
  wire operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse;
  wire MultLoop_or_22_cse;
  wire AccumDotWidth_or_140_cse;
  wire operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_42_cse;
  wire operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse;
  wire MultLoop_or_81_cse;
  wire AccumDotWidth_or_132_cse_1;
  wire AccumDotWidth_or_153_cse;
  wire AccumDotWidth_or_156_cse;
  wire AccumDotWidth_or_25_cse;
  wire MultLoop_or_87_cse;
  wire AccumDotWidth_or_149_cse;
  wire AccumDotWidth_or_139_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse;
  wire MultLoop_or_89_cse;
  wire AccumDotWidth_or_145_cse;
  wire AccumDotWidth_or_152_cse;
  wire AccumDotWidth_or_150_cse;
  wire AccumDotWidth_or_142_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse;
  wire MultLoop_or_93_cse;
  wire ConvFiltWidth_else_or_730_cse;
  wire ConvFiltWidth_else_or_752_cse;
  wire ConvFiltWidth_else_or_751_cse;
  wire AccumDotWidth_or_157_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse;
  wire AccumDotWidth_or_29_cse;
  wire ConvFiltWidth_else_or_787_cse;
  wire MultLoop_or_17_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_53_cse;
  wire nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse;
  wire AccumDotWidth_or_138_cse;
  wire ConvFiltWidth_else_or_847_cse;
  wire ConvFiltWidth_else_or_849_cse;
  wire ConvFiltWidth_else_or_844_cse;
  wire ConvFiltWidth_else_or_871_cse;
  wire ConvFiltWidth_else_or_861_cse;
  wire ConvFiltWidth_else_or_882_cse;
  wire ConvFiltWidth_else_or_892_cse;
  wire ConvFiltWidth_else_or_1020_cse;
  wire ConvFiltWidth_else_or_1081_cse;
  wire ConvFiltWidth_else_or_1171_cse;
  wire ConvFiltWidth_else_or_987_cse;
  wire AccumDotWidth_or_26_cse;
  wire ConvFiltWidth_else_or_1183_cse;

  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[22:0] nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[20:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[22:0] nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[28:0] MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[28:0] MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire signed [29:0] nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_21_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_22_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_23_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_24_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_25_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_26_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_27_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_28_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_29_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_30_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_31_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_32_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_33_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_34_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux_2_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_35_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_36_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_37_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux_3_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_1_mux_2_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_1_mux_3_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_38_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_operator_22_4_true_AC_TRN_AC_WRAP_mux_1_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_39_nl;
  wire[22:0] operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl;
  wire[23:0] nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl;
  wire[21:0] operator_22_4_true_AC_TRN_AC_WRAP_mux1h_40_nl;
  wire[9:0] AccumDotWidth_mux1h_752_nl;
  wire[7:0] AccumDotWidth_mux1h_753_nl;
  wire[9:0] AccumDotWidth_mux1h_755_nl;
  wire[7:0] AccumDotWidth_mux1h_756_nl;
  wire[9:0] AccumDotWidth_mux1h_757_nl;
  wire[7:0] AccumDotWidth_mux1h_758_nl;
  wire[9:0] AccumDotWidth_mux1h_759_nl;
  wire[7:0] AccumDotWidth_mux1h_760_nl;
  wire[9:0] AccumDotWidth_mux_81_nl;
  wire[9:0] AccumDotWidth_AccumDotWidth_mux_18_nl;
  wire[7:0] AccumDotWidth_AccumDotWidth_mux_19_nl;
  wire[9:0] AccumDotWidth_mux1h_761_nl;
  wire[7:0] AccumDotWidth_AccumDotWidth_mux_20_nl;
  wire[28:0] mul_nl;
  wire signed [29:0] nl_mul_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_332_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_333_nl;
  wire[28:0] mul_1_nl;
  wire signed [29:0] nl_mul_1_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_334_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_335_nl;
  wire[28:0] mul_2_nl;
  wire signed [29:0] nl_mul_2_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_336_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_337_nl;
  wire[28:0] mul_3_nl;
  wire signed [29:0] nl_mul_3_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_338_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_339_nl;
  wire[28:0] mul_4_nl;
  wire signed [29:0] nl_mul_4_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_340_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_341_nl;
  wire[28:0] mul_5_nl;
  wire signed [29:0] nl_mul_5_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_342_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_343_nl;
  wire[28:0] mul_6_nl;
  wire signed [29:0] nl_mul_6_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_344_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_345_nl;
  wire[28:0] mul_7_nl;
  wire signed [29:0] nl_mul_7_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_346_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_347_nl;
  wire[28:0] mul_8_nl;
  wire signed [29:0] nl_mul_8_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_348_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_349_nl;
  wire[28:0] mul_9_nl;
  wire signed [29:0] nl_mul_9_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_350_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_351_nl;
  wire[28:0] mul_10_nl;
  wire signed [29:0] nl_mul_10_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_352_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_353_nl;
  wire[28:0] mul_11_nl;
  wire signed [29:0] nl_mul_11_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_354_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_355_nl;
  wire[28:0] mul_12_nl;
  wire signed [29:0] nl_mul_12_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_356_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_357_nl;
  wire[28:0] mul_13_nl;
  wire signed [29:0] nl_mul_13_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_358_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_359_nl;
  wire[28:0] mul_14_nl;
  wire signed [29:0] nl_mul_14_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_360_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_361_nl;
  wire[28:0] mul_15_nl;
  wire signed [29:0] nl_mul_15_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_362_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_363_nl;
  wire[28:0] mul_16_nl;
  wire signed [29:0] nl_mul_16_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_364_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_365_nl;
  wire[28:0] mul_17_nl;
  wire signed [29:0] nl_mul_17_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_366_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_367_nl;
  wire[28:0] mul_18_nl;
  wire signed [29:0] nl_mul_18_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_368_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_369_nl;
  wire[28:0] mul_19_nl;
  wire signed [29:0] nl_mul_19_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_370_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_371_nl;
  wire[28:0] mul_20_nl;
  wire signed [29:0] nl_mul_20_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_372_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_373_nl;
  wire[28:0] mul_21_nl;
  wire signed [29:0] nl_mul_21_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_374_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_375_nl;
  wire[28:0] mul_22_nl;
  wire signed [29:0] nl_mul_22_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_376_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_377_nl;
  wire[28:0] mul_23_nl;
  wire signed [29:0] nl_mul_23_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_89_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_90_nl;
  wire[28:0] mul_24_nl;
  wire signed [29:0] nl_mul_24_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_91_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_92_nl;
  wire[28:0] mul_25_nl;
  wire signed [29:0] nl_mul_25_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_378_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_379_nl;
  wire[28:0] mul_26_nl;
  wire signed [29:0] nl_mul_26_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_380_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_381_nl;
  wire[28:0] mul_27_nl;
  wire signed [29:0] nl_mul_27_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_382_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_383_nl;
  wire[28:0] mul_28_nl;
  wire signed [29:0] nl_mul_28_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_384_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_385_nl;
  wire[28:0] mul_29_nl;
  wire signed [29:0] nl_mul_29_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_386_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_387_nl;
  wire[28:0] mul_30_nl;
  wire signed [29:0] nl_mul_30_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_388_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_389_nl;
  wire[28:0] mul_31_nl;
  wire signed [29:0] nl_mul_31_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_390_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_391_nl;
  wire[28:0] mul_32_nl;
  wire signed [29:0] nl_mul_32_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_392_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_393_nl;
  wire[28:0] mul_33_nl;
  wire signed [29:0] nl_mul_33_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_394_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_395_nl;
  wire[28:0] mul_34_nl;
  wire signed [29:0] nl_mul_34_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_396_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_397_nl;
  wire[28:0] mul_35_nl;
  wire signed [29:0] nl_mul_35_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_398_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_399_nl;
  wire[28:0] mul_36_nl;
  wire signed [29:0] nl_mul_36_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_400_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_401_nl;
  wire[28:0] mul_37_nl;
  wire signed [29:0] nl_mul_37_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_402_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_403_nl;
  wire[28:0] mul_38_nl;
  wire signed [29:0] nl_mul_38_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_404_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_405_nl;
  wire[28:0] mul_39_nl;
  wire signed [29:0] nl_mul_39_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_406_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_407_nl;
  wire[28:0] mul_40_nl;
  wire signed [29:0] nl_mul_40_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_408_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_409_nl;
  wire[28:0] mul_41_nl;
  wire signed [29:0] nl_mul_41_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_410_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_411_nl;
  wire[28:0] mul_42_nl;
  wire signed [29:0] nl_mul_42_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_412_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_413_nl;
  wire[28:0] mul_43_nl;
  wire signed [29:0] nl_mul_43_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_414_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_415_nl;
  wire[28:0] mul_44_nl;
  wire signed [29:0] nl_mul_44_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_416_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_417_nl;
  wire[28:0] mul_45_nl;
  wire signed [29:0] nl_mul_45_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_418_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_419_nl;
  wire[28:0] mul_46_nl;
  wire signed [29:0] nl_mul_46_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_420_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_421_nl;
  wire[28:0] mul_47_nl;
  wire signed [29:0] nl_mul_47_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_422_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_423_nl;
  wire[28:0] mul_48_nl;
  wire signed [29:0] nl_mul_48_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_424_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_425_nl;
  wire[28:0] mul_49_nl;
  wire signed [29:0] nl_mul_49_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_426_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_427_nl;
  wire[28:0] mul_50_nl;
  wire signed [29:0] nl_mul_50_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_428_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_429_nl;
  wire[28:0] mul_51_nl;
  wire signed [29:0] nl_mul_51_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_93_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_94_nl;
  wire[28:0] mul_52_nl;
  wire signed [29:0] nl_mul_52_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_95_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_96_nl;
  wire[28:0] mul_53_nl;
  wire signed [29:0] nl_mul_53_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_430_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_431_nl;
  wire[28:0] mul_54_nl;
  wire signed [29:0] nl_mul_54_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_432_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_433_nl;
  wire[28:0] mul_55_nl;
  wire signed [29:0] nl_mul_55_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_434_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_435_nl;
  wire[28:0] mul_56_nl;
  wire signed [29:0] nl_mul_56_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_436_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_437_nl;
  wire[28:0] mul_57_nl;
  wire signed [29:0] nl_mul_57_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_438_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_439_nl;
  wire[28:0] mul_58_nl;
  wire signed [29:0] nl_mul_58_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_440_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_441_nl;
  wire[28:0] mul_59_nl;
  wire signed [29:0] nl_mul_59_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_442_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_443_nl;
  wire[28:0] mul_60_nl;
  wire signed [29:0] nl_mul_60_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_444_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_445_nl;
  wire[28:0] mul_61_nl;
  wire signed [29:0] nl_mul_61_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_446_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_447_nl;
  wire[28:0] mul_62_nl;
  wire signed [29:0] nl_mul_62_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_448_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_449_nl;
  wire[28:0] mul_63_nl;
  wire signed [29:0] nl_mul_63_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_450_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_451_nl;
  wire[28:0] mul_64_nl;
  wire signed [29:0] nl_mul_64_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_452_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_453_nl;
  wire[28:0] mul_65_nl;
  wire signed [29:0] nl_mul_65_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_454_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_455_nl;
  wire[28:0] mul_66_nl;
  wire signed [29:0] nl_mul_66_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_456_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_457_nl;
  wire[28:0] mul_67_nl;
  wire signed [29:0] nl_mul_67_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_458_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_459_nl;
  wire[28:0] mul_68_nl;
  wire signed [29:0] nl_mul_68_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_460_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_461_nl;
  wire[28:0] mul_69_nl;
  wire signed [29:0] nl_mul_69_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_462_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_463_nl;
  wire[28:0] mul_70_nl;
  wire signed [29:0] nl_mul_70_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_464_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_465_nl;
  wire[28:0] mul_71_nl;
  wire signed [29:0] nl_mul_71_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_466_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_467_nl;
  wire[28:0] mul_72_nl;
  wire signed [29:0] nl_mul_72_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_468_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_469_nl;
  wire[28:0] mul_73_nl;
  wire signed [29:0] nl_mul_73_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_470_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_471_nl;
  wire[28:0] mul_74_nl;
  wire signed [29:0] nl_mul_74_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_472_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_473_nl;
  wire[28:0] mul_75_nl;
  wire signed [29:0] nl_mul_75_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_474_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_475_nl;
  wire[28:0] mul_76_nl;
  wire signed [29:0] nl_mul_76_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_476_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_477_nl;
  wire[28:0] mul_77_nl;
  wire signed [29:0] nl_mul_77_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_478_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_479_nl;
  wire[28:0] mul_78_nl;
  wire signed [29:0] nl_mul_78_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_480_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_481_nl;
  wire[28:0] mul_79_nl;
  wire signed [29:0] nl_mul_79_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_482_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_483_nl;
  wire[28:0] mul_80_nl;
  wire signed [29:0] nl_mul_80_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_484_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_485_nl;
  wire[28:0] mul_81_nl;
  wire signed [29:0] nl_mul_81_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_486_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_487_nl;
  wire[28:0] mul_82_nl;
  wire signed [29:0] nl_mul_82_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_488_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_489_nl;
  wire[28:0] mul_83_nl;
  wire signed [29:0] nl_mul_83_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_97_nl;
  wire[28:0] mul_84_nl;
  wire signed [29:0] nl_mul_84_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_490_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_491_nl;
  wire[28:0] mul_85_nl;
  wire signed [29:0] nl_mul_85_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_492_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_493_nl;
  wire[28:0] mul_86_nl;
  wire signed [29:0] nl_mul_86_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_494_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_495_nl;
  wire[28:0] mul_87_nl;
  wire signed [29:0] nl_mul_87_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_496_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_497_nl;
  wire[28:0] mul_88_nl;
  wire signed [29:0] nl_mul_88_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_498_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_499_nl;
  wire[28:0] mul_89_nl;
  wire signed [29:0] nl_mul_89_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_500_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_501_nl;
  wire[28:0] mul_90_nl;
  wire signed [29:0] nl_mul_90_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_502_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_503_nl;
  wire[28:0] mul_91_nl;
  wire signed [29:0] nl_mul_91_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_504_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_505_nl;
  wire[28:0] mul_92_nl;
  wire signed [29:0] nl_mul_92_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_506_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_507_nl;
  wire[28:0] mul_93_nl;
  wire signed [29:0] nl_mul_93_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_98_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_99_nl;
  wire[28:0] mul_94_nl;
  wire signed [29:0] nl_mul_94_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_100_nl;
  wire[28:0] mul_95_nl;
  wire signed [29:0] nl_mul_95_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_508_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_509_nl;
  wire[28:0] mul_96_nl;
  wire signed [29:0] nl_mul_96_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_510_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_511_nl;
  wire[28:0] mul_97_nl;
  wire signed [29:0] nl_mul_97_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_512_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_513_nl;
  wire[28:0] mul_98_nl;
  wire signed [29:0] nl_mul_98_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_514_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_515_nl;
  wire[28:0] mul_99_nl;
  wire signed [29:0] nl_mul_99_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_516_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_517_nl;
  wire[28:0] mul_100_nl;
  wire signed [29:0] nl_mul_100_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_518_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_519_nl;
  wire[28:0] mul_101_nl;
  wire signed [29:0] nl_mul_101_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_520_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_521_nl;
  wire[28:0] mul_102_nl;
  wire signed [29:0] nl_mul_102_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_522_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_523_nl;
  wire[28:0] mul_103_nl;
  wire signed [29:0] nl_mul_103_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_524_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_525_nl;
  wire[28:0] mul_104_nl;
  wire signed [29:0] nl_mul_104_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_526_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_527_nl;
  wire[28:0] mul_105_nl;
  wire signed [29:0] nl_mul_105_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_528_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_529_nl;
  wire[28:0] mul_106_nl;
  wire signed [29:0] nl_mul_106_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_530_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_531_nl;
  wire[28:0] mul_107_nl;
  wire signed [29:0] nl_mul_107_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_532_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_533_nl;
  wire[28:0] mul_108_nl;
  wire signed [29:0] nl_mul_108_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_534_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_535_nl;
  wire[28:0] mul_109_nl;
  wire signed [29:0] nl_mul_109_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_536_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_537_nl;
  wire[28:0] mul_110_nl;
  wire signed [29:0] nl_mul_110_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_538_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_539_nl;
  wire[28:0] mul_111_nl;
  wire signed [29:0] nl_mul_111_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_101_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_102_nl;
  wire[28:0] mul_112_nl;
  wire signed [29:0] nl_mul_112_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_103_nl;
  wire[28:0] mul_113_nl;
  wire signed [29:0] nl_mul_113_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_104_nl;
  wire[28:0] mul_114_nl;
  wire signed [29:0] nl_mul_114_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_105_nl;
  wire[28:0] mul_115_nl;
  wire signed [29:0] nl_mul_115_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_540_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_541_nl;
  wire[28:0] mul_116_nl;
  wire signed [29:0] nl_mul_116_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_542_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_543_nl;
  wire[28:0] mul_117_nl;
  wire signed [29:0] nl_mul_117_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_544_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_106_nl;
  wire[28:0] mul_118_nl;
  wire signed [29:0] nl_mul_118_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_545_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_107_nl;
  wire[28:0] mul_119_nl;
  wire signed [29:0] nl_mul_119_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_108_nl;
  wire[28:0] mul_120_nl;
  wire signed [29:0] nl_mul_120_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_109_nl;
  wire[28:0] mul_121_nl;
  wire signed [29:0] nl_mul_121_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_110_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_111_nl;
  wire[28:0] mul_122_nl;
  wire signed [29:0] nl_mul_122_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_546_nl;
  wire[28:0] mul_123_nl;
  wire signed [29:0] nl_mul_123_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_112_nl;
  wire[28:0] mul_124_nl;
  wire signed [29:0] nl_mul_124_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_547_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_113_nl;
  wire[28:0] mul_125_nl;
  wire signed [29:0] nl_mul_125_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_548_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_114_nl;
  wire[28:0] mul_126_nl;
  wire signed [29:0] nl_mul_126_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_549_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_115_nl;
  wire[28:0] mul_127_nl;
  wire signed [29:0] nl_mul_127_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_550_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_116_nl;
  wire[28:0] mul_128_nl;
  wire signed [29:0] nl_mul_128_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_551_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_117_nl;
  wire[28:0] mul_129_nl;
  wire signed [29:0] nl_mul_129_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_118_nl;
  wire[28:0] mul_130_nl;
  wire signed [29:0] nl_mul_130_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_119_nl;
  wire[28:0] mul_131_nl;
  wire signed [29:0] nl_mul_131_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_120_nl;
  wire[28:0] mul_132_nl;
  wire signed [29:0] nl_mul_132_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_552_nl;
  wire[28:0] mul_133_nl;
  wire signed [29:0] nl_mul_133_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_553_nl;
  wire[28:0] mul_134_nl;
  wire signed [29:0] nl_mul_134_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_121_nl;
  wire[28:0] mul_135_nl;
  wire signed [29:0] nl_mul_135_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_554_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_555_nl;
  wire[28:0] mul_136_nl;
  wire signed [29:0] nl_mul_136_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_556_nl;
  wire[28:0] mul_137_nl;
  wire signed [29:0] nl_mul_137_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_557_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_122_nl;
  wire[28:0] mul_138_nl;
  wire signed [29:0] nl_mul_138_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_558_nl;
  wire[28:0] mul_139_nl;
  wire signed [29:0] nl_mul_139_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_559_nl;
  wire[28:0] mul_140_nl;
  wire signed [29:0] nl_mul_140_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_560_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_123_nl;
  wire[28:0] mul_141_nl;
  wire signed [29:0] nl_mul_141_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_561_nl;
  wire[28:0] mul_142_nl;
  wire signed [29:0] nl_mul_142_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_562_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_563_nl;
  wire[28:0] mul_143_nl;
  wire signed [29:0] nl_mul_143_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_564_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_565_nl;
  wire[28:0] mul_144_nl;
  wire signed [29:0] nl_mul_144_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_566_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_124_nl;
  wire[28:0] mul_145_nl;
  wire signed [29:0] nl_mul_145_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_125_nl;
  wire[28:0] mul_146_nl;
  wire signed [29:0] nl_mul_146_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_567_nl;
  wire[28:0] mul_147_nl;
  wire signed [29:0] nl_mul_147_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_126_nl;
  wire[28:0] mul_148_nl;
  wire signed [29:0] nl_mul_148_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_127_nl;
  wire[28:0] mul_149_nl;
  wire signed [29:0] nl_mul_149_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_128_nl;
  wire[28:0] mul_150_nl;
  wire signed [29:0] nl_mul_150_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_129_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_130_nl;
  wire[28:0] mul_151_nl;
  wire signed [29:0] nl_mul_151_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_568_nl;
  wire[28:0] mul_152_nl;
  wire signed [29:0] nl_mul_152_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_569_nl;
  wire[28:0] mul_153_nl;
  wire signed [29:0] nl_mul_153_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_131_nl;
  wire[28:0] mul_154_nl;
  wire signed [29:0] nl_mul_154_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_132_nl;
  wire[28:0] mul_155_nl;
  wire signed [29:0] nl_mul_155_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_570_nl;
  wire[28:0] mul_156_nl;
  wire signed [29:0] nl_mul_156_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_133_nl;
  wire[28:0] mul_157_nl;
  wire signed [29:0] nl_mul_157_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_571_nl;
  wire[28:0] mul_158_nl;
  wire signed [29:0] nl_mul_158_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_572_nl;
  wire[28:0] mul_159_nl;
  wire signed [29:0] nl_mul_159_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_573_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_134_nl;
  wire[21:0] MultLoop_mux1h_310_nl;
  wire[21:0] MultLoop_mux1h_311_nl;
  wire[21:0] MultLoop_mux1h_312_nl;
  wire[21:0] MultLoop_mux1h_313_nl;
  wire[21:0] MultLoop_acc_1290_nl;
  wire[22:0] nl_MultLoop_acc_1290_nl;
  wire[21:0] MultLoop_mux1h_314_nl;
  wire[21:0] MultLoop_mux1h_315_nl;
  wire[21:0] MultLoop_mux1h_316_nl;
  wire[21:0] MultLoop_mux1h_317_nl;
  wire[21:0] MultLoop_mux1h_318_nl;
  wire[21:0] MultLoop_mux1h_319_nl;
  wire[21:0] MultLoop_mux1h_320_nl;
  wire[21:0] MultLoop_mux1h_321_nl;
  wire[21:0] MultLoop_mux1h_322_nl;
  wire[21:0] MultLoop_mux1h_323_nl;
  wire[21:0] MultLoop_mux1h_324_nl;
  wire[21:0] MultLoop_mux1h_325_nl;
  wire[21:0] MultLoop_mux1h_326_nl;
  wire[21:0] MultLoop_mux1h_327_nl;
  wire[21:0] MultLoop_mux1h_328_nl;
  wire[21:0] MultLoop_mux1h_329_nl;
  wire[21:0] MultLoop_mux1h_330_nl;
  wire[21:0] MultLoop_mux1h_331_nl;
  wire[21:0] MultLoop_mux1h_332_nl;
  wire[21:0] MultLoop_mux1h_333_nl;
  wire[28:0] MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux_82_nl;
  wire[21:0] MultLoop_acc_1291_nl;
  wire[22:0] nl_MultLoop_acc_1291_nl;
  wire[21:0] AccumDotWidth_mux_83_nl;
  wire[21:0] MultLoop_acc_1292_nl;
  wire[22:0] nl_MultLoop_acc_1292_nl;
  wire[21:0] MultLoop_mux1h_334_nl;
  wire[21:0] MultLoop_mux1h_335_nl;
  wire[21:0] MultLoop_mux1h_336_nl;
  wire[21:0] MultLoop_mux1h_337_nl;
  wire[21:0] MultLoop_mux1h_338_nl;
  wire[21:0] MultLoop_acc_1293_nl;
  wire[22:0] nl_MultLoop_acc_1293_nl;
  wire[21:0] MultLoop_acc_1294_nl;
  wire[24:0] nl_MultLoop_acc_1294_nl;
  wire[21:0] MultLoop_acc_1304_nl;
  wire[22:0] nl_MultLoop_acc_1304_nl;
  wire[21:0] MultLoop_acc_1305_nl;
  wire[22:0] nl_MultLoop_acc_1305_nl;
  wire[21:0] MultLoop_acc_1297_nl;
  wire[22:0] nl_MultLoop_acc_1297_nl;
  wire[21:0] MultLoop_acc_1298_nl;
  wire[22:0] nl_MultLoop_acc_1298_nl;
  wire[21:0] MultLoop_acc_1300_nl;
  wire[22:0] nl_MultLoop_acc_1300_nl;
  wire[21:0] MultLoop_acc_1301_nl;
  wire[22:0] nl_MultLoop_acc_1301_nl;
  wire[21:0] MultLoop_acc_1307_nl;
  wire[22:0] nl_MultLoop_acc_1307_nl;
  wire[21:0] MultLoop_acc_1308_nl;
  wire[22:0] nl_MultLoop_acc_1308_nl;
  wire[21:0] MultLoop_mux1h_339_nl;
  wire[21:0] MultLoop_mux1h_340_nl;
  wire[21:0] MultLoop_mux1h_341_nl;
  wire[21:0] MultLoop_mux1h_342_nl;
  wire[21:0] MultLoop_mux1h_343_nl;
  wire[21:0] MultLoop_mux1h_344_nl;
  wire[21:0] MultLoop_mux1h_345_nl;
  wire[21:0] MultLoop_mux1h_346_nl;
  wire[21:0] MultLoop_mux1h_347_nl;
  wire[21:0] MultLoop_acc_1309_nl;
  wire[23:0] nl_MultLoop_acc_1309_nl;
  wire[21:0] MultLoop_acc_1310_nl;
  wire[22:0] nl_MultLoop_acc_1310_nl;
  wire[21:0] MultLoop_acc_1311_nl;
  wire[22:0] nl_MultLoop_acc_1311_nl;
  wire[21:0] MultLoop_acc_1312_nl;
  wire[22:0] nl_MultLoop_acc_1312_nl;
  wire[21:0] MultLoop_acc_1315_nl;
  wire[22:0] nl_MultLoop_acc_1315_nl;
  wire[21:0] MultLoop_acc_1316_nl;
  wire[22:0] nl_MultLoop_acc_1316_nl;
  wire[21:0] MultLoop_mux1h_348_nl;
  wire[21:0] MultLoop_mux1h_349_nl;
  wire[21:0] MultLoop_mux1h_350_nl;
  wire[21:0] MultLoop_mux1h_351_nl;
  wire[21:0] MultLoop_acc_1317_nl;
  wire[22:0] nl_MultLoop_acc_1317_nl;
  wire[21:0] MultLoop_acc_1318_nl;
  wire[22:0] nl_MultLoop_acc_1318_nl;
  wire[21:0] MultLoop_mux1h_352_nl;
  wire[21:0] MultLoop_acc_1319_nl;
  wire[22:0] nl_MultLoop_acc_1319_nl;
  wire[21:0] MultLoop_acc_1320_nl;
  wire[22:0] nl_MultLoop_acc_1320_nl;
  wire[21:0] MultLoop_mux1h_353_nl;
  wire[21:0] MultLoop_acc_1321_nl;
  wire[22:0] nl_MultLoop_acc_1321_nl;
  wire[21:0] MultLoop_acc_1322_nl;
  wire[22:0] nl_MultLoop_acc_1322_nl;
  wire[21:0] MultLoop_acc_1323_nl;
  wire[22:0] nl_MultLoop_acc_1323_nl;
  wire[21:0] MultLoop_mux1h_354_nl;
  wire[21:0] MultLoop_mux1h_355_nl;
  wire[21:0] MultLoop_mux1h_356_nl;
  wire[21:0] MultLoop_MultLoop_mux_10_nl;
  wire[21:0] MultLoop_mux1h_357_nl;
  wire[21:0] MultLoop_MultLoop_mux_11_nl;
  wire[21:0] MultLoop_mux1h_358_nl;
  wire[21:0] MultLoop_acc_1324_nl;
  wire[22:0] nl_MultLoop_acc_1324_nl;
  wire[21:0] MultLoop_acc_1325_nl;
  wire[22:0] nl_MultLoop_acc_1325_nl;
  wire[21:0] MultLoop_mux1h_359_nl;
  wire[21:0] MultLoop_acc_1326_nl;
  wire[22:0] nl_MultLoop_acc_1326_nl;
  wire[21:0] MultLoop_mux1h_360_nl;
  wire[21:0] MultLoop_mux1h_361_nl;
  wire[21:0] MultLoop_acc_1327_nl;
  wire[22:0] nl_MultLoop_acc_1327_nl;
  wire[21:0] MultLoop_acc_1328_nl;
  wire[24:0] nl_MultLoop_acc_1328_nl;
  wire[21:0] MultLoop_acc_1335_nl;
  wire[22:0] nl_MultLoop_acc_1335_nl;
  wire[21:0] MultLoop_acc_1336_nl;
  wire[22:0] nl_MultLoop_acc_1336_nl;
  wire[28:0] MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1331_nl;
  wire[22:0] nl_MultLoop_acc_1331_nl;
  wire[21:0] MultLoop_acc_1332_nl;
  wire[22:0] nl_MultLoop_acc_1332_nl;
  wire[21:0] MultLoop_acc_1338_nl;
  wire[22:0] nl_MultLoop_acc_1338_nl;
  wire[28:0] MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1339_nl;
  wire[22:0] nl_MultLoop_acc_1339_nl;
  wire[28:0] MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_362_nl;
  wire[21:0] MultLoop_mux1h_363_nl;
  wire[21:0] MultLoop_mux_78_nl;
  wire[21:0] MultLoop_mux_79_nl;
  wire[21:0] MultLoop_MultLoop_mux_12_nl;
  wire[21:0] MultLoop_MultLoop_mux_13_nl;
  wire[21:0] MultLoop_mux1h_364_nl;
  wire[21:0] MultLoop_mux1h_365_nl;
  wire[21:0] MultLoop_mux1h_366_nl;
  wire[21:0] MultLoop_acc_1340_nl;
  wire[22:0] nl_MultLoop_acc_1340_nl;
  wire[21:0] MultLoop_mux1h_367_nl;
  wire[21:0] AccumDotWidth_mux1h_762_nl;
  wire[21:0] AccumDotWidth_mux1h_763_nl;
  wire[21:0] AccumDotWidth_mux1h_764_nl;
  wire[21:0] AccumDotWidth_mux1h_765_nl;
  wire[21:0] AccumDotWidth_mux1h_766_nl;
  wire[21:0] MultLoop_acc_1341_nl;
  wire[22:0] nl_MultLoop_acc_1341_nl;
  wire[21:0] AccumDotWidth_mux1h_767_nl;
  wire[21:0] MultLoop_mux_80_nl;
  wire[21:0] MultLoop_mux_81_nl;
  wire[21:0] MultLoop_mux_82_nl;
  wire[21:0] MultLoop_mux_83_nl;
  wire[21:0] MultLoop_mux1h_368_nl;
  wire[21:0] MultLoop_mux1h_369_nl;
  wire[21:0] MultLoop_mux1h_370_nl;
  wire[21:0] MultLoop_acc_1342_nl;
  wire[22:0] nl_MultLoop_acc_1342_nl;
  wire[21:0] MultLoop_acc_1343_nl;
  wire[22:0] nl_MultLoop_acc_1343_nl;
  wire[21:0] MultLoop_acc_1344_nl;
  wire[23:0] nl_MultLoop_acc_1344_nl;
  wire[21:0] MultLoop_acc_1346_nl;
  wire[22:0] nl_MultLoop_acc_1346_nl;
  wire[28:0] MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1347_nl;
  wire[22:0] nl_MultLoop_acc_1347_nl;
  wire[28:0] MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1349_nl;
  wire[22:0] nl_MultLoop_acc_1349_nl;
  wire[28:0] MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1350_nl;
  wire[22:0] nl_MultLoop_acc_1350_nl;
  wire[28:0] MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_371_nl;
  wire[28:0] MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1351_nl;
  wire[23:0] nl_MultLoop_acc_1351_nl;
  wire[21:0] MultLoop_acc_1353_nl;
  wire[22:0] nl_MultLoop_acc_1353_nl;
  wire[21:0] MultLoop_acc_1354_nl;
  wire[22:0] nl_MultLoop_acc_1354_nl;
  wire[21:0] MultLoop_acc_1355_nl;
  wire[22:0] nl_MultLoop_acc_1355_nl;
  wire[21:0] AccumDotWidth_mux1h_768_nl;
  wire[21:0] AccumDotWidth_mux1h_769_nl;
  wire[21:0] AccumDotWidth_mux1h_770_nl;
  wire[21:0] AccumDotWidth_mux1h_771_nl;
  wire[21:0] AccumDotWidth_mux1h_772_nl;
  wire[21:0] AccumDotWidth_acc_2401_nl;
  wire[22:0] nl_AccumDotWidth_acc_2401_nl;
  wire[21:0] AccumDotWidth_mux1h_773_nl;
  wire[21:0] AccumDotWidth_mux1h_774_nl;
  wire[21:0] AccumDotWidth_mux1h_775_nl;
  wire[21:0] MultLoop_acc_1356_nl;
  wire[22:0] nl_MultLoop_acc_1356_nl;
  wire[21:0] AccumDotWidth_mux1h_776_nl;
  wire[21:0] MultLoop_acc_1357_nl;
  wire[22:0] nl_MultLoop_acc_1357_nl;
  wire[21:0] AccumDotWidth_mux1h_777_nl;
  wire[21:0] AccumDotWidth_mux_84_nl;
  wire[21:0] MultLoop_acc_1358_nl;
  wire[22:0] nl_MultLoop_acc_1358_nl;
  wire[21:0] AccumDotWidth_mux_85_nl;
  wire[21:0] MultLoop_acc_1359_nl;
  wire[22:0] nl_MultLoop_acc_1359_nl;
  wire[21:0] AccumDotWidth_mux1h_778_nl;
  wire[21:0] MultLoop_acc_1360_nl;
  wire[22:0] nl_MultLoop_acc_1360_nl;
  wire[21:0] AccumDotWidth_mux1h_779_nl;
  wire[21:0] MultLoop_acc_1361_nl;
  wire[22:0] nl_MultLoop_acc_1361_nl;
  wire[21:0] AccumDotWidth_mux1h_780_nl;
  wire[21:0] MultLoop_acc_1362_nl;
  wire[22:0] nl_MultLoop_acc_1362_nl;
  wire[21:0] AccumDotWidth_mux1h_781_nl;
  wire[21:0] MultLoop_acc_1363_nl;
  wire[22:0] nl_MultLoop_acc_1363_nl;
  wire[21:0] AccumDotWidth_mux1h_782_nl;
  wire[21:0] AccumDotWidth_mux1h_783_nl;
  wire[21:0] AccumDotWidth_mux_86_nl;
  wire[21:0] AccumDotWidth_mux_87_nl;
  wire[21:0] AccumDotWidth_mux1h_784_nl;
  wire[21:0] AccumDotWidth_acc_2402_nl;
  wire[22:0] nl_AccumDotWidth_acc_2402_nl;
  wire[21:0] AccumDotWidth_mux1h_785_nl;
  wire[21:0] AccumDotWidth_acc_2403_nl;
  wire[22:0] nl_AccumDotWidth_acc_2403_nl;
  wire[21:0] AccumDotWidth_mux1h_786_nl;
  wire[21:0] AccumDotWidth_mux1h_787_nl;
  wire[21:0] AccumDotWidth_mux_88_nl;
  wire[21:0] MultLoop_acc_1364_nl;
  wire[22:0] nl_MultLoop_acc_1364_nl;
  wire[21:0] AccumDotWidth_mux_89_nl;
  wire[21:0] MultLoop_acc_1365_nl;
  wire[22:0] nl_MultLoop_acc_1365_nl;
  wire[21:0] AccumDotWidth_mux1h_788_nl;
  wire[21:0] AccumDotWidth_mux1h_789_nl;
  wire[21:0] AccumDotWidth_mux_90_nl;
  wire[21:0] AccumDotWidth_mux_91_nl;
  wire[21:0] AccumDotWidth_mux1h_790_nl;
  wire[21:0] AccumDotWidth_acc_2404_nl;
  wire[22:0] nl_AccumDotWidth_acc_2404_nl;
  wire[21:0] AccumDotWidth_mux1h_791_nl;
  wire[21:0] AccumDotWidth_mux1h_792_nl;
  wire[21:0] AccumDotWidth_mux1h_793_nl;
  wire[21:0] AccumDotWidth_mux1h_794_nl;
  wire[21:0] AccumDotWidth_mux1h_795_nl;
  wire[21:0] AccumDotWidth_mux1h_796_nl;
  wire[21:0] AccumDotWidth_mux1h_797_nl;
  wire[21:0] AccumDotWidth_mux1h_798_nl;
  wire[21:0] AccumDotWidth_mux1h_799_nl;
  wire[21:0] AccumDotWidth_acc_2405_nl;
  wire[22:0] nl_AccumDotWidth_acc_2405_nl;
  wire[21:0] AccumDotWidth_mux1h_800_nl;
  wire[21:0] AccumDotWidth_mux1h_801_nl;
  wire[21:0] AccumDotWidth_mux1h_802_nl;
  wire[21:0] AccumDotWidth_mux1h_803_nl;
  wire[21:0] AccumDotWidth_mux1h_804_nl;
  wire[21:0] AccumDotWidth_mux1h_805_nl;
  wire[21:0] AccumDotWidth_mux1h_806_nl;
  wire[21:0] AccumDotWidth_mux1h_807_nl;
  wire[21:0] AccumDotWidth_mux1h_808_nl;
  wire[21:0] AccumDotWidth_acc_2406_nl;
  wire[22:0] nl_AccumDotWidth_acc_2406_nl;
  wire[21:0] AccumDotWidth_mux1h_809_nl;
  wire[21:0] AccumDotWidth_acc_2407_nl;
  wire[22:0] nl_AccumDotWidth_acc_2407_nl;
  wire[21:0] AccumDotWidth_mux1h_810_nl;
  wire[21:0] AccumDotWidth_mux1h_811_nl;
  wire[21:0] AccumDotWidth_mux1h_812_nl;
  wire[21:0] AccumDotWidth_mux1h_813_nl;
  wire[21:0] AccumDotWidth_mux1h_814_nl;
  wire[21:0] AccumDotWidth_mux1h_815_nl;
  wire[21:0] AccumDotWidth_mux1h_816_nl;
  wire[0:0] AccumDotWidth_or_151_nl;
  wire[21:0] AccumDotWidth_mux1h_817_nl;
  wire[21:0] MultLoop_acc_1366_nl;
  wire[22:0] nl_MultLoop_acc_1366_nl;
  wire[28:0] MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_818_nl;
  wire[21:0] AccumDotWidth_mux1h_819_nl;
  wire[21:0] AccumDotWidth_mux1h_820_nl;
  wire[21:0] AccumDotWidth_acc_2408_nl;
  wire[22:0] nl_AccumDotWidth_acc_2408_nl;
  wire[21:0] MultLoop_acc_1367_nl;
  wire[22:0] nl_MultLoop_acc_1367_nl;
  wire[21:0] MultLoop_acc_1368_nl;
  wire[22:0] nl_MultLoop_acc_1368_nl;
  wire[21:0] AccumDotWidth_mux1h_821_nl;
  wire[21:0] MultLoop_acc_1369_nl;
  wire[22:0] nl_MultLoop_acc_1369_nl;
  wire[21:0] AccumDotWidth_mux1h_822_nl;
  wire[21:0] AccumDotWidth_acc_2409_nl;
  wire[22:0] nl_AccumDotWidth_acc_2409_nl;
  wire[21:0] AccumDotWidth_mux1h_823_nl;
  wire[21:0] AccumDotWidth_acc_2410_nl;
  wire[22:0] nl_AccumDotWidth_acc_2410_nl;
  wire[21:0] AccumDotWidth_acc_2411_nl;
  wire[22:0] nl_AccumDotWidth_acc_2411_nl;
  wire[21:0] AccumDotWidth_mux1h_824_nl;
  wire[21:0] MultLoop_acc_1370_nl;
  wire[22:0] nl_MultLoop_acc_1370_nl;
  wire[21:0] AccumDotWidth_mux1h_825_nl;
  wire[21:0] MultLoop_acc_1371_nl;
  wire[22:0] nl_MultLoop_acc_1371_nl;
  wire[21:0] AccumDotWidth_mux1h_826_nl;
  wire[21:0] MultLoop_acc_1372_nl;
  wire[22:0] nl_MultLoop_acc_1372_nl;
  wire[21:0] AccumDotWidth_mux1h_827_nl;
  wire[21:0] MultLoop_acc_1373_nl;
  wire[22:0] nl_MultLoop_acc_1373_nl;
  wire[21:0] MultLoop_mux1h_372_nl;
  wire[21:0] MultLoop_mux1h_373_nl;
  wire[21:0] AccumDotWidth_mux1h_828_nl;
  wire[21:0] AccumDotWidth_mux1h_829_nl;
  wire[21:0] AccumDotWidth_mux1h_830_nl;
  wire[21:0] AccumDotWidth_acc_2412_nl;
  wire[22:0] nl_AccumDotWidth_acc_2412_nl;
  wire[21:0] AccumDotWidth_mux1h_831_nl;
  wire[21:0] AccumDotWidth_mux1h_832_nl;
  wire[21:0] AccumDotWidth_acc_2413_nl;
  wire[22:0] nl_AccumDotWidth_acc_2413_nl;
  wire[21:0] AccumDotWidth_mux1h_833_nl;
  wire[21:0] MultLoop_mux1h_374_nl;
  wire[28:0] MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_375_nl;
  wire[21:0] MultLoop_acc_1374_nl;
  wire[22:0] nl_MultLoop_acc_1374_nl;
  wire[21:0] AccumDotWidth_mux1h_834_nl;
  wire[21:0] AccumDotWidth_mux1h_835_nl;
  wire[21:0] AccumDotWidth_mux1h_836_nl;
  wire[21:0] MultLoop_acc_1375_nl;
  wire[22:0] nl_MultLoop_acc_1375_nl;
  wire[21:0] MultLoop_acc_1376_nl;
  wire[22:0] nl_MultLoop_acc_1376_nl;
  wire[21:0] AccumDotWidth_mux1h_837_nl;
  wire[21:0] MultLoop_acc_1377_nl;
  wire[22:0] nl_MultLoop_acc_1377_nl;
  wire[21:0] MultLoop_acc_1378_nl;
  wire[22:0] nl_MultLoop_acc_1378_nl;
  wire[21:0] AccumDotWidth_mux1h_838_nl;
  wire[21:0] MultLoop_acc_1379_nl;
  wire[22:0] nl_MultLoop_acc_1379_nl;
  wire[21:0] MultLoop_acc_1380_nl;
  wire[22:0] nl_MultLoop_acc_1380_nl;
  wire[21:0] AccumDotWidth_mux1h_839_nl;
  wire[21:0] MultLoop_mux1h_376_nl;
  wire[21:0] MultLoop_mux1h_377_nl;
  wire[21:0] MultLoop_mux1h_378_nl;
  wire[21:0] MultLoop_mux1h_379_nl;
  wire[21:0] MultLoop_mux_84_nl;
  wire[21:0] MultLoop_acc_1381_nl;
  wire[22:0] nl_MultLoop_acc_1381_nl;
  wire[21:0] MultLoop_mux1h_380_nl;
  wire[21:0] MultLoop_mux1h_381_nl;
  wire[21:0] MultLoop_mux_85_nl;
  wire[21:0] MultLoop_mux_86_nl;
  wire[21:0] MultLoop_acc_1382_nl;
  wire[22:0] nl_MultLoop_acc_1382_nl;
  wire[21:0] MultLoop_mux_87_nl;
  wire[21:0] MultLoop_mux1h_382_nl;
  wire[21:0] MultLoop_mux1h_383_nl;
  wire[21:0] MultLoop_mux1h_384_nl;
  wire[21:0] MultLoop_mux1h_385_nl;
  wire[21:0] MultLoop_acc_1383_nl;
  wire[22:0] nl_MultLoop_acc_1383_nl;
  wire[21:0] MultLoop_mux1h_386_nl;
  wire[21:0] MultLoop_mux1h_387_nl;
  wire[21:0] MultLoop_mux1h_388_nl;
  wire[21:0] MultLoop_mux1h_389_nl;
  wire[21:0] MultLoop_mux_88_nl;
  wire[21:0] MultLoop_acc_1384_nl;
  wire[22:0] nl_MultLoop_acc_1384_nl;
  wire[21:0] MultLoop_acc_1385_nl;
  wire[22:0] nl_MultLoop_acc_1385_nl;
  wire[21:0] MultLoop_acc_1386_nl;
  wire[22:0] nl_MultLoop_acc_1386_nl;
  wire[21:0] MultLoop_mux1h_390_nl;
  wire[21:0] MultLoop_mux1h_391_nl;
  wire[21:0] MultLoop_mux1h_392_nl;
  wire[21:0] MultLoop_acc_1387_nl;
  wire[22:0] nl_MultLoop_acc_1387_nl;
  wire[21:0] MultLoop_mux1h_393_nl;
  wire[21:0] MultLoop_acc_1388_nl;
  wire[22:0] nl_MultLoop_acc_1388_nl;
  wire[21:0] MultLoop_mux1h_394_nl;
  wire[21:0] MultLoop_acc_1389_nl;
  wire[22:0] nl_MultLoop_acc_1389_nl;
  wire[21:0] MultLoop_mux1h_395_nl;
  wire[21:0] MultLoop_acc_1390_nl;
  wire[22:0] nl_MultLoop_acc_1390_nl;
  wire[21:0] MultLoop_mux1h_396_nl;
  wire[21:0] MultLoop_mux1h_397_nl;
  wire[21:0] MultLoop_acc_1391_nl;
  wire[22:0] nl_MultLoop_acc_1391_nl;
  wire[21:0] MultLoop_acc_1392_nl;
  wire[22:0] nl_MultLoop_acc_1392_nl;
  wire[21:0] MultLoop_mux1h_398_nl;
  wire[21:0] MultLoop_mux1h_399_nl;
  wire[21:0] MultLoop_mux1h_400_nl;
  wire[21:0] MultLoop_acc_1393_nl;
  wire[22:0] nl_MultLoop_acc_1393_nl;
  wire[21:0] MultLoop_acc_1394_nl;
  wire[22:0] nl_MultLoop_acc_1394_nl;
  wire[21:0] MultLoop_mux1h_401_nl;
  wire[21:0] MultLoop_acc_1395_nl;
  wire[22:0] nl_MultLoop_acc_1395_nl;
  wire[21:0] MultLoop_mux1h_402_nl;
  wire[21:0] MultLoop_mux1h_403_nl;
  wire[21:0] MultLoop_mux1h_404_nl;
  wire[21:0] MultLoop_acc_1396_nl;
  wire[22:0] nl_MultLoop_acc_1396_nl;
  wire[21:0] MultLoop_mux1h_405_nl;
  wire[21:0] MultLoop_mux1h_406_nl;
  wire[21:0] MultLoop_mux1h_407_nl;
  wire[21:0] MultLoop_mux1h_408_nl;
  wire[21:0] MultLoop_mux1h_409_nl;
  wire[21:0] MultLoop_mux1h_410_nl;
  wire[21:0] MultLoop_mux1h_411_nl;
  wire[21:0] MultLoop_mux1h_412_nl;
  wire[21:0] MultLoop_acc_1397_nl;
  wire[22:0] nl_MultLoop_acc_1397_nl;
  wire[21:0] MultLoop_acc_1398_nl;
  wire[22:0] nl_MultLoop_acc_1398_nl;
  wire[21:0] MultLoop_mux1h_413_nl;
  wire[21:0] MultLoop_acc_1399_nl;
  wire[22:0] nl_MultLoop_acc_1399_nl;
  wire[21:0] MultLoop_acc_1400_nl;
  wire[22:0] nl_MultLoop_acc_1400_nl;
  wire[21:0] MultLoop_acc_1401_nl;
  wire[22:0] nl_MultLoop_acc_1401_nl;
  wire[21:0] MultLoop_mux1h_414_nl;
  wire[21:0] MultLoop_mux1h_415_nl;
  wire[21:0] MultLoop_mux1h_416_nl;
  wire[21:0] MultLoop_acc_1402_nl;
  wire[22:0] nl_MultLoop_acc_1402_nl;
  wire[21:0] MultLoop_acc_1403_nl;
  wire[24:0] nl_MultLoop_acc_1403_nl;
  wire[21:0] MultLoop_acc_1413_nl;
  wire[22:0] nl_MultLoop_acc_1413_nl;
  wire[28:0] MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1414_nl;
  wire[22:0] nl_MultLoop_acc_1414_nl;
  wire[28:0] MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1406_nl;
  wire[22:0] nl_MultLoop_acc_1406_nl;
  wire[28:0] MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1407_nl;
  wire[22:0] nl_MultLoop_acc_1407_nl;
  wire[28:0] MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1409_nl;
  wire[22:0] nl_MultLoop_acc_1409_nl;
  wire[28:0] MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1410_nl;
  wire[22:0] nl_MultLoop_acc_1410_nl;
  wire[28:0] MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1416_nl;
  wire[22:0] nl_MultLoop_acc_1416_nl;
  wire[28:0] MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1417_nl;
  wire[22:0] nl_MultLoop_acc_1417_nl;
  wire[28:0] MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_417_nl;
  wire[21:0] MultLoop_mux1h_418_nl;
  wire[21:0] MultLoop_mux1h_419_nl;
  wire[21:0] MultLoop_mux1h_420_nl;
  wire[21:0] MultLoop_mux1h_421_nl;
  wire[21:0] MultLoop_mux1h_422_nl;
  wire[21:0] MultLoop_mux1h_423_nl;
  wire[21:0] MultLoop_acc_1418_nl;
  wire[22:0] nl_MultLoop_acc_1418_nl;
  wire[21:0] MultLoop_acc_1419_nl;
  wire[22:0] nl_MultLoop_acc_1419_nl;
  wire[21:0] MultLoop_mux1h_424_nl;
  wire[21:0] MultLoop_mux1h_425_nl;
  wire[21:0] MultLoop_mux1h_426_nl;
  wire[21:0] MultLoop_mux1h_427_nl;
  wire[21:0] MultLoop_mux1h_428_nl;
  wire[21:0] MultLoop_mux1h_429_nl;
  wire[21:0] AccumDotWidth_mux1h_840_nl;
  wire[21:0] AccumDotWidth_mux1h_841_nl;
  wire[21:0] AccumDotWidth_mux1h_842_nl;
  wire[21:0] AccumDotWidth_mux1h_843_nl;
  wire[21:0] AccumDotWidth_mux1h_844_nl;
  wire[21:0] AccumDotWidth_mux1h_845_nl;
  wire[21:0] AccumDotWidth_acc_2414_nl;
  wire[22:0] nl_AccumDotWidth_acc_2414_nl;
  wire[9:0] AccumDotWidth_acc_2415_nl;
  wire[10:0] nl_AccumDotWidth_acc_2415_nl;
  wire[21:0] AccumDotWidth_mux1h_846_nl;
  wire[21:0] AccumDotWidth_acc_2416_nl;
  wire[22:0] nl_AccumDotWidth_acc_2416_nl;
  wire[21:0] AccumDotWidth_mux1h_847_nl;
  wire[21:0] AccumDotWidth_acc_2417_nl;
  wire[22:0] nl_AccumDotWidth_acc_2417_nl;
  wire[21:0] AccumDotWidth_mux1h_848_nl;
  wire[21:0] AccumDotWidth_acc_2418_nl;
  wire[22:0] nl_AccumDotWidth_acc_2418_nl;
  wire[21:0] AccumDotWidth_mux1h_849_nl;
  wire[21:0] AccumDotWidth_acc_2419_nl;
  wire[22:0] nl_AccumDotWidth_acc_2419_nl;
  wire[21:0] AccumDotWidth_mux_92_nl;
  wire[21:0] AccumDotWidth_mux_93_nl;
  wire[21:0] AccumDotWidth_mux1h_850_nl;
  wire[21:0] AccumDotWidth_mux1h_851_nl;
  wire[21:0] AccumDotWidth_mux1h_852_nl;
  wire[21:0] AccumDotWidth_acc_2420_nl;
  wire[22:0] nl_AccumDotWidth_acc_2420_nl;
  wire[21:0] AccumDotWidth_mux1h_853_nl;
  wire[21:0] AccumDotWidth_acc_2421_nl;
  wire[22:0] nl_AccumDotWidth_acc_2421_nl;
  wire[21:0] AccumDotWidth_mux1h_854_nl;
  wire[21:0] AccumDotWidth_acc_2422_nl;
  wire[22:0] nl_AccumDotWidth_acc_2422_nl;
  wire[21:0] AccumDotWidth_mux1h_855_nl;
  wire[21:0] AccumDotWidth_acc_2423_nl;
  wire[22:0] nl_AccumDotWidth_acc_2423_nl;
  wire[21:0] AccumDotWidth_mux1h_856_nl;
  wire[21:0] AccumDotWidth_mux1h_857_nl;
  wire[21:0] AccumDotWidth_mux1h_858_nl;
  wire[21:0] AccumDotWidth_mux1h_859_nl;
  wire[21:0] MultLoop_acc_1420_nl;
  wire[22:0] nl_MultLoop_acc_1420_nl;
  wire[21:0] AccumDotWidth_mux1h_860_nl;
  wire[21:0] AccumDotWidth_mux1h_861_nl;
  wire[21:0] AccumDotWidth_mux1h_862_nl;
  wire[21:0] AccumDotWidth_mux1h_863_nl;
  wire[21:0] AccumDotWidth_mux1h_864_nl;
  wire[21:0] AccumDotWidth_mux1h_865_nl;
  wire[21:0] MultLoop_acc_1421_nl;
  wire[22:0] nl_MultLoop_acc_1421_nl;
  wire[21:0] AccumDotWidth_mux1h_866_nl;
  wire[21:0] AccumDotWidth_mux1h_867_nl;
  wire[21:0] MultLoop_acc_1422_nl;
  wire[22:0] nl_MultLoop_acc_1422_nl;
  wire[21:0] AccumDotWidth_mux1h_868_nl;
  wire[21:0] MultLoop_acc_1423_nl;
  wire[22:0] nl_MultLoop_acc_1423_nl;
  wire[21:0] AccumDotWidth_mux1h_869_nl;
  wire[21:0] AccumDotWidth_mux1h_870_nl;
  wire[21:0] AccumDotWidth_mux1h_871_nl;
  wire[21:0] AccumDotWidth_mux_94_nl;
  wire[21:0] AccumDotWidth_mux_95_nl;
  wire[21:0] AccumDotWidth_mux1h_872_nl;
  wire[21:0] AccumDotWidth_mux1h_873_nl;
  wire[21:0] MultLoop_acc_1424_nl;
  wire[22:0] nl_MultLoop_acc_1424_nl;
  wire[21:0] AccumDotWidth_mux1h_874_nl;
  wire[21:0] MultLoop_acc_1425_nl;
  wire[22:0] nl_MultLoop_acc_1425_nl;
  wire[21:0] AccumDotWidth_mux1h_875_nl;
  wire[21:0] MultLoop_acc_1426_nl;
  wire[22:0] nl_MultLoop_acc_1426_nl;
  wire[21:0] AccumDotWidth_mux1h_876_nl;
  wire[21:0] MultLoop_acc_1427_nl;
  wire[22:0] nl_MultLoop_acc_1427_nl;
  wire[21:0] AccumDotWidth_mux1h_877_nl;
  wire[21:0] MultLoop_acc_1428_nl;
  wire[22:0] nl_MultLoop_acc_1428_nl;
  wire[21:0] AccumDotWidth_mux1h_878_nl;
  wire[21:0] MultLoop_acc_1429_nl;
  wire[22:0] nl_MultLoop_acc_1429_nl;
  wire[10:0] AccumDotWidth_mux1h_879_nl;
  wire[9:0] AccumDotWidth_acc_2424_nl;
  wire[10:0] nl_AccumDotWidth_acc_2424_nl;
  wire[9:0] AccumDotWidth_acc_2425_nl;
  wire[10:0] nl_AccumDotWidth_acc_2425_nl;
  wire[9:0] AccumDotWidth_acc_2426_nl;
  wire[10:0] nl_AccumDotWidth_acc_2426_nl;
  wire[9:0] AccumDotWidth_acc_2427_nl;
  wire[10:0] nl_AccumDotWidth_acc_2427_nl;
  wire[10:0] AccumDotWidth_mux1h_880_nl;
  wire[21:0] AccumDotWidth_mux1h_881_nl;
  wire[21:0] AccumDotWidth_acc_2428_nl;
  wire[22:0] nl_AccumDotWidth_acc_2428_nl;
  wire[21:0] MultLoop_acc_1430_nl;
  wire[22:0] nl_MultLoop_acc_1430_nl;
  wire[21:0] AccumDotWidth_mux1h_882_nl;
  wire[21:0] AccumDotWidth_acc_2429_nl;
  wire[22:0] nl_AccumDotWidth_acc_2429_nl;
  wire[9:0] AccumDotWidth_acc_2430_nl;
  wire[10:0] nl_AccumDotWidth_acc_2430_nl;
  wire[21:0] MultLoop_acc_1431_nl;
  wire[22:0] nl_MultLoop_acc_1431_nl;
  wire[21:0] AccumDotWidth_mux1h_883_nl;
  wire[21:0] AccumDotWidth_mux1h_884_nl;
  wire[21:0] MultLoop_acc_1432_nl;
  wire[22:0] nl_MultLoop_acc_1432_nl;
  wire[28:0] MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_885_nl;
  wire[21:0] AccumDotWidth_acc_2431_nl;
  wire[22:0] nl_AccumDotWidth_acc_2431_nl;
  wire[21:0] MultLoop_acc_1433_nl;
  wire[22:0] nl_MultLoop_acc_1433_nl;
  wire[10:0] AccumDotWidth_mux1h_886_nl;
  wire[9:0] AccumDotWidth_acc_2432_nl;
  wire[10:0] nl_AccumDotWidth_acc_2432_nl;
  wire[9:0] AccumDotWidth_acc_2433_nl;
  wire[10:0] nl_AccumDotWidth_acc_2433_nl;
  wire[9:0] AccumDotWidth_acc_2434_nl;
  wire[10:0] nl_AccumDotWidth_acc_2434_nl;
  wire[9:0] AccumDotWidth_acc_2435_nl;
  wire[10:0] nl_AccumDotWidth_acc_2435_nl;
  wire[10:0] AccumDotWidth_mux1h_887_nl;
  wire[21:0] AccumDotWidth_mux1h_888_nl;
  wire[21:0] AccumDotWidth_mux1h_889_nl;
  wire[21:0] MultLoop_acc_1434_nl;
  wire[22:0] nl_MultLoop_acc_1434_nl;
  wire[21:0] AccumDotWidth_mux1h_890_nl;
  wire[21:0] AccumDotWidth_mux1h_891_nl;
  wire[21:0] AccumDotWidth_mux1h_892_nl;
  wire[21:0] MultLoop_acc_1435_nl;
  wire[22:0] nl_MultLoop_acc_1435_nl;
  wire[21:0] AccumDotWidth_mux1h_893_nl;
  wire[21:0] MultLoop_acc_1436_nl;
  wire[22:0] nl_MultLoop_acc_1436_nl;
  wire[28:0] MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_894_nl;
  wire[21:0] MultLoop_acc_1437_nl;
  wire[22:0] nl_MultLoop_acc_1437_nl;
  wire[28:0] MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_895_nl;
  wire[21:0] MultLoop_acc_1438_nl;
  wire[22:0] nl_MultLoop_acc_1438_nl;
  wire[28:0] MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_896_nl;
  wire[21:0] MultLoop_acc_1439_nl;
  wire[22:0] nl_MultLoop_acc_1439_nl;
  wire[28:0] MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[10:0] AccumDotWidth_mux1h_897_nl;
  wire[10:0] AccumDotWidth_mux1h_898_nl;
  wire[21:0] AccumDotWidth_mux1h_899_nl;
  wire[21:0] MultLoop_acc_1440_nl;
  wire[22:0] nl_MultLoop_acc_1440_nl;
  wire[21:0] AccumDotWidth_mux1h_900_nl;
  wire[9:0] AccumDotWidth_acc_2436_nl;
  wire[10:0] nl_AccumDotWidth_acc_2436_nl;
  wire[9:0] AccumDotWidth_acc_2437_nl;
  wire[10:0] nl_AccumDotWidth_acc_2437_nl;
  wire[21:0] MultLoop_acc_1441_nl;
  wire[22:0] nl_MultLoop_acc_1441_nl;
  wire[21:0] AccumDotWidth_mux1h_901_nl;
  wire[21:0] MultLoop_acc_1442_nl;
  wire[22:0] nl_MultLoop_acc_1442_nl;
  wire[28:0] MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_902_nl;
  wire[21:0] MultLoop_acc_1443_nl;
  wire[22:0] nl_MultLoop_acc_1443_nl;
  wire[28:0] MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[10:0] AccumDotWidth_mux1h_903_nl;
  wire[10:0] AccumDotWidth_mux1h_904_nl;
  wire[21:0] AccumDotWidth_mux1h_905_nl;
  wire[21:0] MultLoop_acc_1444_nl;
  wire[22:0] nl_MultLoop_acc_1444_nl;
  wire[28:0] MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[10:0] AccumDotWidth_mux1h_906_nl;
  wire[0:0] AccumDotWidth_or_172_nl;
  wire[10:0] AccumDotWidth_mux1h_907_nl;
  wire[21:0] AccumDotWidth_mux1h_908_nl;
  wire[21:0] MultLoop_acc_1445_nl;
  wire[22:0] nl_MultLoop_acc_1445_nl;
  wire[28:0] MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[10:0] AccumDotWidth_mux1h_909_nl;
  wire[9:0] AccumDotWidth_acc_2438_nl;
  wire[10:0] nl_AccumDotWidth_acc_2438_nl;
  wire[9:0] AccumDotWidth_acc_2439_nl;
  wire[10:0] nl_AccumDotWidth_acc_2439_nl;
  wire[9:0] AccumDotWidth_acc_2440_nl;
  wire[10:0] nl_AccumDotWidth_acc_2440_nl;
  wire[9:0] AccumDotWidth_acc_2441_nl;
  wire[10:0] nl_AccumDotWidth_acc_2441_nl;
  wire[9:0] AccumDotWidth_acc_2442_nl;
  wire[10:0] nl_AccumDotWidth_acc_2442_nl;
  wire[10:0] AccumDotWidth_mux1h_910_nl;
  wire[21:0] AccumDotWidth_mux1h_911_nl;
  wire[21:0] MultLoop_acc_1446_nl;
  wire[22:0] nl_MultLoop_acc_1446_nl;
  wire[9:0] AccumDotWidth_mux1h_912_nl;
  wire[9:0] AccumDotWidth_acc_2443_nl;
  wire[10:0] nl_AccumDotWidth_acc_2443_nl;
  wire[9:0] AccumDotWidth_acc_2444_nl;
  wire[10:0] nl_AccumDotWidth_acc_2444_nl;
  wire[9:0] AccumDotWidth_acc_2445_nl;
  wire[10:0] nl_AccumDotWidth_acc_2445_nl;
  wire[9:0] AccumDotWidth_acc_2446_nl;
  wire[10:0] nl_AccumDotWidth_acc_2446_nl;
  wire[9:0] AccumDotWidth_acc_2447_nl;
  wire[10:0] nl_AccumDotWidth_acc_2447_nl;
  wire[9:0] AccumDotWidth_acc_2448_nl;
  wire[10:0] nl_AccumDotWidth_acc_2448_nl;
  wire[10:0] AccumDotWidth_mux1h_913_nl;
  wire[20:0] AccumDotWidth_mux1h_914_nl;
  wire[9:0] AccumDotWidth_mux1h_915_nl;
  wire[9:0] AccumDotWidth_acc_2449_nl;
  wire[10:0] nl_AccumDotWidth_acc_2449_nl;
  wire[9:0] AccumDotWidth_acc_2450_nl;
  wire[10:0] nl_AccumDotWidth_acc_2450_nl;
  wire[9:0] AccumDotWidth_acc_2451_nl;
  wire[10:0] nl_AccumDotWidth_acc_2451_nl;
  wire[9:0] AccumDotWidth_acc_2452_nl;
  wire[10:0] nl_AccumDotWidth_acc_2452_nl;
  wire[9:0] AccumDotWidth_acc_2453_nl;
  wire[10:0] nl_AccumDotWidth_acc_2453_nl;
  wire[9:0] AccumDotWidth_acc_2454_nl;
  wire[10:0] nl_AccumDotWidth_acc_2454_nl;
  wire[10:0] AccumDotWidth_mux1h_916_nl;
  wire[20:0] AccumDotWidth_mux1h_917_nl;
  wire[9:0] AccumDotWidth_mux1h_918_nl;
  wire[9:0] AccumDotWidth_acc_2455_nl;
  wire[10:0] nl_AccumDotWidth_acc_2455_nl;
  wire[9:0] AccumDotWidth_acc_2456_nl;
  wire[10:0] nl_AccumDotWidth_acc_2456_nl;
  wire[9:0] AccumDotWidth_acc_2457_nl;
  wire[10:0] nl_AccumDotWidth_acc_2457_nl;
  wire[9:0] AccumDotWidth_acc_2458_nl;
  wire[10:0] nl_AccumDotWidth_acc_2458_nl;
  wire[10:0] AccumDotWidth_mux1h_919_nl;
  wire[20:0] AccumDotWidth_mux1h_920_nl;
  wire[9:0] AccumDotWidth_mux1h_921_nl;
  wire[9:0] AccumDotWidth_acc_2459_nl;
  wire[10:0] nl_AccumDotWidth_acc_2459_nl;
  wire[9:0] AccumDotWidth_acc_2460_nl;
  wire[10:0] nl_AccumDotWidth_acc_2460_nl;
  wire[9:0] AccumDotWidth_acc_2461_nl;
  wire[10:0] nl_AccumDotWidth_acc_2461_nl;
  wire[9:0] AccumDotWidth_acc_2462_nl;
  wire[10:0] nl_AccumDotWidth_acc_2462_nl;
  wire[9:0] AccumDotWidth_acc_2463_nl;
  wire[10:0] nl_AccumDotWidth_acc_2463_nl;
  wire[10:0] AccumDotWidth_mux1h_922_nl;
  wire[20:0] AccumDotWidth_mux1h_923_nl;
  wire[21:0] AccumDotWidth_mux1h_924_nl;
  wire[21:0] AccumDotWidth_acc_2464_nl;
  wire[22:0] nl_AccumDotWidth_acc_2464_nl;
  wire[9:0] AccumDotWidth_mux1h_925_nl;
  wire[9:0] AccumDotWidth_acc_2465_nl;
  wire[10:0] nl_AccumDotWidth_acc_2465_nl;
  wire[9:0] AccumDotWidth_acc_2466_nl;
  wire[10:0] nl_AccumDotWidth_acc_2466_nl;
  wire[9:0] AccumDotWidth_acc_2467_nl;
  wire[10:0] nl_AccumDotWidth_acc_2467_nl;
  wire[10:0] AccumDotWidth_mux1h_926_nl;
  wire[20:0] AccumDotWidth_mux1h_927_nl;
  wire[9:0] AccumDotWidth_acc_2468_nl;
  wire[10:0] nl_AccumDotWidth_acc_2468_nl;
  wire[9:0] AccumDotWidth_acc_2469_nl;
  wire[10:0] nl_AccumDotWidth_acc_2469_nl;
  wire[9:0] AccumDotWidth_acc_2470_nl;
  wire[10:0] nl_AccumDotWidth_acc_2470_nl;
  wire[9:0] AccumDotWidth_acc_2471_nl;
  wire[10:0] nl_AccumDotWidth_acc_2471_nl;
  wire[20:0] AccumDotWidth_mux1h_928_nl;
  wire[21:0] AccumDotWidth_mux_96_nl;
  wire[21:0] AccumDotWidth_acc_2472_nl;
  wire[22:0] nl_AccumDotWidth_acc_2472_nl;
  wire[9:0] AccumDotWidth_mux_97_nl;
  wire[9:0] AccumDotWidth_acc_2473_nl;
  wire[10:0] nl_AccumDotWidth_acc_2473_nl;
  wire[9:0] AccumDotWidth_acc_2474_nl;
  wire[10:0] nl_AccumDotWidth_acc_2474_nl;
  wire[10:0] AccumDotWidth_mux_98_nl;
  wire[9:0] AccumDotWidth_mux1h_929_nl;
  wire[9:0] AccumDotWidth_acc_2475_nl;
  wire[10:0] nl_AccumDotWidth_acc_2475_nl;
  wire[9:0] AccumDotWidth_acc_2476_nl;
  wire[10:0] nl_AccumDotWidth_acc_2476_nl;
  wire[9:0] AccumDotWidth_acc_2477_nl;
  wire[10:0] nl_AccumDotWidth_acc_2477_nl;
  wire[9:0] AccumDotWidth_acc_2478_nl;
  wire[10:0] nl_AccumDotWidth_acc_2478_nl;
  wire[9:0] AccumDotWidth_acc_2479_nl;
  wire[10:0] nl_AccumDotWidth_acc_2479_nl;
  wire[9:0] AccumDotWidth_acc_2480_nl;
  wire[10:0] nl_AccumDotWidth_acc_2480_nl;
  wire[10:0] AccumDotWidth_mux1h_930_nl;
  wire[20:0] AccumDotWidth_mux1h_931_nl;
  wire[20:0] AccumDotWidth_mux1h_932_nl;
  wire[9:0] AccumDotWidth_acc_2481_nl;
  wire[10:0] nl_AccumDotWidth_acc_2481_nl;
  wire[9:0] AccumDotWidth_acc_2482_nl;
  wire[10:0] nl_AccumDotWidth_acc_2482_nl;
  wire[20:0] AccumDotWidth_mux1h_933_nl;
  wire[20:0] AccumDotWidth_mux1h_934_nl;
  wire[9:0] AccumDotWidth_acc_2483_nl;
  wire[10:0] nl_AccumDotWidth_acc_2483_nl;
  wire[9:0] AccumDotWidth_acc_2484_nl;
  wire[10:0] nl_AccumDotWidth_acc_2484_nl;
  wire[20:0] AccumDotWidth_mux1h_935_nl;
  wire[20:0] AccumDotWidth_mux1h_936_nl;
  wire[20:0] AccumDotWidth_mux1h_937_nl;
  wire[20:0] AccumDotWidth_mux1h_938_nl;
  wire[9:0] AccumDotWidth_acc_2485_nl;
  wire[10:0] nl_AccumDotWidth_acc_2485_nl;
  wire[20:0] AccumDotWidth_mux1h_939_nl;
  wire[20:0] AccumDotWidth_mux1h_940_nl;
  wire[9:0] AccumDotWidth_acc_2486_nl;
  wire[10:0] nl_AccumDotWidth_acc_2486_nl;
  wire[9:0] AccumDotWidth_acc_2487_nl;
  wire[10:0] nl_AccumDotWidth_acc_2487_nl;
  wire[20:0] AccumDotWidth_mux1h_941_nl;
  wire[20:0] AccumDotWidth_mux1h_942_nl;
  wire[9:0] AccumDotWidth_acc_2488_nl;
  wire[10:0] nl_AccumDotWidth_acc_2488_nl;
  wire[20:0] AccumDotWidth_mux1h_943_nl;
  wire[20:0] AccumDotWidth_mux1h_944_nl;
  wire[20:0] AccumDotWidth_mux1h_945_nl;
  wire[20:0] AccumDotWidth_mux1h_946_nl;
  wire[20:0] AccumDotWidth_mux1h_947_nl;
  wire[20:0] AccumDotWidth_mux1h_948_nl;
  wire[20:0] AccumDotWidth_mux1h_949_nl;
  wire[20:0] AccumDotWidth_mux1h_950_nl;
  wire[20:0] AccumDotWidth_mux1h_951_nl;
  wire[20:0] AccumDotWidth_mux1h_952_nl;
  wire[20:0] AccumDotWidth_mux1h_953_nl;
  wire[20:0] AccumDotWidth_mux1h_954_nl;
  wire[20:0] AccumDotWidth_mux1h_955_nl;
  wire[20:0] AccumDotWidth_mux1h_956_nl;
  wire[20:0] AccumDotWidth_mux1h_957_nl;
  wire[20:0] AccumDotWidth_mux1h_958_nl;
  wire[20:0] AccumDotWidth_mux1h_959_nl;
  wire[20:0] AccumDotWidth_mux1h_960_nl;
  wire[20:0] AccumDotWidth_mux1h_961_nl;
  wire[20:0] AccumDotWidth_mux1h_962_nl;
  wire[20:0] AccumDotWidth_mux1h_963_nl;
  wire[20:0] AccumDotWidth_mux1h_964_nl;
  wire[20:0] AccumDotWidth_mux1h_965_nl;
  wire[20:0] AccumDotWidth_mux1h_966_nl;
  wire[20:0] AccumDotWidth_mux1h_967_nl;
  wire[20:0] AccumDotWidth_mux1h_968_nl;
  wire[20:0] AccumDotWidth_mux1h_969_nl;
  wire[20:0] AccumDotWidth_mux1h_970_nl;
  wire[20:0] AccumDotWidth_mux1h_971_nl;
  wire[20:0] AccumDotWidth_mux1h_972_nl;
  wire[20:0] AccumDotWidth_mux1h_973_nl;
  wire[20:0] AccumDotWidth_mux1h_974_nl;
  wire[20:0] AccumDotWidth_mux1h_975_nl;
  wire[20:0] AccumDotWidth_mux1h_976_nl;
  wire[20:0] AccumDotWidth_mux1h_977_nl;
  wire[20:0] AccumDotWidth_mux1h_978_nl;
  wire[20:0] AccumDotWidth_mux1h_979_nl;
  wire[20:0] AccumDotWidth_mux1h_980_nl;
  wire[20:0] AccumDotWidth_mux1h_981_nl;
  wire[20:0] AccumDotWidth_mux1h_982_nl;
  wire[20:0] AccumDotWidth_mux1h_983_nl;
  wire[20:0] AccumDotWidth_mux1h_984_nl;
  wire[20:0] AccumDotWidth_mux1h_985_nl;
  wire[20:0] AccumDotWidth_mux1h_986_nl;
  wire[20:0] AccumDotWidth_mux1h_987_nl;
  wire[20:0] AccumDotWidth_mux1h_988_nl;
  wire[20:0] AccumDotWidth_mux1h_989_nl;
  wire[20:0] AccumDotWidth_mux1h_990_nl;
  wire[20:0] AccumDotWidth_mux1h_991_nl;
  wire[20:0] AccumDotWidth_mux1h_992_nl;
  wire[20:0] AccumDotWidth_mux1h_993_nl;
  wire[20:0] AccumDotWidth_mux1h_994_nl;
  wire[20:0] AccumDotWidth_mux1h_995_nl;
  wire[20:0] AccumDotWidth_mux1h_996_nl;
  wire[20:0] AccumDotWidth_mux1h_997_nl;
  wire[20:0] AccumDotWidth_mux1h_998_nl;
  wire[20:0] AccumDotWidth_mux1h_999_nl;
  wire[20:0] AccumDotWidth_mux_99_nl;
  wire[20:0] AccumDotWidth_mux_100_nl;
  wire[20:0] AccumDotWidth_mux1h_1000_nl;
  wire[20:0] AccumDotWidth_mux1h_1001_nl;
  wire[20:0] AccumDotWidth_mux1h_1002_nl;
  wire[20:0] AccumDotWidth_mux1h_1003_nl;
  wire[20:0] AccumDotWidth_mux1h_1004_nl;
  wire[20:0] AccumDotWidth_mux1h_1005_nl;
  wire[20:0] AccumDotWidth_mux1h_1006_nl;
  wire[20:0] AccumDotWidth_mux1h_1007_nl;
  wire[20:0] AccumDotWidth_mux1h_1008_nl;
  wire[20:0] AccumDotWidth_mux1h_1009_nl;
  wire[20:0] AccumDotWidth_mux1h_1010_nl;
  wire[20:0] AccumDotWidth_mux1h_1011_nl;
  wire[20:0] AccumDotWidth_mux1h_1012_nl;
  wire[20:0] AccumDotWidth_mux1h_1013_nl;
  wire[20:0] AccumDotWidth_mux1h_1014_nl;
  wire[20:0] AccumDotWidth_mux1h_1015_nl;
  wire[20:0] AccumDotWidth_mux1h_1016_nl;
  wire[20:0] AccumDotWidth_mux1h_1017_nl;
  wire[20:0] AccumDotWidth_mux1h_1018_nl;
  wire[20:0] AccumDotWidth_mux1h_1019_nl;
  wire[20:0] AccumDotWidth_mux1h_1020_nl;
  wire[20:0] AccumDotWidth_mux1h_1021_nl;
  wire[20:0] AccumDotWidth_mux1h_1022_nl;
  wire[20:0] AccumDotWidth_mux1h_1023_nl;
  wire[20:0] AccumDotWidth_mux1h_1024_nl;
  wire[20:0] AccumDotWidth_mux1h_1025_nl;
  wire[20:0] AccumDotWidth_mux1h_1026_nl;
  wire[20:0] AccumDotWidth_mux1h_1027_nl;
  wire[20:0] AccumDotWidth_mux1h_1028_nl;
  wire[20:0] AccumDotWidth_mux1h_1029_nl;
  wire[20:0] AccumDotWidth_mux1h_1030_nl;
  wire[20:0] AccumDotWidth_mux1h_1031_nl;
  wire[20:0] AccumDotWidth_mux1h_1032_nl;
  wire[20:0] AccumDotWidth_mux1h_1033_nl;
  wire[21:0] AccumDotWidth_mux1h_1034_nl;
  wire[20:0] AccumDotWidth_mux1h_1035_nl;
  wire[9:0] AccumDotWidth_acc_2489_nl;
  wire[10:0] nl_AccumDotWidth_acc_2489_nl;
  wire[20:0] AccumDotWidth_mux1h_1036_nl;
  wire[20:0] AccumDotWidth_mux1h_1037_nl;
  wire[20:0] AccumDotWidth_mux1h_1038_nl;
  wire[20:0] AccumDotWidth_mux1h_1039_nl;
  wire[20:0] AccumDotWidth_mux1h_1040_nl;
  wire[20:0] AccumDotWidth_mux1h_1041_nl;
  wire[20:0] AccumDotWidth_mux_101_nl;
  wire[20:0] AccumDotWidth_mux_102_nl;
  wire[21:0] AccumDotWidth_mux1h_1042_nl;
  wire[21:0] AccumDotWidth_acc_2490_nl;
  wire[22:0] nl_AccumDotWidth_acc_2490_nl;
  wire[20:0] AccumDotWidth_mux1h_1043_nl;
  wire[9:0] AccumDotWidth_acc_2491_nl;
  wire[10:0] nl_AccumDotWidth_acc_2491_nl;
  wire[20:0] AccumDotWidth_mux1h_1044_nl;
  wire[20:0] AccumDotWidth_mux1h_1045_nl;
  wire[20:0] AccumDotWidth_mux_103_nl;
  wire[20:0] AccumDotWidth_mux_104_nl;
  wire[20:0] AccumDotWidth_mux_105_nl;
  wire[20:0] AccumDotWidth_mux_106_nl;
  wire[20:0] AccumDotWidth_mux_107_nl;
  wire[20:0] AccumDotWidth_mux_108_nl;
  wire[20:0] AccumDotWidth_mux1h_1046_nl;
  wire[20:0] AccumDotWidth_mux1h_1047_nl;
  wire[20:0] AccumDotWidth_mux1h_1048_nl;
  wire[20:0] AccumDotWidth_mux1h_1049_nl;
  wire[20:0] AccumDotWidth_mux1h_1050_nl;
  wire[20:0] AccumDotWidth_mux1h_1051_nl;
  wire[20:0] AccumDotWidth_mux1h_1052_nl;
  wire[20:0] AccumDotWidth_mux1h_1053_nl;
  wire[20:0] AccumDotWidth_mux1h_1054_nl;
  wire[20:0] AccumDotWidth_mux1h_1055_nl;
  wire[20:0] AccumDotWidth_mux1h_1056_nl;
  wire[20:0] AccumDotWidth_mux1h_1057_nl;
  wire[20:0] AccumDotWidth_mux1h_1058_nl;
  wire[20:0] AccumDotWidth_mux1h_1059_nl;
  wire[20:0] AccumDotWidth_mux1h_1060_nl;
  wire[20:0] AccumDotWidth_mux1h_1061_nl;
  wire[20:0] AccumDotWidth_mux_109_nl;
  wire[20:0] AccumDotWidth_mux_110_nl;
  wire[20:0] AccumDotWidth_mux_111_nl;
  wire[20:0] AccumDotWidth_mux_112_nl;
  wire[20:0] AccumDotWidth_mux1h_1062_nl;
  wire[20:0] AccumDotWidth_mux1h_1063_nl;
  wire[20:0] AccumDotWidth_mux1h_1064_nl;
  wire[20:0] AccumDotWidth_mux1h_1065_nl;
  wire[20:0] AccumDotWidth_mux1h_1066_nl;
  wire[20:0] AccumDotWidth_mux1h_1067_nl;
  wire[9:0] AccumDotWidth_mux_113_nl;
  wire[9:0] AccumDotWidth_acc_2492_nl;
  wire[10:0] nl_AccumDotWidth_acc_2492_nl;
  wire[9:0] AccumDotWidth_acc_2493_nl;
  wire[10:0] nl_AccumDotWidth_acc_2493_nl;
  wire[10:0] AccumDotWidth_mux_114_nl;
  wire[9:0] AccumDotWidth_mux_115_nl;
  wire[9:0] AccumDotWidth_acc_2494_nl;
  wire[10:0] nl_AccumDotWidth_acc_2494_nl;
  wire[9:0] AccumDotWidth_acc_2495_nl;
  wire[10:0] nl_AccumDotWidth_acc_2495_nl;
  wire[10:0] AccumDotWidth_mux_116_nl;
  wire[9:0] AccumDotWidth_mux_117_nl;
  wire[9:0] AccumDotWidth_acc_2496_nl;
  wire[10:0] nl_AccumDotWidth_acc_2496_nl;
  wire[9:0] AccumDotWidth_acc_2497_nl;
  wire[10:0] nl_AccumDotWidth_acc_2497_nl;
  wire[20:0] AccumDotWidth_mux_118_nl;
  wire[9:0] AccumDotWidth_mux1h_1068_nl;
  wire[9:0] AccumDotWidth_acc_2498_nl;
  wire[10:0] nl_AccumDotWidth_acc_2498_nl;
  wire[9:0] AccumDotWidth_acc_2499_nl;
  wire[10:0] nl_AccumDotWidth_acc_2499_nl;
  wire[9:0] AccumDotWidth_acc_2500_nl;
  wire[10:0] nl_AccumDotWidth_acc_2500_nl;
  wire[10:0] AccumDotWidth_AccumDotWidth_mux_21_nl;
  wire[9:0] AccumDotWidth_mux1h_1069_nl;
  wire[9:0] AccumDotWidth_acc_2501_nl;
  wire[10:0] nl_AccumDotWidth_acc_2501_nl;
  wire[9:0] AccumDotWidth_acc_2502_nl;
  wire[10:0] nl_AccumDotWidth_acc_2502_nl;
  wire[9:0] AccumDotWidth_acc_2503_nl;
  wire[10:0] nl_AccumDotWidth_acc_2503_nl;
  wire[20:0] AccumDotWidth_mux1h_1070_nl;
  wire[20:0] AccumDotWidth_mux1h_1071_nl;
  wire[20:0] AccumDotWidth_mux1h_1072_nl;
  wire[20:0] AccumDotWidth_mux1h_1073_nl;
  wire[20:0] AccumDotWidth_mux_119_nl;
  wire[20:0] AccumDotWidth_mux_120_nl;
  wire[20:0] AccumDotWidth_mux_121_nl;
  wire[20:0] AccumDotWidth_mux_122_nl;
  wire[20:0] AccumDotWidth_mux_123_nl;
  wire[20:0] AccumDotWidth_mux_124_nl;
  wire[20:0] AccumDotWidth_mux_125_nl;
  wire[20:0] AccumDotWidth_mux_126_nl;
  wire[21:0] MultLoop_mux1h_430_nl;
  wire[21:0] MultLoop_acc_1447_nl;
  wire[22:0] nl_MultLoop_acc_1447_nl;
  wire[21:0] MultLoop_acc_1448_nl;
  wire[22:0] nl_MultLoop_acc_1448_nl;
  wire[21:0] MultLoop_acc_1449_nl;
  wire[22:0] nl_MultLoop_acc_1449_nl;
  wire[21:0] MultLoop_mux1h_431_nl;
  wire[21:0] MultLoop_acc_1450_nl;
  wire[22:0] nl_MultLoop_acc_1450_nl;
  wire[21:0] MultLoop_mux_89_nl;
  wire[21:0] MultLoop_mux_90_nl;
  wire[21:0] MultLoop_mux1h_432_nl;
  wire[21:0] MultLoop_mux1h_433_nl;
  wire[21:0] MultLoop_mux1h_434_nl;
  wire[21:0] MultLoop_mux1h_435_nl;
  wire[21:0] MultLoop_mux_91_nl;
  wire[21:0] MultLoop_mux_92_nl;
  wire[21:0] MultLoop_mux1h_436_nl;
  wire[21:0] MultLoop_mux1h_437_nl;
  wire[21:0] MultLoop_mux1h_438_nl;
  wire[21:0] MultLoop_mux1h_439_nl;
  wire[21:0] MultLoop_mux1h_440_nl;
  wire[21:0] MultLoop_mux1h_441_nl;
  wire[21:0] AccumDotWidth_mux_127_nl;
  wire[21:0] AccumDotWidth_mux_128_nl;
  wire[21:0] AccumDotWidth_mux_129_nl;
  wire[21:0] AccumDotWidth_mux_130_nl;
  wire[21:0] MultLoop_mux1h_442_nl;
  wire[21:0] MultLoop_mux1h_443_nl;
  wire[21:0] MultLoop_mux1h_444_nl;
  wire[21:0] MultLoop_mux1h_445_nl;
  wire[21:0] MultLoop_MultLoop_mux_14_nl;
  wire[21:0] MultLoop_mux1h_446_nl;
  wire[21:0] MultLoop_mux1h_447_nl;
  wire[21:0] MultLoop_mux1h_448_nl;
  wire[21:0] AccumDotWidth_mux1h_1074_nl;
  wire[21:0] AccumDotWidth_mux1h_1075_nl;
  wire[21:0] MultLoop_mux1h_449_nl;
  wire[21:0] MultLoop_mux1h_450_nl;
  wire[21:0] MultLoop_mux1h_451_nl;
  wire[21:0] MultLoop_mux1h_452_nl;
  wire[21:0] AccumDotWidth_mux1h_1076_nl;
  wire[21:0] AccumDotWidth_mux1h_1077_nl;
  wire[21:0] MultLoop_acc_1451_nl;
  wire[22:0] nl_MultLoop_acc_1451_nl;
  wire[21:0] MultLoop_acc_1452_nl;
  wire[22:0] nl_MultLoop_acc_1452_nl;
  wire[21:0] MultLoop_acc_1453_nl;
  wire[22:0] nl_MultLoop_acc_1453_nl;
  wire[21:0] AccumDotWidth_mux1h_1078_nl;
  wire[21:0] AccumDotWidth_acc_2504_nl;
  wire[22:0] nl_AccumDotWidth_acc_2504_nl;
  wire[21:0] AccumDotWidth_mux1h_1079_nl;
  wire[21:0] MultLoop_acc_1454_nl;
  wire[22:0] nl_MultLoop_acc_1454_nl;
  wire[21:0] MultLoop_acc_1455_nl;
  wire[22:0] nl_MultLoop_acc_1455_nl;
  wire[28:0] MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1456_nl;
  wire[22:0] nl_MultLoop_acc_1456_nl;
  wire[28:0] MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_453_nl;
  wire[21:0] MultLoop_mux1h_454_nl;
  wire[21:0] AccumDotWidth_mux1h_1080_nl;
  wire[21:0] AccumDotWidth_acc_2505_nl;
  wire[22:0] nl_AccumDotWidth_acc_2505_nl;
  wire[21:0] MultLoop_acc_1457_nl;
  wire[22:0] nl_MultLoop_acc_1457_nl;
  wire[21:0] MultLoop_acc_1458_nl;
  wire[22:0] nl_MultLoop_acc_1458_nl;
  wire[28:0] MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1459_nl;
  wire[22:0] nl_MultLoop_acc_1459_nl;
  wire[28:0] MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1081_nl;
  wire[21:0] MultLoop_mux1h_455_nl;
  wire[21:0] MultLoop_acc_1460_nl;
  wire[22:0] nl_MultLoop_acc_1460_nl;
  wire[21:0] MultLoop_acc_1461_nl;
  wire[23:0] nl_MultLoop_acc_1461_nl;
  wire[21:0] MultLoop_acc_1462_nl;
  wire[22:0] nl_MultLoop_acc_1462_nl;
  wire[21:0] MultLoop_acc_1465_nl;
  wire[22:0] nl_MultLoop_acc_1465_nl;
  wire[21:0] MultLoop_acc_1466_nl;
  wire[22:0] nl_MultLoop_acc_1466_nl;
  wire[21:0] MultLoop_mux1h_456_nl;
  wire[21:0] MultLoop_acc_1467_nl;
  wire[22:0] nl_MultLoop_acc_1467_nl;
  wire[21:0] AccumDotWidth_mux1h_1082_nl;
  wire[21:0] AccumDotWidth_acc_2506_nl;
  wire[22:0] nl_AccumDotWidth_acc_2506_nl;
  wire[21:0] MultLoop_acc_1468_nl;
  wire[22:0] nl_MultLoop_acc_1468_nl;
  wire[21:0] AccumDotWidth_mux1h_1083_nl;
  wire[21:0] AccumDotWidth_acc_2507_nl;
  wire[22:0] nl_AccumDotWidth_acc_2507_nl;
  wire[21:0] MultLoop_mux1h_457_nl;
  wire[21:0] MultLoop_mux1h_458_nl;
  wire[21:0] MultLoop_mux_93_nl;
  wire[21:0] MultLoop_acc_1469_nl;
  wire[22:0] nl_MultLoop_acc_1469_nl;
  wire[21:0] MultLoop_acc_1470_nl;
  wire[22:0] nl_MultLoop_acc_1470_nl;
  wire[21:0] MultLoop_acc_1471_nl;
  wire[22:0] nl_MultLoop_acc_1471_nl;
  wire[21:0] MultLoop_mux_94_nl;
  wire[21:0] AccumDotWidth_mux1h_1084_nl;
  wire[21:0] AccumDotWidth_acc_2508_nl;
  wire[22:0] nl_AccumDotWidth_acc_2508_nl;
  wire[21:0] AccumDotWidth_mux1h_1085_nl;
  wire[21:0] AccumDotWidth_acc_2509_nl;
  wire[22:0] nl_AccumDotWidth_acc_2509_nl;
  wire[21:0] AccumDotWidth_mux_131_nl;
  wire[21:0] AccumDotWidth_mux_132_nl;
  wire[21:0] AccumDotWidth_mux1h_1086_nl;
  wire[21:0] AccumDotWidth_acc_2510_nl;
  wire[22:0] nl_AccumDotWidth_acc_2510_nl;
  wire[21:0] AccumDotWidth_mux1h_1087_nl;
  wire[21:0] MultLoop_acc_1472_nl;
  wire[22:0] nl_MultLoop_acc_1472_nl;
  wire[21:0] AccumDotWidth_mux1h_1088_nl;
  wire[21:0] MultLoop_acc_1473_nl;
  wire[22:0] nl_MultLoop_acc_1473_nl;
  wire[21:0] MultLoop_acc_1474_nl;
  wire[22:0] nl_MultLoop_acc_1474_nl;
  wire[21:0] AccumDotWidth_mux1h_1089_nl;
  wire[21:0] MultLoop_acc_1475_nl;
  wire[22:0] nl_MultLoop_acc_1475_nl;
  wire[21:0] MultLoop_acc_1476_nl;
  wire[22:0] nl_MultLoop_acc_1476_nl;
  wire[21:0] MultLoop_acc_1477_nl;
  wire[22:0] nl_MultLoop_acc_1477_nl;
  wire[21:0] MultLoop_mux1h_459_nl;
  wire[21:0] MultLoop_mux1h_460_nl;
  wire[21:0] AccumDotWidth_mux1h_1090_nl;
  wire[21:0] AccumDotWidth_mux1h_1091_nl;
  wire[21:0] AccumDotWidth_mux1h_1092_nl;
  wire[21:0] AccumDotWidth_acc_2511_nl;
  wire[22:0] nl_AccumDotWidth_acc_2511_nl;
  wire[21:0] AccumDotWidth_mux1h_1093_nl;
  wire[21:0] MultLoop_mux1h_461_nl;
  wire[21:0] MultLoop_mux1h_462_nl;
  wire[21:0] AccumDotWidth_mux1h_1094_nl;
  wire[21:0] MultLoop_acc_1478_nl;
  wire[23:0] nl_MultLoop_acc_1478_nl;
  wire[21:0] MultLoop_acc_1480_nl;
  wire[22:0] nl_MultLoop_acc_1480_nl;
  wire[21:0] MultLoop_acc_1481_nl;
  wire[22:0] nl_MultLoop_acc_1481_nl;
  wire[21:0] MultLoop_acc_1483_nl;
  wire[22:0] nl_MultLoop_acc_1483_nl;
  wire[21:0] MultLoop_acc_1484_nl;
  wire[22:0] nl_MultLoop_acc_1484_nl;
  wire[21:0] AccumDotWidth_mux1h_1095_nl;
  wire[21:0] MultLoop_acc_1485_nl;
  wire[22:0] nl_MultLoop_acc_1485_nl;
  wire[21:0] MultLoop_acc_1486_nl;
  wire[22:0] nl_MultLoop_acc_1486_nl;
  wire[21:0] MultLoop_acc_1487_nl;
  wire[22:0] nl_MultLoop_acc_1487_nl;
  wire[21:0] AccumDotWidth_mux1h_1096_nl;
  wire[21:0] AccumDotWidth_mux1h_1097_nl;
  wire[21:0] AccumDotWidth_mux1h_1098_nl;
  wire[21:0] AccumDotWidth_mux1h_1099_nl;
  wire[21:0] AccumDotWidth_mux1h_1100_nl;
  wire[21:0] MultLoop_acc_1488_nl;
  wire[23:0] nl_MultLoop_acc_1488_nl;
  wire[21:0] MultLoop_acc_1490_nl;
  wire[22:0] nl_MultLoop_acc_1490_nl;
  wire[21:0] MultLoop_acc_1491_nl;
  wire[22:0] nl_MultLoop_acc_1491_nl;
  wire[21:0] MultLoop_acc_1493_nl;
  wire[22:0] nl_MultLoop_acc_1493_nl;
  wire[21:0] MultLoop_acc_1494_nl;
  wire[22:0] nl_MultLoop_acc_1494_nl;
  wire[21:0] AccumDotWidth_mux1h_1101_nl;
  wire[21:0] MultLoop_acc_1495_nl;
  wire[23:0] nl_MultLoop_acc_1495_nl;
  wire[21:0] MultLoop_acc_1497_nl;
  wire[22:0] nl_MultLoop_acc_1497_nl;
  wire[21:0] MultLoop_acc_1498_nl;
  wire[22:0] nl_MultLoop_acc_1498_nl;
  wire[21:0] MultLoop_acc_1500_nl;
  wire[22:0] nl_MultLoop_acc_1500_nl;
  wire[21:0] MultLoop_acc_1501_nl;
  wire[22:0] nl_MultLoop_acc_1501_nl;
  wire[21:0] AccumDotWidth_mux1h_1102_nl;
  wire[21:0] MultLoop_acc_1502_nl;
  wire[22:0] nl_MultLoop_acc_1502_nl;
  wire[21:0] AccumDotWidth_mux1h_1103_nl;
  wire[21:0] MultLoop_acc_1503_nl;
  wire[22:0] nl_MultLoop_acc_1503_nl;
  wire[21:0] MultLoop_acc_1504_nl;
  wire[22:0] nl_MultLoop_acc_1504_nl;
  wire[21:0] MultLoop_acc_1505_nl;
  wire[22:0] nl_MultLoop_acc_1505_nl;
  wire[21:0] AccumDotWidth_mux1h_1104_nl;
  wire[21:0] MultLoop_acc_1506_nl;
  wire[22:0] nl_MultLoop_acc_1506_nl;
  wire[21:0] MultLoop_acc_1507_nl;
  wire[22:0] nl_MultLoop_acc_1507_nl;
  wire[21:0] MultLoop_acc_1508_nl;
  wire[22:0] nl_MultLoop_acc_1508_nl;
  wire[21:0] AccumDotWidth_mux1h_1105_nl;
  wire[21:0] AccumDotWidth_mux1h_1106_nl;
  wire[21:0] AccumDotWidth_mux1h_1107_nl;
  wire[21:0] AccumDotWidth_mux1h_1108_nl;
  wire[21:0] AccumDotWidth_mux1h_1109_nl;
  wire[21:0] MultLoop_acc_1509_nl;
  wire[22:0] nl_MultLoop_acc_1509_nl;
  wire[21:0] MultLoop_mux1h_463_nl;
  wire[21:0] MultLoop_mux1h_464_nl;
  wire[21:0] MultLoop_mux1h_465_nl;
  wire[21:0] MultLoop_mux1h_466_nl;
  wire[21:0] MultLoop_mux1h_467_nl;
  wire[21:0] MultLoop_mux1h_468_nl;
  wire[21:0] AccumDotWidth_mux_133_nl;
  wire[21:0] MultLoop_acc_1510_nl;
  wire[22:0] nl_MultLoop_acc_1510_nl;
  wire[21:0] AccumDotWidth_mux_134_nl;
  wire[21:0] MultLoop_acc_1511_nl;
  wire[22:0] nl_MultLoop_acc_1511_nl;
  wire[21:0] AccumDotWidth_mux1h_1110_nl;
  wire[21:0] AccumDotWidth_mux1h_1111_nl;
  wire[21:0] MultLoop_acc_1512_nl;
  wire[22:0] nl_MultLoop_acc_1512_nl;
  wire[21:0] MultLoop_acc_1513_nl;
  wire[22:0] nl_MultLoop_acc_1513_nl;
  wire[21:0] MultLoop_acc_1514_nl;
  wire[22:0] nl_MultLoop_acc_1514_nl;
  wire[21:0] MultLoop_acc_1515_nl;
  wire[22:0] nl_MultLoop_acc_1515_nl;
  wire[21:0] MultLoop_mux1h_469_nl;
  wire[21:0] MultLoop_acc_1516_nl;
  wire[22:0] nl_MultLoop_acc_1516_nl;
  wire[21:0] MultLoop_mux1h_470_nl;
  wire[21:0] MultLoop_acc_1517_nl;
  wire[22:0] nl_MultLoop_acc_1517_nl;
  wire[21:0] MultLoop_acc_1518_nl;
  wire[22:0] nl_MultLoop_acc_1518_nl;
  wire[21:0] MultLoop_acc_1519_nl;
  wire[22:0] nl_MultLoop_acc_1519_nl;
  wire[21:0] MultLoop_acc_1520_nl;
  wire[22:0] nl_MultLoop_acc_1520_nl;
  wire[21:0] AccumDotWidth_mux1h_1112_nl;
  wire[21:0] AccumDotWidth_acc_2512_nl;
  wire[22:0] nl_AccumDotWidth_acc_2512_nl;
  wire[21:0] AccumDotWidth_mux1h_1113_nl;
  wire[21:0] AccumDotWidth_mux1h_1114_nl;
  wire[21:0] AccumDotWidth_acc_2513_nl;
  wire[22:0] nl_AccumDotWidth_acc_2513_nl;
  wire[21:0] AccumDotWidth_mux1h_1115_nl;
  wire[21:0] AccumDotWidth_acc_2514_nl;
  wire[22:0] nl_AccumDotWidth_acc_2514_nl;
  wire[21:0] MultLoop_mux1h_471_nl;
  wire[21:0] MultLoop_mux1h_472_nl;
  wire[21:0] MultLoop_acc_1521_nl;
  wire[22:0] nl_MultLoop_acc_1521_nl;
  wire[21:0] AccumDotWidth_mux_135_nl;
  wire[21:0] AccumDotWidth_mux_136_nl;
  wire[21:0] AccumDotWidth_mux_137_nl;
  wire[21:0] AccumDotWidth_mux_138_nl;
  wire[21:0] MultLoop_mux1h_473_nl;
  wire[21:0] AccumDotWidth_acc_2515_nl;
  wire[22:0] nl_AccumDotWidth_acc_2515_nl;
  wire[21:0] MultLoop_mux1h_474_nl;
  wire[21:0] AccumDotWidth_mux1h_1116_nl;
  wire[21:0] AccumDotWidth_acc_2516_nl;
  wire[22:0] nl_AccumDotWidth_acc_2516_nl;
  wire[21:0] AccumDotWidth_mux1h_1117_nl;
  wire[21:0] AccumDotWidth_acc_2517_nl;
  wire[22:0] nl_AccumDotWidth_acc_2517_nl;
  wire[21:0] AccumDotWidth_acc_2518_nl;
  wire[22:0] nl_AccumDotWidth_acc_2518_nl;
  wire[21:0] MultLoop_mux1h_475_nl;
  wire[21:0] AccumDotWidth_acc_2519_nl;
  wire[22:0] nl_AccumDotWidth_acc_2519_nl;
  wire[21:0] AccumDotWidth_acc_2520_nl;
  wire[22:0] nl_AccumDotWidth_acc_2520_nl;
  wire[21:0] MultLoop_mux1h_476_nl;
  wire[21:0] AccumDotWidth_acc_2521_nl;
  wire[22:0] nl_AccumDotWidth_acc_2521_nl;
  wire[21:0] MultLoop_mux1h_477_nl;
  wire[21:0] AccumDotWidth_acc_2522_nl;
  wire[22:0] nl_AccumDotWidth_acc_2522_nl;
  wire[21:0] MultLoop_mux1h_478_nl;
  wire[21:0] AccumDotWidth_acc_2523_nl;
  wire[22:0] nl_AccumDotWidth_acc_2523_nl;
  wire[21:0] AccumDotWidth_mux1h_1118_nl;
  wire[21:0] AccumDotWidth_mux1h_1119_nl;
  wire[21:0] AccumDotWidth_mux1h_1120_nl;
  wire[21:0] AccumDotWidth_acc_2524_nl;
  wire[22:0] nl_AccumDotWidth_acc_2524_nl;
  wire[21:0] AccumDotWidth_acc_2525_nl;
  wire[22:0] nl_AccumDotWidth_acc_2525_nl;
  wire[21:0] AccumDotWidth_acc_2526_nl;
  wire[22:0] nl_AccumDotWidth_acc_2526_nl;
  wire[21:0] AccumDotWidth_mux1h_1121_nl;
  wire[21:0] AccumDotWidth_acc_2527_nl;
  wire[22:0] nl_AccumDotWidth_acc_2527_nl;
  wire[21:0] AccumDotWidth_acc_2528_nl;
  wire[22:0] nl_AccumDotWidth_acc_2528_nl;
  wire[9:0] AccumDotWidth_acc_2529_nl;
  wire[10:0] nl_AccumDotWidth_acc_2529_nl;
  wire[21:0] AccumDotWidth_acc_2530_nl;
  wire[22:0] nl_AccumDotWidth_acc_2530_nl;
  wire[21:0] AccumDotWidth_acc_2531_nl;
  wire[22:0] nl_AccumDotWidth_acc_2531_nl;
  wire[21:0] MultLoop_mux1h_479_nl;
  wire[21:0] AccumDotWidth_acc_2532_nl;
  wire[22:0] nl_AccumDotWidth_acc_2532_nl;
  wire[21:0] AccumDotWidth_acc_2533_nl;
  wire[22:0] nl_AccumDotWidth_acc_2533_nl;
  wire[21:0] AccumDotWidth_acc_2534_nl;
  wire[22:0] nl_AccumDotWidth_acc_2534_nl;
  wire[21:0] MultLoop_mux1h_480_nl;
  wire[21:0] AccumDotWidth_acc_2535_nl;
  wire[22:0] nl_AccumDotWidth_acc_2535_nl;
  wire[9:0] AccumDotWidth_acc_2536_nl;
  wire[10:0] nl_AccumDotWidth_acc_2536_nl;
  wire[21:0] AccumDotWidth_acc_2537_nl;
  wire[22:0] nl_AccumDotWidth_acc_2537_nl;
  wire[21:0] AccumDotWidth_acc_2538_nl;
  wire[22:0] nl_AccumDotWidth_acc_2538_nl;
  wire[21:0] AccumDotWidth_acc_2539_nl;
  wire[22:0] nl_AccumDotWidth_acc_2539_nl;
  wire[21:0] MultLoop_mux1h_481_nl;
  wire[21:0] MultLoop_mux1h_482_nl;
  wire[21:0] MultLoop_mux_95_nl;
  wire[21:0] MultLoop_acc_1522_nl;
  wire[22:0] nl_MultLoop_acc_1522_nl;
  wire[21:0] MultLoop_mux_96_nl;
  wire[21:0] MultLoop_acc_1523_nl;
  wire[22:0] nl_MultLoop_acc_1523_nl;
  wire[21:0] MultLoop_mux1h_483_nl;
  wire[21:0] MultLoop_mux1h_484_nl;
  wire[21:0] MultLoop_mux1h_485_nl;
  wire[21:0] MultLoop_mux1h_486_nl;
  wire[21:0] MultLoop_mux1h_487_nl;
  wire[21:0] MultLoop_mux1h_488_nl;
  wire[21:0] AccumDotWidth_mux1h_1122_nl;
  wire[21:0] AccumDotWidth_mux1h_1123_nl;
  wire[21:0] AccumDotWidth_acc_2540_nl;
  wire[22:0] nl_AccumDotWidth_acc_2540_nl;
  wire[9:0] AccumDotWidth_acc_2541_nl;
  wire[10:0] nl_AccumDotWidth_acc_2541_nl;
  wire[21:0] MultLoop_mux1h_489_nl;
  wire[21:0] MultLoop_mux1h_490_nl;
  wire[21:0] MultLoop_mux1h_491_nl;
  wire[21:0] MultLoop_mux1h_492_nl;
  wire[21:0] AccumDotWidth_mux1h_1124_nl;
  wire[21:0] AccumDotWidth_acc_2542_nl;
  wire[22:0] nl_AccumDotWidth_acc_2542_nl;
  wire[21:0] AccumDotWidth_acc_2543_nl;
  wire[22:0] nl_AccumDotWidth_acc_2543_nl;
  wire[21:0] AccumDotWidth_acc_2544_nl;
  wire[22:0] nl_AccumDotWidth_acc_2544_nl;
  wire[21:0] AccumDotWidth_acc_2545_nl;
  wire[22:0] nl_AccumDotWidth_acc_2545_nl;
  wire[21:0] AccumDotWidth_mux1h_1125_nl;
  wire[21:0] AccumDotWidth_acc_2546_nl;
  wire[22:0] nl_AccumDotWidth_acc_2546_nl;
  wire[21:0] AccumDotWidth_acc_2547_nl;
  wire[22:0] nl_AccumDotWidth_acc_2547_nl;
  wire[21:0] AccumDotWidth_acc_2548_nl;
  wire[22:0] nl_AccumDotWidth_acc_2548_nl;
  wire[21:0] AccumDotWidth_acc_2549_nl;
  wire[22:0] nl_AccumDotWidth_acc_2549_nl;
  wire[21:0] MultLoop_mux1h_493_nl;
  wire[28:0] MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_494_nl;
  wire[28:0] MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux1h_495_nl;
  wire[21:0] MultLoop_mux1h_496_nl;
  wire[21:0] MultLoop_mux1h_497_nl;
  wire[21:0] MultLoop_mux1h_498_nl;
  wire[21:0] MultLoop_mux1h_499_nl;
  wire[0:0] MultLoop_or_107_nl;
  wire[21:0] MultLoop_mux1h_500_nl;
  wire[21:0] AccumDotWidth_mux1h_1126_nl;
  wire[21:0] AccumDotWidth_mux1h_1127_nl;
  wire[21:0] MultLoop_acc_1524_nl;
  wire[22:0] nl_MultLoop_acc_1524_nl;
  wire[21:0] AccumDotWidth_mux1h_1128_nl;
  wire[21:0] AccumDotWidth_mux1h_1129_nl;
  wire[21:0] MultLoop_acc_1525_nl;
  wire[23:0] nl_MultLoop_acc_1525_nl;
  wire[21:0] MultLoop_acc_1527_nl;
  wire[22:0] nl_MultLoop_acc_1527_nl;
  wire[21:0] MultLoop_acc_1528_nl;
  wire[22:0] nl_MultLoop_acc_1528_nl;
  wire[21:0] MultLoop_acc_1530_nl;
  wire[22:0] nl_MultLoop_acc_1530_nl;
  wire[21:0] MultLoop_acc_1531_nl;
  wire[22:0] nl_MultLoop_acc_1531_nl;
  wire[21:0] AccumDotWidth_mux1h_1130_nl;
  wire[21:0] AccumDotWidth_mux1h_1131_nl;
  wire[21:0] MultLoop_acc_1532_nl;
  wire[22:0] nl_MultLoop_acc_1532_nl;
  wire[21:0] AccumDotWidth_mux1h_1132_nl;
  wire[21:0] MultLoop_acc_1533_nl;
  wire[22:0] nl_MultLoop_acc_1533_nl;
  wire[21:0] AccumDotWidth_mux1h_1133_nl;
  wire[21:0] MultLoop_acc_1534_nl;
  wire[22:0] nl_MultLoop_acc_1534_nl;
  wire[21:0] AccumDotWidth_mux1h_1134_nl;
  wire[21:0] MultLoop_acc_1535_nl;
  wire[22:0] nl_MultLoop_acc_1535_nl;
  wire[21:0] AccumDotWidth_mux1h_1135_nl;
  wire[21:0] MultLoop_acc_1536_nl;
  wire[22:0] nl_MultLoop_acc_1536_nl;
  wire[21:0] AccumDotWidth_mux_139_nl;
  wire[21:0] AccumDotWidth_mux_140_nl;
  wire[21:0] AccumDotWidth_mux1h_1136_nl;
  wire[21:0] AccumDotWidth_mux1h_1137_nl;
  wire[21:0] AccumDotWidth_mux_141_nl;
  wire[21:0] MultLoop_acc_1537_nl;
  wire[22:0] nl_MultLoop_acc_1537_nl;
  wire[21:0] AccumDotWidth_mux_142_nl;
  wire[21:0] MultLoop_acc_1538_nl;
  wire[22:0] nl_MultLoop_acc_1538_nl;
  wire[21:0] AccumDotWidth_mux1h_1138_nl;
  wire[21:0] MultLoop_acc_1539_nl;
  wire[22:0] nl_MultLoop_acc_1539_nl;
  wire[21:0] AccumDotWidth_mux1h_1139_nl;
  wire[21:0] MultLoop_acc_1540_nl;
  wire[22:0] nl_MultLoop_acc_1540_nl;
  wire[21:0] AccumDotWidth_mux1h_1140_nl;
  wire[21:0] MultLoop_acc_1541_nl;
  wire[22:0] nl_MultLoop_acc_1541_nl;
  wire[21:0] AccumDotWidth_mux1h_1141_nl;
  wire[21:0] MultLoop_acc_1542_nl;
  wire[22:0] nl_MultLoop_acc_1542_nl;
  wire[21:0] AccumDotWidth_mux1h_1142_nl;
  wire[21:0] AccumDotWidth_acc_2550_nl;
  wire[22:0] nl_AccumDotWidth_acc_2550_nl;
  wire[21:0] AccumDotWidth_mux1h_1143_nl;
  wire[21:0] MultLoop_acc_1543_nl;
  wire[22:0] nl_MultLoop_acc_1543_nl;
  wire[21:0] AccumDotWidth_mux1h_1144_nl;
  wire[21:0] AccumDotWidth_mux1h_1145_nl;
  wire[21:0] MultLoop_acc_1544_nl;
  wire[22:0] nl_MultLoop_acc_1544_nl;
  wire[21:0] AccumDotWidth_mux1h_1146_nl;
  wire[21:0] AccumDotWidth_acc_2551_nl;
  wire[22:0] nl_AccumDotWidth_acc_2551_nl;
  wire[21:0] MultLoop_acc_1545_nl;
  wire[22:0] nl_MultLoop_acc_1545_nl;
  wire[21:0] AccumDotWidth_mux1h_1147_nl;
  wire[21:0] AccumDotWidth_acc_2552_nl;
  wire[22:0] nl_AccumDotWidth_acc_2552_nl;
  wire[21:0] MultLoop_acc_1546_nl;
  wire[22:0] nl_MultLoop_acc_1546_nl;
  wire[21:0] AccumDotWidth_mux1h_1148_nl;
  wire[21:0] AccumDotWidth_mux1h_1149_nl;
  wire[21:0] AccumDotWidth_mux1h_1150_nl;
  wire[21:0] AccumDotWidth_mux1h_1151_nl;
  wire[21:0] AccumDotWidth_mux1h_1152_nl;
  wire[21:0] AccumDotWidth_mux1h_1153_nl;
  wire[21:0] AccumDotWidth_mux1h_1154_nl;
  wire[21:0] AccumDotWidth_mux1h_1155_nl;
  wire[21:0] AccumDotWidth_mux1h_1156_nl;
  wire[21:0] AccumDotWidth_acc_2553_nl;
  wire[22:0] nl_AccumDotWidth_acc_2553_nl;
  wire[21:0] AccumDotWidth_acc_2554_nl;
  wire[22:0] nl_AccumDotWidth_acc_2554_nl;
  wire[21:0] AccumDotWidth_acc_2555_nl;
  wire[22:0] nl_AccumDotWidth_acc_2555_nl;
  wire[21:0] AccumDotWidth_acc_2556_nl;
  wire[22:0] nl_AccumDotWidth_acc_2556_nl;
  wire[21:0] AccumDotWidth_acc_2557_nl;
  wire[22:0] nl_AccumDotWidth_acc_2557_nl;
  wire[21:0] AccumDotWidth_acc_2558_nl;
  wire[22:0] nl_AccumDotWidth_acc_2558_nl;
  wire[21:0] AccumDotWidth_acc_2559_nl;
  wire[22:0] nl_AccumDotWidth_acc_2559_nl;
  wire[21:0] AccumDotWidth_mux1h_1157_nl;
  wire[21:0] AccumDotWidth_acc_2560_nl;
  wire[22:0] nl_AccumDotWidth_acc_2560_nl;
  wire[21:0] AccumDotWidth_acc_2561_nl;
  wire[22:0] nl_AccumDotWidth_acc_2561_nl;
  wire[21:0] AccumDotWidth_acc_2562_nl;
  wire[22:0] nl_AccumDotWidth_acc_2562_nl;
  wire[21:0] AccumDotWidth_acc_2563_nl;
  wire[22:0] nl_AccumDotWidth_acc_2563_nl;
  wire[21:0] AccumDotWidth_acc_2564_nl;
  wire[22:0] nl_AccumDotWidth_acc_2564_nl;
  wire[21:0] AccumDotWidth_acc_2565_nl;
  wire[22:0] nl_AccumDotWidth_acc_2565_nl;
  wire[21:0] AccumDotWidth_acc_2566_nl;
  wire[22:0] nl_AccumDotWidth_acc_2566_nl;
  wire[21:0] AccumDotWidth_mux1h_1158_nl;
  wire[21:0] AccumDotWidth_mux1h_1159_nl;
  wire[21:0] AccumDotWidth_mux1h_1160_nl;
  wire[21:0] AccumDotWidth_acc_2567_nl;
  wire[23:0] nl_AccumDotWidth_acc_2567_nl;
  wire[21:0] AccumDotWidth_mux1h_1161_nl;
  wire[21:0] AccumDotWidth_acc_2570_nl;
  wire[23:0] nl_AccumDotWidth_acc_2570_nl;
  wire[21:0] AccumDotWidth_mux1h_1162_nl;
  wire[21:0] AccumDotWidth_mux1h_1163_nl;
  wire[21:0] AccumDotWidth_mux1h_1164_nl;
  wire[21:0] AccumDotWidth_mux1h_1165_nl;
  wire[21:0] MultLoop_acc_1547_nl;
  wire[22:0] nl_MultLoop_acc_1547_nl;
  wire[21:0] AccumDotWidth_mux1h_1166_nl;
  wire[21:0] AccumDotWidth_acc_2573_nl;
  wire[22:0] nl_AccumDotWidth_acc_2573_nl;
  wire[21:0] AccumDotWidth_mux1h_1167_nl;
  wire[21:0] AccumDotWidth_mux1h_1168_nl;
  wire[21:0] AccumDotWidth_acc_2574_nl;
  wire[22:0] nl_AccumDotWidth_acc_2574_nl;
  wire[21:0] AccumDotWidth_mux1h_1169_nl;
  wire[21:0] AccumDotWidth_acc_2575_nl;
  wire[22:0] nl_AccumDotWidth_acc_2575_nl;
  wire[9:0] AccumDotWidth_acc_2576_nl;
  wire[10:0] nl_AccumDotWidth_acc_2576_nl;
  wire[21:0] AccumDotWidth_mux1h_1170_nl;
  wire[21:0] AccumDotWidth_mux1h_1171_nl;
  wire[21:0] AccumDotWidth_mux1h_1172_nl;
  wire[21:0] AccumDotWidth_mux1h_1173_nl;
  wire[21:0] AccumDotWidth_mux1h_1174_nl;
  wire[21:0] AccumDotWidth_mux1h_1175_nl;
  wire[21:0] AccumDotWidth_mux1h_1176_nl;
  wire[21:0] AccumDotWidth_acc_2577_nl;
  wire[22:0] nl_AccumDotWidth_acc_2577_nl;
  wire[21:0] AccumDotWidth_mux1h_1177_nl;
  wire[21:0] AccumDotWidth_mux1h_1178_nl;
  wire[21:0] AccumDotWidth_mux1h_1179_nl;
  wire[21:0] AccumDotWidth_mux1h_1180_nl;
  wire[21:0] AccumDotWidth_mux1h_1181_nl;
  wire[21:0] MultLoop_acc_1548_nl;
  wire[23:0] nl_MultLoop_acc_1548_nl;
  wire[21:0] MultLoop_acc_1550_nl;
  wire[22:0] nl_MultLoop_acc_1550_nl;
  wire[21:0] MultLoop_acc_1551_nl;
  wire[22:0] nl_MultLoop_acc_1551_nl;
  wire[21:0] MultLoop_acc_1553_nl;
  wire[22:0] nl_MultLoop_acc_1553_nl;
  wire[21:0] MultLoop_acc_1554_nl;
  wire[22:0] nl_MultLoop_acc_1554_nl;
  wire[21:0] AccumDotWidth_mux1h_1182_nl;
  wire[21:0] AccumDotWidth_mux1h_1183_nl;
  wire[21:0] AccumDotWidth_mux1h_1184_nl;
  wire[21:0] MultLoop_acc_1555_nl;
  wire[22:0] nl_MultLoop_acc_1555_nl;
  wire[21:0] MultLoop_acc_1556_nl;
  wire[22:0] nl_MultLoop_acc_1556_nl;
  wire[21:0] MultLoop_acc_1557_nl;
  wire[22:0] nl_MultLoop_acc_1557_nl;
  wire[21:0] MultLoop_acc_1558_nl;
  wire[22:0] nl_MultLoop_acc_1558_nl;
  wire[21:0] AccumDotWidth_mux1h_1185_nl;
  wire[21:0] MultLoop_acc_1559_nl;
  wire[23:0] nl_MultLoop_acc_1559_nl;
  wire[21:0] MultLoop_acc_1561_nl;
  wire[22:0] nl_MultLoop_acc_1561_nl;
  wire[21:0] MultLoop_acc_1562_nl;
  wire[22:0] nl_MultLoop_acc_1562_nl;
  wire[21:0] MultLoop_acc_1564_nl;
  wire[22:0] nl_MultLoop_acc_1564_nl;
  wire[21:0] MultLoop_acc_1565_nl;
  wire[22:0] nl_MultLoop_acc_1565_nl;
  wire[21:0] AccumDotWidth_mux1h_1186_nl;
  wire[21:0] AccumDotWidth_mux1h_1187_nl;
  wire[21:0] AccumDotWidth_mux1h_1188_nl;
  wire[21:0] MultLoop_acc_1566_nl;
  wire[23:0] nl_MultLoop_acc_1566_nl;
  wire[21:0] MultLoop_acc_1568_nl;
  wire[22:0] nl_MultLoop_acc_1568_nl;
  wire[21:0] MultLoop_acc_1569_nl;
  wire[22:0] nl_MultLoop_acc_1569_nl;
  wire[21:0] MultLoop_acc_1571_nl;
  wire[22:0] nl_MultLoop_acc_1571_nl;
  wire[28:0] MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1572_nl;
  wire[22:0] nl_MultLoop_acc_1572_nl;
  wire[28:0] MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1189_nl;
  wire[21:0] MultLoop_acc_1573_nl;
  wire[23:0] nl_MultLoop_acc_1573_nl;
  wire[21:0] MultLoop_acc_1575_nl;
  wire[22:0] nl_MultLoop_acc_1575_nl;
  wire[28:0] MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1576_nl;
  wire[22:0] nl_MultLoop_acc_1576_nl;
  wire[28:0] MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1578_nl;
  wire[22:0] nl_MultLoop_acc_1578_nl;
  wire[28:0] MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1579_nl;
  wire[22:0] nl_MultLoop_acc_1579_nl;
  wire[28:0] MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1190_nl;
  wire[21:0] AccumDotWidth_acc_2578_nl;
  wire[23:0] nl_AccumDotWidth_acc_2578_nl;
  wire[21:0] AccumDotWidth_mux1h_1191_nl;
  wire[21:0] AccumDotWidth_mux1h_1192_nl;
  wire[21:0] MultLoop_acc_1580_nl;
  wire[23:0] nl_MultLoop_acc_1580_nl;
  wire[21:0] MultLoop_acc_1582_nl;
  wire[22:0] nl_MultLoop_acc_1582_nl;
  wire[28:0] MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1583_nl;
  wire[22:0] nl_MultLoop_acc_1583_nl;
  wire[28:0] MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1585_nl;
  wire[22:0] nl_MultLoop_acc_1585_nl;
  wire[28:0] MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1586_nl;
  wire[22:0] nl_MultLoop_acc_1586_nl;
  wire[28:0] MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1193_nl;
  wire[21:0] MultLoop_acc_1587_nl;
  wire[23:0] nl_MultLoop_acc_1587_nl;
  wire[21:0] MultLoop_acc_1589_nl;
  wire[22:0] nl_MultLoop_acc_1589_nl;
  wire[28:0] MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1590_nl;
  wire[22:0] nl_MultLoop_acc_1590_nl;
  wire[28:0] MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1592_nl;
  wire[22:0] nl_MultLoop_acc_1592_nl;
  wire[28:0] MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1593_nl;
  wire[22:0] nl_MultLoop_acc_1593_nl;
  wire[21:0] MultLoop_mux1h_501_nl;
  wire[21:0] AccumDotWidth_acc_2581_nl;
  wire[22:0] nl_AccumDotWidth_acc_2581_nl;
  wire[21:0] MultLoop_mux1h_502_nl;
  wire[21:0] AccumDotWidth_acc_2582_nl;
  wire[22:0] nl_AccumDotWidth_acc_2582_nl;
  wire[21:0] AccumDotWidth_acc_2583_nl;
  wire[22:0] nl_AccumDotWidth_acc_2583_nl;
  wire[21:0] AccumDotWidth_mux1h_1194_nl;
  wire[21:0] AccumDotWidth_acc_2584_nl;
  wire[22:0] nl_AccumDotWidth_acc_2584_nl;
  wire[21:0] AccumDotWidth_mux1h_1195_nl;
  wire[21:0] AccumDotWidth_acc_2585_nl;
  wire[22:0] nl_AccumDotWidth_acc_2585_nl;
  wire[21:0] AccumDotWidth_acc_2586_nl;
  wire[22:0] nl_AccumDotWidth_acc_2586_nl;
  wire[21:0] AccumDotWidth_mux1h_1196_nl;
  wire[21:0] AccumDotWidth_acc_2587_nl;
  wire[22:0] nl_AccumDotWidth_acc_2587_nl;
  wire[21:0] AccumDotWidth_mux1h_1197_nl;
  wire[21:0] AccumDotWidth_acc_2588_nl;
  wire[22:0] nl_AccumDotWidth_acc_2588_nl;
  wire[21:0] AccumDotWidth_mux1h_1198_nl;
  wire[21:0] MultLoop_acc_1594_nl;
  wire[22:0] nl_MultLoop_acc_1594_nl;
  wire[21:0] AccumDotWidth_mux1h_1199_nl;
  wire[21:0] MultLoop_acc_1595_nl;
  wire[22:0] nl_MultLoop_acc_1595_nl;
  wire[21:0] MultLoop_mux1h_503_nl;
  wire[21:0] AccumDotWidth_acc_2589_nl;
  wire[22:0] nl_AccumDotWidth_acc_2589_nl;
  wire[21:0] MultLoop_mux1h_504_nl;
  wire[21:0] AccumDotWidth_acc_2590_nl;
  wire[22:0] nl_AccumDotWidth_acc_2590_nl;
  wire[21:0] AccumDotWidth_mux1h_1200_nl;
  wire[21:0] AccumDotWidth_acc_2591_nl;
  wire[22:0] nl_AccumDotWidth_acc_2591_nl;
  wire[21:0] AccumDotWidth_acc_2592_nl;
  wire[22:0] nl_AccumDotWidth_acc_2592_nl;
  wire[21:0] AccumDotWidth_mux1h_1201_nl;
  wire[21:0] AccumDotWidth_acc_2593_nl;
  wire[22:0] nl_AccumDotWidth_acc_2593_nl;
  wire[21:0] AccumDotWidth_acc_2594_nl;
  wire[22:0] nl_AccumDotWidth_acc_2594_nl;
  wire[21:0] MultLoop_mux1h_505_nl;
  wire[21:0] AccumDotWidth_acc_2595_nl;
  wire[22:0] nl_AccumDotWidth_acc_2595_nl;
  wire[21:0] MultLoop_mux1h_506_nl;
  wire[21:0] AccumDotWidth_acc_2596_nl;
  wire[22:0] nl_AccumDotWidth_acc_2596_nl;
  wire[21:0] AccumDotWidth_mux1h_1202_nl;
  wire[21:0] AccumDotWidth_acc_2597_nl;
  wire[22:0] nl_AccumDotWidth_acc_2597_nl;
  wire[21:0] AccumDotWidth_mux1h_1203_nl;
  wire[21:0] AccumDotWidth_acc_2598_nl;
  wire[22:0] nl_AccumDotWidth_acc_2598_nl;
  wire[21:0] AccumDotWidth_mux1h_1204_nl;
  wire[21:0] AccumDotWidth_acc_2599_nl;
  wire[22:0] nl_AccumDotWidth_acc_2599_nl;
  wire[21:0] AccumDotWidth_acc_2600_nl;
  wire[22:0] nl_AccumDotWidth_acc_2600_nl;
  wire[21:0] AccumDotWidth_acc_2601_nl;
  wire[22:0] nl_AccumDotWidth_acc_2601_nl;
  wire[21:0] AccumDotWidth_acc_2602_nl;
  wire[22:0] nl_AccumDotWidth_acc_2602_nl;
  wire[28:0] MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1205_nl;
  wire[21:0] AccumDotWidth_acc_2603_nl;
  wire[22:0] nl_AccumDotWidth_acc_2603_nl;
  wire[21:0] AccumDotWidth_acc_2604_nl;
  wire[22:0] nl_AccumDotWidth_acc_2604_nl;
  wire[21:0] AccumDotWidth_acc_2605_nl;
  wire[22:0] nl_AccumDotWidth_acc_2605_nl;
  wire[21:0] AccumDotWidth_acc_2606_nl;
  wire[22:0] nl_AccumDotWidth_acc_2606_nl;
  wire[28:0] MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1206_nl;
  wire[21:0] AccumDotWidth_acc_2607_nl;
  wire[22:0] nl_AccumDotWidth_acc_2607_nl;
  wire[21:0] AccumDotWidth_acc_2608_nl;
  wire[22:0] nl_AccumDotWidth_acc_2608_nl;
  wire[21:0] AccumDotWidth_acc_2609_nl;
  wire[22:0] nl_AccumDotWidth_acc_2609_nl;
  wire[21:0] AccumDotWidth_acc_2610_nl;
  wire[22:0] nl_AccumDotWidth_acc_2610_nl;
  wire[28:0] MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1207_nl;
  wire[21:0] AccumDotWidth_acc_2611_nl;
  wire[22:0] nl_AccumDotWidth_acc_2611_nl;
  wire[21:0] AccumDotWidth_acc_2612_nl;
  wire[22:0] nl_AccumDotWidth_acc_2612_nl;
  wire[21:0] AccumDotWidth_acc_2613_nl;
  wire[22:0] nl_AccumDotWidth_acc_2613_nl;
  wire[21:0] AccumDotWidth_acc_2614_nl;
  wire[22:0] nl_AccumDotWidth_acc_2614_nl;
  wire[28:0] MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1208_nl;
  wire[21:0] AccumDotWidth_acc_2615_nl;
  wire[22:0] nl_AccumDotWidth_acc_2615_nl;
  wire[28:0] MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1209_nl;
  wire[21:0] AccumDotWidth_acc_2616_nl;
  wire[22:0] nl_AccumDotWidth_acc_2616_nl;
  wire[28:0] MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1210_nl;
  wire[28:0] MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1211_nl;
  wire[28:0] MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1212_nl;
  wire[21:0] AccumDotWidth_acc_2617_nl;
  wire[22:0] nl_AccumDotWidth_acc_2617_nl;
  wire[21:0] AccumDotWidth_mux1h_1213_nl;
  wire[21:0] AccumDotWidth_mux1h_1214_nl;
  wire[21:0] AccumDotWidth_acc_2618_nl;
  wire[22:0] nl_AccumDotWidth_acc_2618_nl;
  wire[21:0] AccumDotWidth_mux1h_1215_nl;
  wire[21:0] AccumDotWidth_acc_2619_nl;
  wire[22:0] nl_AccumDotWidth_acc_2619_nl;
  wire[21:0] AccumDotWidth_mux1h_1216_nl;
  wire[21:0] AccumDotWidth_mux1h_1217_nl;
  wire[21:0] AccumDotWidth_mux1h_1218_nl;
  wire[21:0] MultLoop_acc_1596_nl;
  wire[22:0] nl_MultLoop_acc_1596_nl;
  wire[21:0] AccumDotWidth_mux1h_1219_nl;
  wire[21:0] MultLoop_acc_1597_nl;
  wire[22:0] nl_MultLoop_acc_1597_nl;
  wire[21:0] AccumDotWidth_mux1h_1220_nl;
  wire[21:0] AccumDotWidth_mux1h_1221_nl;
  wire[21:0] MultLoop_mux_97_nl;
  wire[28:0] MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_mux_98_nl;
  wire[21:0] AccumDotWidth_mux1h_1222_nl;
  wire[21:0] MultLoop_acc_1598_nl;
  wire[22:0] nl_MultLoop_acc_1598_nl;
  wire[10:0] MultLoop_acc_1599_nl;
  wire[11:0] nl_MultLoop_acc_1599_nl;
  wire[21:0] AccumDotWidth_mux1h_1223_nl;
  wire[21:0] MultLoop_acc_1600_nl;
  wire[22:0] nl_MultLoop_acc_1600_nl;
  wire[21:0] AccumDotWidth_mux1h_1224_nl;
  wire[21:0] AccumDotWidth_acc_2620_nl;
  wire[24:0] nl_AccumDotWidth_acc_2620_nl;
  wire[9:0] AccumDotWidth_acc_2625_nl;
  wire[10:0] nl_AccumDotWidth_acc_2625_nl;
  wire[21:0] AccumDotWidth_acc_2626_nl;
  wire[22:0] nl_AccumDotWidth_acc_2626_nl;
  wire[21:0] AccumDotWidth_acc_2627_nl;
  wire[23:0] nl_AccumDotWidth_acc_2627_nl;
  wire[9:0] AccumDotWidth_acc_2629_nl;
  wire[10:0] nl_AccumDotWidth_acc_2629_nl;
  wire[21:0] MultLoop_acc_1601_nl;
  wire[22:0] nl_MultLoop_acc_1601_nl;
  wire[10:0] MultLoop_acc_1602_nl;
  wire[11:0] nl_MultLoop_acc_1602_nl;
  wire[21:0] AccumDotWidth_mux1h_1225_nl;
  wire[21:0] AccumDotWidth_mux1h_1226_nl;
  wire[21:0] AccumDotWidth_acc_2630_nl;
  wire[24:0] nl_AccumDotWidth_acc_2630_nl;
  wire[9:0] AccumDotWidth_acc_2635_nl;
  wire[10:0] nl_AccumDotWidth_acc_2635_nl;
  wire[21:0] AccumDotWidth_acc_2636_nl;
  wire[22:0] nl_AccumDotWidth_acc_2636_nl;
  wire[21:0] AccumDotWidth_acc_2637_nl;
  wire[23:0] nl_AccumDotWidth_acc_2637_nl;
  wire[21:0] AccumDotWidth_acc_2640_nl;
  wire[24:0] nl_AccumDotWidth_acc_2640_nl;
  wire[9:0] AccumDotWidth_acc_2645_nl;
  wire[10:0] nl_AccumDotWidth_acc_2645_nl;
  wire[21:0] MultLoop_acc_1603_nl;
  wire[22:0] nl_MultLoop_acc_1603_nl;
  wire[10:0] MultLoop_acc_1604_nl;
  wire[11:0] nl_MultLoop_acc_1604_nl;
  wire[21:0] AccumDotWidth_mux1h_1227_nl;
  wire[21:0] AccumDotWidth_acc_2646_nl;
  wire[22:0] nl_AccumDotWidth_acc_2646_nl;
  wire[21:0] AccumDotWidth_acc_2647_nl;
  wire[23:0] nl_AccumDotWidth_acc_2647_nl;
  wire[21:0] AccumDotWidth_mux1h_1228_nl;
  wire[21:0] MultLoop_acc_1605_nl;
  wire[22:0] nl_MultLoop_acc_1605_nl;
  wire[10:0] MultLoop_acc_1606_nl;
  wire[11:0] nl_MultLoop_acc_1606_nl;
  wire[28:0] MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1229_nl;
  wire[21:0] MultLoop_acc_1607_nl;
  wire[22:0] nl_MultLoop_acc_1607_nl;
  wire[28:0] MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[28:0] MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1230_nl;
  wire[21:0] AccumDotWidth_acc_2650_nl;
  wire[24:0] nl_AccumDotWidth_acc_2650_nl;
  wire[9:0] AccumDotWidth_acc_2655_nl;
  wire[10:0] nl_AccumDotWidth_acc_2655_nl;
  wire[21:0] AccumDotWidth_acc_2656_nl;
  wire[24:0] nl_AccumDotWidth_acc_2656_nl;
  wire[21:0] AccumDotWidth_acc_2660_nl;
  wire[23:0] nl_AccumDotWidth_acc_2660_nl;
  wire[21:0] AccumDotWidth_acc_2663_nl;
  wire[24:0] nl_AccumDotWidth_acc_2663_nl;
  wire[9:0] AccumDotWidth_acc_2668_nl;
  wire[10:0] nl_AccumDotWidth_acc_2668_nl;
  wire[21:0] AccumDotWidth_mux1h_1231_nl;
  wire[21:0] AccumDotWidth_acc_2669_nl;
  wire[24:0] nl_AccumDotWidth_acc_2669_nl;
  wire[21:0] AccumDotWidth_acc_2673_nl;
  wire[23:0] nl_AccumDotWidth_acc_2673_nl;
  wire[21:0] MultLoop_acc_1608_nl;
  wire[22:0] nl_MultLoop_acc_1608_nl;
  wire[21:0] AccumDotWidth_mux1h_1232_nl;
  wire[21:0] AccumDotWidth_acc_2676_nl;
  wire[22:0] nl_AccumDotWidth_acc_2676_nl;
  wire[21:0] AccumDotWidth_mux1h_1233_nl;
  wire[21:0] AccumDotWidth_acc_2677_nl;
  wire[22:0] nl_AccumDotWidth_acc_2677_nl;
  wire[29:0] mul_160_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_805_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_806_nl;
  wire[29:0] mul_161_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_807_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_808_nl;
  wire[29:0] mul_162_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_809_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_810_nl;
  wire[29:0] mul_163_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_811_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_812_nl;
  wire[29:0] mul_164_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_813_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_36_nl;
  wire[29:0] mul_165_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_814_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_815_nl;
  wire[29:0] mul_166_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_816_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_817_nl;
  wire[29:0] mul_167_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_818_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_819_nl;
  wire[29:0] mul_168_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_820_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_821_nl;
  wire[29:0] mul_169_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_822_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_823_nl;
  wire[29:0] mul_170_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_824_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_825_nl;
  wire[29:0] mul_171_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_826_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_827_nl;
  wire[29:0] mul_172_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_828_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_829_nl;
  wire[29:0] mul_173_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_830_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_831_nl;
  wire[29:0] mul_174_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_832_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_833_nl;
  wire[29:0] mul_175_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_834_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_835_nl;
  wire[29:0] mul_176_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_836_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_837_nl;
  wire[29:0] mul_177_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_838_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_839_nl;
  wire[29:0] mul_178_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_840_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_841_nl;
  wire[29:0] mul_179_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_842_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_843_nl;
  wire[29:0] mul_180_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_844_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_845_nl;
  wire[29:0] mul_181_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_846_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_847_nl;
  wire[29:0] mul_182_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_848_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_849_nl;
  wire[29:0] mul_183_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_850_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_851_nl;
  wire[29:0] mul_184_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_852_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_853_nl;
  wire[29:0] mul_185_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_854_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_855_nl;
  wire[29:0] mul_186_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_856_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_857_nl;
  wire[29:0] mul_187_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_858_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_859_nl;
  wire[29:0] mul_188_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_860_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_861_nl;
  wire[29:0] mul_189_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_862_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_863_nl;
  wire[29:0] mul_190_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_864_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_865_nl;
  wire[29:0] mul_191_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_866_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_867_nl;
  wire[29:0] mul_192_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_868_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_869_nl;
  wire[29:0] mul_193_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_870_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_871_nl;
  wire[29:0] mul_194_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_872_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_873_nl;
  wire[29:0] mul_195_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_874_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_875_nl;
  wire[29:0] mul_196_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_876_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_877_nl;
  wire[29:0] mul_197_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_878_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_879_nl;
  wire[29:0] mul_198_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_880_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_881_nl;
  wire[29:0] mul_199_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_882_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_883_nl;
  wire[29:0] mul_200_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_884_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_885_nl;
  wire[29:0] mul_201_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_886_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_887_nl;
  wire[29:0] mul_202_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_888_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_889_nl;
  wire[29:0] mul_203_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_890_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_891_nl;
  wire[29:0] mul_204_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_892_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_893_nl;
  wire[29:0] mul_205_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_894_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_895_nl;
  wire[29:0] mul_206_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_896_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_897_nl;
  wire[29:0] mul_207_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_898_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_899_nl;
  wire[29:0] mul_208_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_900_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_901_nl;
  wire[29:0] mul_209_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_902_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_903_nl;
  wire[29:0] mul_210_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_904_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_37_nl;
  wire[29:0] mul_211_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_905_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_906_nl;
  wire[29:0] mul_212_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_574_nl;
  wire[21:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_575_nl;
  wire[0:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_52_nl;
  wire[29:0] mul_213_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_907_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_38_nl;
  wire[29:0] mul_214_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_908_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_39_nl;
  wire[29:0] mul_215_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_576_nl;
  wire[21:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_577_nl;
  wire[29:0] mul_216_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_909_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_910_nl;
  wire[29:0] mul_217_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_911_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_912_nl;
  wire[29:0] mul_218_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_913_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_914_nl;
  wire[29:0] mul_219_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_915_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_916_nl;
  wire[29:0] mul_220_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_917_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_918_nl;
  wire[29:0] mul_221_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_919_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_920_nl;
  wire[29:0] mul_222_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_921_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_922_nl;
  wire[28:0] mul_223_nl;
  wire signed [29:0] nl_mul_223_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_578_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_579_nl;
  wire[28:0] mul_224_nl;
  wire signed [29:0] nl_mul_224_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_580_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_581_nl;
  wire[28:0] mul_225_nl;
  wire signed [29:0] nl_mul_225_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_582_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_583_nl;
  wire[28:0] mul_226_nl;
  wire signed [29:0] nl_mul_226_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_584_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_585_nl;
  wire[28:0] mul_227_nl;
  wire signed [29:0] nl_mul_227_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_135_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_136_nl;
  wire[28:0] mul_228_nl;
  wire signed [29:0] nl_mul_228_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_586_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_587_nl;
  wire[28:0] mul_229_nl;
  wire signed [29:0] nl_mul_229_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_588_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_589_nl;
  wire[28:0] mul_230_nl;
  wire signed [29:0] nl_mul_230_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_590_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_591_nl;
  wire[28:0] mul_231_nl;
  wire signed [29:0] nl_mul_231_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_137_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_138_nl;
  wire[28:0] mul_232_nl;
  wire signed [29:0] nl_mul_232_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_139_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_140_nl;
  wire[28:0] mul_233_nl;
  wire signed [29:0] nl_mul_233_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_592_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_593_nl;
  wire[28:0] mul_234_nl;
  wire signed [29:0] nl_mul_234_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_594_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_595_nl;
  wire[28:0] mul_235_nl;
  wire signed [29:0] nl_mul_235_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_596_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_597_nl;
  wire[28:0] mul_236_nl;
  wire signed [29:0] nl_mul_236_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_598_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_599_nl;
  wire[28:0] mul_237_nl;
  wire signed [29:0] nl_mul_237_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_600_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_601_nl;
  wire[28:0] mul_238_nl;
  wire signed [29:0] nl_mul_238_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_602_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_603_nl;
  wire[28:0] mul_239_nl;
  wire signed [29:0] nl_mul_239_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_604_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_605_nl;
  wire[28:0] mul_240_nl;
  wire signed [29:0] nl_mul_240_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_606_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_607_nl;
  wire[28:0] mul_241_nl;
  wire signed [29:0] nl_mul_241_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_608_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_609_nl;
  wire[28:0] mul_242_nl;
  wire signed [29:0] nl_mul_242_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_610_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_611_nl;
  wire[28:0] mul_243_nl;
  wire signed [29:0] nl_mul_243_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_612_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_613_nl;
  wire[28:0] mul_244_nl;
  wire signed [29:0] nl_mul_244_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_614_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_615_nl;
  wire[28:0] mul_245_nl;
  wire signed [29:0] nl_mul_245_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_141_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_142_nl;
  wire[28:0] mul_246_nl;
  wire signed [29:0] nl_mul_246_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_143_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_144_nl;
  wire[28:0] mul_247_nl;
  wire signed [29:0] nl_mul_247_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_616_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_617_nl;
  wire[28:0] mul_248_nl;
  wire signed [29:0] nl_mul_248_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_618_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_619_nl;
  wire[28:0] mul_249_nl;
  wire signed [29:0] nl_mul_249_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_620_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_621_nl;
  wire[28:0] mul_250_nl;
  wire signed [29:0] nl_mul_250_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_622_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_623_nl;
  wire[28:0] mul_251_nl;
  wire signed [29:0] nl_mul_251_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_624_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_625_nl;
  wire[28:0] mul_252_nl;
  wire signed [29:0] nl_mul_252_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_626_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_627_nl;
  wire[28:0] mul_253_nl;
  wire signed [29:0] nl_mul_253_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_628_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_629_nl;
  wire[28:0] mul_254_nl;
  wire signed [29:0] nl_mul_254_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_630_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_631_nl;
  wire[28:0] mul_255_nl;
  wire signed [29:0] nl_mul_255_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_632_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_633_nl;
  wire[28:0] mul_256_nl;
  wire signed [29:0] nl_mul_256_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_634_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_635_nl;
  wire[28:0] mul_257_nl;
  wire signed [29:0] nl_mul_257_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_636_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_637_nl;
  wire[28:0] mul_258_nl;
  wire signed [29:0] nl_mul_258_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_638_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_639_nl;
  wire[28:0] mul_259_nl;
  wire signed [29:0] nl_mul_259_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_640_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_145_nl;
  wire[28:0] mul_260_nl;
  wire signed [29:0] nl_mul_260_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_641_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_146_nl;
  wire[28:0] mul_261_nl;
  wire signed [29:0] nl_mul_261_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_642_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_147_nl;
  wire[28:0] mul_262_nl;
  wire signed [29:0] nl_mul_262_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_643_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_8_nl;
  wire[28:0] mul_263_nl;
  wire signed [29:0] nl_mul_263_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_644_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_9_nl;
  wire[28:0] mul_264_nl;
  wire signed [29:0] nl_mul_264_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_645_nl;
  wire[28:0] mul_265_nl;
  wire signed [29:0] nl_mul_265_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_646_nl;
  wire[28:0] mul_266_nl;
  wire signed [29:0] nl_mul_266_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_647_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_10_nl;
  wire[28:0] mul_267_nl;
  wire signed [29:0] nl_mul_267_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_648_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_11_nl;
  wire[28:0] mul_268_nl;
  wire signed [29:0] nl_mul_268_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_649_nl;
  wire[20:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_12_nl;
  wire[28:0] mul_269_nl;
  wire signed [29:0] nl_mul_269_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_148_nl;
  wire[28:0] mul_270_nl;
  wire signed [29:0] nl_mul_270_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_149_nl;
  wire[28:0] mul_271_nl;
  wire signed [29:0] nl_mul_271_nl;
  wire[7:0] nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_150_nl;
  wire[20:0] AccumDotWidth_mux1h_1234_nl;
  wire[9:0] AccumDotWidth_acc_2678_nl;
  wire[10:0] nl_AccumDotWidth_acc_2678_nl;
  wire[20:0] AccumDotWidth_mux1h_1235_nl;
  wire[20:0] AccumDotWidth_mux1h_1236_nl;
  wire[9:0] AccumDotWidth_acc_2679_nl;
  wire[10:0] nl_AccumDotWidth_acc_2679_nl;
  wire[9:0] AccumDotWidth_acc_2680_nl;
  wire[10:0] nl_AccumDotWidth_acc_2680_nl;
  wire[20:0] AccumDotWidth_mux1h_1237_nl;
  wire[20:0] AccumDotWidth_mux1h_1238_nl;
  wire[20:0] AccumDotWidth_mux1h_1239_nl;
  wire[9:0] AccumDotWidth_mux1h_1240_nl;
  wire[9:0] AccumDotWidth_acc_2681_nl;
  wire[10:0] nl_AccumDotWidth_acc_2681_nl;
  wire[9:0] AccumDotWidth_acc_2682_nl;
  wire[10:0] nl_AccumDotWidth_acc_2682_nl;
  wire[10:0] AccumDotWidth_mux1h_1241_nl;
  wire[20:0] AccumDotWidth_mux1h_1242_nl;
  wire[20:0] AccumDotWidth_mux1h_1243_nl;
  wire[9:0] AccumDotWidth_acc_2683_nl;
  wire[10:0] nl_AccumDotWidth_acc_2683_nl;
  wire[9:0] AccumDotWidth_acc_2684_nl;
  wire[10:0] nl_AccumDotWidth_acc_2684_nl;
  wire[20:0] AccumDotWidth_mux1h_1244_nl;
  wire[9:0] AccumDotWidth_mux1h_1245_nl;
  wire[9:0] AccumDotWidth_acc_2730_nl;
  wire[10:0] nl_AccumDotWidth_acc_2730_nl;
  wire[9:0] AccumDotWidth_mux1h_754_nl;
  wire[7:0] AccumDotWidth_AccumDotWidth_mux_17_nl;
  wire[9:0] AccumDotWidth_acc_2685_nl;
  wire[10:0] nl_AccumDotWidth_acc_2685_nl;
  wire[0:0] AccumDotWidth_or_209_nl;
  wire[10:0] AccumDotWidth_mux1h_1246_nl;
  wire[20:0] AccumDotWidth_mux1h_1247_nl;
  wire[9:0] AccumDotWidth_mux1h_1248_nl;
  wire[9:0] AccumDotWidth_acc_2686_nl;
  wire[10:0] nl_AccumDotWidth_acc_2686_nl;
  wire[9:0] AccumDotWidth_acc_2687_nl;
  wire[10:0] nl_AccumDotWidth_acc_2687_nl;
  wire[10:0] AccumDotWidth_mux1h_1249_nl;
  wire[20:0] AccumDotWidth_mux1h_1250_nl;
  wire[9:0] AccumDotWidth_mux1h_1251_nl;
  wire[9:0] AccumDotWidth_acc_2728_nl;
  wire[10:0] nl_AccumDotWidth_acc_2728_nl;
  wire[9:0] AccumDotWidth_mux_79_nl;
  wire[7:0] AccumDotWidth_mux_80_nl;
  wire[9:0] AccumDotWidth_acc_2688_nl;
  wire[10:0] nl_AccumDotWidth_acc_2688_nl;
  wire[10:0] AccumDotWidth_mux1h_1252_nl;
  wire[20:0] AccumDotWidth_mux1h_1253_nl;
  wire[20:0] AccumDotWidth_mux1h_1254_nl;
  wire[20:0] AccumDotWidth_mux1h_1255_nl;
  wire[20:0] AccumDotWidth_mux1h_1256_nl;
  wire[20:0] AccumDotWidth_mux1h_1257_nl;
  wire[20:0] AccumDotWidth_mux1h_1258_nl;
  wire[20:0] AccumDotWidth_mux1h_1259_nl;
  wire[20:0] AccumDotWidth_mux1h_1260_nl;
  wire[20:0] AccumDotWidth_mux1h_1261_nl;
  wire[20:0] AccumDotWidth_mux1h_1262_nl;
  wire[20:0] AccumDotWidth_mux1h_1263_nl;
  wire[20:0] AccumDotWidth_mux1h_1264_nl;
  wire[20:0] AccumDotWidth_mux1h_1265_nl;
  wire[20:0] AccumDotWidth_mux1h_1266_nl;
  wire[20:0] AccumDotWidth_mux1h_1267_nl;
  wire[20:0] AccumDotWidth_mux1h_1268_nl;
  wire[20:0] AccumDotWidth_mux1h_1269_nl;
  wire[20:0] AccumDotWidth_mux1h_1270_nl;
  wire[20:0] AccumDotWidth_mux1h_1271_nl;
  wire[20:0] AccumDotWidth_mux1h_1272_nl;
  wire[20:0] AccumDotWidth_mux1h_1273_nl;
  wire[20:0] AccumDotWidth_mux1h_1274_nl;
  wire[20:0] AccumDotWidth_mux1h_1275_nl;
  wire[20:0] AccumDotWidth_mux1h_1276_nl;
  wire[20:0] AccumDotWidth_mux1h_1277_nl;
  wire[20:0] AccumDotWidth_mux1h_1278_nl;
  wire[20:0] AccumDotWidth_mux1h_1279_nl;
  wire[20:0] AccumDotWidth_mux1h_1280_nl;
  wire[20:0] AccumDotWidth_mux1h_1281_nl;
  wire[20:0] AccumDotWidth_mux1h_1282_nl;
  wire[20:0] AccumDotWidth_mux1h_1283_nl;
  wire[20:0] AccumDotWidth_mux1h_1284_nl;
  wire[20:0] AccumDotWidth_mux1h_1285_nl;
  wire[20:0] AccumDotWidth_mux1h_1286_nl;
  wire[20:0] AccumDotWidth_mux1h_1287_nl;
  wire[20:0] AccumDotWidth_mux1h_1288_nl;
  wire[20:0] AccumDotWidth_mux1h_1289_nl;
  wire[20:0] AccumDotWidth_mux1h_1290_nl;
  wire[20:0] AccumDotWidth_mux1h_1291_nl;
  wire[20:0] AccumDotWidth_mux1h_1292_nl;
  wire[20:0] AccumDotWidth_mux1h_1293_nl;
  wire[20:0] AccumDotWidth_mux1h_1294_nl;
  wire[20:0] AccumDotWidth_mux1h_1295_nl;
  wire[20:0] AccumDotWidth_mux1h_1296_nl;
  wire[20:0] AccumDotWidth_mux1h_1297_nl;
  wire[20:0] AccumDotWidth_mux1h_1298_nl;
  wire[20:0] AccumDotWidth_mux1h_1299_nl;
  wire[20:0] AccumDotWidth_mux1h_1300_nl;
  wire[20:0] AccumDotWidth_mux1h_1301_nl;
  wire[20:0] AccumDotWidth_mux1h_1302_nl;
  wire[20:0] AccumDotWidth_mux1h_1303_nl;
  wire[20:0] AccumDotWidth_mux1h_1304_nl;
  wire[20:0] AccumDotWidth_mux1h_1305_nl;
  wire[20:0] AccumDotWidth_mux1h_1306_nl;
  wire[20:0] AccumDotWidth_mux1h_1307_nl;
  wire[20:0] AccumDotWidth_mux1h_1308_nl;
  wire[20:0] AccumDotWidth_mux1h_1309_nl;
  wire[20:0] AccumDotWidth_mux1h_1310_nl;
  wire[20:0] AccumDotWidth_mux1h_1311_nl;
  wire[20:0] AccumDotWidth_mux1h_1312_nl;
  wire[20:0] AccumDotWidth_mux1h_1313_nl;
  wire[20:0] AccumDotWidth_mux1h_1314_nl;
  wire[20:0] AccumDotWidth_mux1h_1315_nl;
  wire[20:0] AccumDotWidth_mux1h_1316_nl;
  wire[20:0] AccumDotWidth_mux1h_1317_nl;
  wire[20:0] AccumDotWidth_mux1h_1318_nl;
  wire[20:0] AccumDotWidth_mux1h_1319_nl;
  wire[20:0] AccumDotWidth_mux1h_1320_nl;
  wire[20:0] AccumDotWidth_mux1h_1321_nl;
  wire[20:0] AccumDotWidth_mux1h_1322_nl;
  wire[20:0] AccumDotWidth_mux1h_1323_nl;
  wire[20:0] AccumDotWidth_mux1h_1324_nl;
  wire[20:0] AccumDotWidth_mux1h_1325_nl;
  wire[20:0] AccumDotWidth_mux1h_1326_nl;
  wire[20:0] AccumDotWidth_mux1h_1327_nl;
  wire[20:0] AccumDotWidth_mux1h_1328_nl;
  wire[20:0] AccumDotWidth_mux1h_1329_nl;
  wire[20:0] AccumDotWidth_mux1h_1330_nl;
  wire[20:0] AccumDotWidth_mux1h_1331_nl;
  wire[20:0] AccumDotWidth_mux1h_1332_nl;
  wire[20:0] AccumDotWidth_mux1h_1333_nl;
  wire[20:0] AccumDotWidth_mux1h_1334_nl;
  wire[20:0] AccumDotWidth_mux1h_1335_nl;
  wire[20:0] AccumDotWidth_mux1h_1336_nl;
  wire[20:0] AccumDotWidth_mux1h_1337_nl;
  wire[20:0] AccumDotWidth_mux1h_1338_nl;
  wire[20:0] AccumDotWidth_mux1h_1339_nl;
  wire[20:0] AccumDotWidth_mux1h_1340_nl;
  wire[20:0] AccumDotWidth_mux1h_1341_nl;
  wire[20:0] AccumDotWidth_mux1h_1342_nl;
  wire[20:0] AccumDotWidth_mux1h_1343_nl;
  wire[20:0] AccumDotWidth_mux1h_1344_nl;
  wire[20:0] AccumDotWidth_mux1h_1345_nl;
  wire[20:0] AccumDotWidth_mux1h_1346_nl;
  wire[20:0] AccumDotWidth_mux1h_1347_nl;
  wire[20:0] AccumDotWidth_mux1h_1348_nl;
  wire[20:0] AccumDotWidth_mux1h_1349_nl;
  wire[20:0] AccumDotWidth_mux1h_1350_nl;
  wire[20:0] AccumDotWidth_mux1h_1351_nl;
  wire[20:0] AccumDotWidth_mux1h_1352_nl;
  wire[20:0] AccumDotWidth_mux1h_1353_nl;
  wire[20:0] AccumDotWidth_mux1h_1354_nl;
  wire[20:0] AccumDotWidth_mux1h_1355_nl;
  wire[20:0] AccumDotWidth_mux1h_1356_nl;
  wire[20:0] AccumDotWidth_mux1h_1357_nl;
  wire[20:0] AccumDotWidth_mux1h_1358_nl;
  wire[20:0] AccumDotWidth_mux1h_1359_nl;
  wire[20:0] AccumDotWidth_mux1h_1360_nl;
  wire[20:0] AccumDotWidth_mux1h_1361_nl;
  wire[20:0] AccumDotWidth_mux1h_1362_nl;
  wire[20:0] AccumDotWidth_mux1h_1363_nl;
  wire[20:0] AccumDotWidth_mux1h_1364_nl;
  wire[20:0] AccumDotWidth_mux1h_1365_nl;
  wire[20:0] AccumDotWidth_mux1h_1366_nl;
  wire[20:0] AccumDotWidth_mux1h_1367_nl;
  wire[20:0] AccumDotWidth_mux1h_1368_nl;
  wire[20:0] AccumDotWidth_mux1h_1369_nl;
  wire[20:0] AccumDotWidth_mux1h_1370_nl;
  wire[20:0] AccumDotWidth_mux1h_1371_nl;
  wire[20:0] AccumDotWidth_mux1h_1372_nl;
  wire[20:0] AccumDotWidth_mux1h_1373_nl;
  wire[20:0] AccumDotWidth_mux1h_1374_nl;
  wire[20:0] AccumDotWidth_mux1h_1375_nl;
  wire[20:0] AccumDotWidth_mux1h_1376_nl;
  wire[20:0] AccumDotWidth_mux1h_1377_nl;
  wire[20:0] AccumDotWidth_mux_143_nl;
  wire[20:0] AccumDotWidth_mux_144_nl;
  wire[21:0] AccumDotWidth_mux1h_1378_nl;
  wire[21:0] AccumDotWidth_mux1h_1379_nl;
  wire[21:0] AccumDotWidth_mux1h_1380_nl;
  wire[21:0] MultLoop_acc_1609_nl;
  wire[22:0] nl_MultLoop_acc_1609_nl;
  wire[21:0] MultLoop_acc_1610_nl;
  wire[22:0] nl_MultLoop_acc_1610_nl;
  wire[21:0] MultLoop_acc_1611_nl;
  wire[22:0] nl_MultLoop_acc_1611_nl;
  wire[21:0] MultLoop_acc_1612_nl;
  wire[22:0] nl_MultLoop_acc_1612_nl;
  wire[21:0] AccumDotWidth_mux1h_1381_nl;
  wire[21:0] MultLoop_acc_1613_nl;
  wire[22:0] nl_MultLoop_acc_1613_nl;
  wire[21:0] MultLoop_mux1h_507_nl;
  wire[21:0] MultLoop_mux1h_508_nl;
  wire[21:0] AccumDotWidth_mux1h_1382_nl;
  wire[21:0] MultLoop_acc_1614_nl;
  wire[23:0] nl_MultLoop_acc_1614_nl;
  wire[21:0] MultLoop_acc_1616_nl;
  wire[22:0] nl_MultLoop_acc_1616_nl;
  wire[21:0] MultLoop_acc_1617_nl;
  wire[22:0] nl_MultLoop_acc_1617_nl;
  wire[21:0] AccumDotWidth_mux1h_1383_nl;
  wire[21:0] AccumDotWidth_mux1h_1384_nl;
  wire[21:0] MultLoop_acc_1618_nl;
  wire[22:0] nl_MultLoop_acc_1618_nl;
  wire[21:0] MultLoop_acc_1619_nl;
  wire[22:0] nl_MultLoop_acc_1619_nl;
  wire[21:0] MultLoop_acc_1620_nl;
  wire[22:0] nl_MultLoop_acc_1620_nl;
  wire[21:0] MultLoop_acc_1621_nl;
  wire[22:0] nl_MultLoop_acc_1621_nl;
  wire[21:0] AccumDotWidth_mux1h_1385_nl;
  wire[21:0] MultLoop_acc_1622_nl;
  wire[23:0] nl_MultLoop_acc_1622_nl;
  wire[21:0] MultLoop_acc_1624_nl;
  wire[22:0] nl_MultLoop_acc_1624_nl;
  wire[21:0] MultLoop_acc_1625_nl;
  wire[22:0] nl_MultLoop_acc_1625_nl;
  wire[21:0] MultLoop_acc_1627_nl;
  wire[22:0] nl_MultLoop_acc_1627_nl;
  wire[21:0] MultLoop_acc_1628_nl;
  wire[22:0] nl_MultLoop_acc_1628_nl;
  wire[21:0] AccumDotWidth_mux1h_1386_nl;
  wire[21:0] AccumDotWidth_mux1h_1387_nl;
  wire[21:0] MultLoop_acc_1629_nl;
  wire[23:0] nl_MultLoop_acc_1629_nl;
  wire[21:0] MultLoop_acc_1631_nl;
  wire[22:0] nl_MultLoop_acc_1631_nl;
  wire[21:0] MultLoop_acc_1632_nl;
  wire[22:0] nl_MultLoop_acc_1632_nl;
  wire[21:0] MultLoop_acc_1634_nl;
  wire[22:0] nl_MultLoop_acc_1634_nl;
  wire[21:0] MultLoop_acc_1635_nl;
  wire[22:0] nl_MultLoop_acc_1635_nl;
  wire[21:0] MultLoop_mux1h_509_nl;
  wire[21:0] MultLoop_mux1h_510_nl;
  wire[21:0] AccumDotWidth_mux1h_1388_nl;
  wire[21:0] AccumDotWidth_mux1h_1389_nl;
  wire[21:0] AccumDotWidth_mux1h_1390_nl;
  wire[21:0] MultLoop_acc_1636_nl;
  wire[22:0] nl_MultLoop_acc_1636_nl;
  wire[21:0] AccumDotWidth_mux1h_1391_nl;
  wire[21:0] AccumDotWidth_mux_145_nl;
  wire[21:0] AccumDotWidth_mux_146_nl;
  wire[21:0] MultLoop_mux1h_511_nl;
  wire[21:0] MultLoop_mux1h_512_nl;
  wire[21:0] AccumDotWidth_mux1h_1392_nl;
  wire[21:0] AccumDotWidth_mux1h_1393_nl;
  wire[21:0] AccumDotWidth_mux_147_nl;
  wire[21:0] AccumDotWidth_mux_148_nl;
  wire[21:0] MultLoop_mux_99_nl;
  wire[21:0] MultLoop_mux_100_nl;
  wire[21:0] AccumDotWidth_mux1h_1394_nl;
  wire[21:0] AccumDotWidth_mux1h_1395_nl;
  wire[21:0] AccumDotWidth_mux1h_1396_nl;
  wire[21:0] AccumDotWidth_mux1h_1397_nl;
  wire[21:0] MultLoop_mux1h_513_nl;
  wire[21:0] MultLoop_mux1h_514_nl;
  wire[21:0] MultLoop_mux1h_515_nl;
  wire[21:0] MultLoop_mux1h_516_nl;
  wire[21:0] MultLoop_mux1h_517_nl;
  wire[21:0] MultLoop_mux1h_518_nl;
  wire[21:0] MultLoop_mux1h_519_nl;
  wire[21:0] MultLoop_mux1h_520_nl;
  wire[21:0] MultLoop_mux1h_521_nl;
  wire[21:0] MultLoop_mux1h_522_nl;
  wire[21:0] MultLoop_acc_1637_nl;
  wire[22:0] nl_MultLoop_acc_1637_nl;
  wire[21:0] AccumDotWidth_mux1h_1398_nl;
  wire[21:0] AccumDotWidth_mux1h_1399_nl;
  wire[21:0] MultLoop_mux1h_523_nl;
  wire[21:0] MultLoop_mux1h_524_nl;
  wire[21:0] MultLoop_mux1h_525_nl;
  wire[21:0] MultLoop_mux1h_526_nl;
  wire[21:0] AccumDotWidth_mux1h_1400_nl;
  wire[21:0] AccumDotWidth_mux1h_1401_nl;
  wire[21:0] MultLoop_mux1h_527_nl;
  wire[21:0] MultLoop_mux1h_528_nl;
  wire[21:0] MultLoop_mux1h_529_nl;
  wire[21:0] MultLoop_mux1h_530_nl;
  wire[21:0] AccumDotWidth_mux1h_1402_nl;
  wire[21:0] AccumDotWidth_mux1h_1403_nl;
  wire[21:0] MultLoop_mux1h_531_nl;
  wire[0:0] MultLoop_or_113_nl;
  wire[21:0] MultLoop_mux1h_532_nl;
  wire[21:0] AccumDotWidth_mux_149_nl;
  wire[21:0] AccumDotWidth_mux_150_nl;
  wire[21:0] MultLoop_mux1h_533_nl;
  wire[21:0] MultLoop_mux1h_534_nl;
  wire[21:0] MultLoop_mux1h_535_nl;
  wire[21:0] MultLoop_mux1h_536_nl;
  wire[21:0] MultLoop_acc_1638_nl;
  wire[22:0] nl_MultLoop_acc_1638_nl;
  wire[21:0] MultLoop_mux1h_537_nl;
  wire[0:0] MultLoop_or_114_nl;
  wire[21:0] MultLoop_mux1h_538_nl;
  wire[21:0] MultLoop_mux1h_539_nl;
  wire[21:0] MultLoop_mux1h_540_nl;
  wire[21:0] MultLoop_mux1h_541_nl;
  wire[21:0] MultLoop_MultLoop_mux_15_nl;
  wire[21:0] MultLoop_mux1h_542_nl;
  wire[21:0] MultLoop_acc_1639_nl;
  wire[22:0] nl_MultLoop_acc_1639_nl;
  wire[21:0] MultLoop_acc_1640_nl;
  wire[22:0] nl_MultLoop_acc_1640_nl;
  wire[21:0] MultLoop_mux1h_543_nl;
  wire[21:0] MultLoop_acc_1641_nl;
  wire[22:0] nl_MultLoop_acc_1641_nl;
  wire[21:0] MultLoop_mux1h_544_nl;
  wire[21:0] MultLoop_mux1h_545_nl;
  wire[21:0] MultLoop_mux1h_546_nl;
  wire[21:0] MultLoop_mux1h_547_nl;
  wire[21:0] MultLoop_mux1h_548_nl;
  wire[21:0] MultLoop_mux1h_549_nl;
  wire[21:0] MultLoop_mux1h_550_nl;
  wire[21:0] MultLoop_mux1h_551_nl;
  wire[21:0] AccumDotWidth_mux_151_nl;
  wire[21:0] AccumDotWidth_mux_152_nl;
  wire[21:0] MultLoop_mux_101_nl;
  wire[21:0] MultLoop_mux_102_nl;
  wire[21:0] AccumDotWidth_mux1h_1404_nl;
  wire[21:0] AccumDotWidth_mux1h_1405_nl;
  wire[21:0] MultLoop_mux1h_552_nl;
  wire[21:0] MultLoop_mux1h_553_nl;
  wire[21:0] AccumDotWidth_mux1h_1406_nl;
  wire[21:0] AccumDotWidth_mux1h_1407_nl;
  wire[21:0] MultLoop_mux1h_554_nl;
  wire[21:0] MultLoop_mux1h_555_nl;
  wire[21:0] AccumDotWidth_mux1h_1408_nl;
  wire[21:0] AccumDotWidth_acc_2689_nl;
  wire[22:0] nl_AccumDotWidth_acc_2689_nl;
  wire[21:0] AccumDotWidth_acc_2690_nl;
  wire[22:0] nl_AccumDotWidth_acc_2690_nl;
  wire[21:0] AccumDotWidth_mux1h_1409_nl;
  wire[21:0] AccumDotWidth_acc_2691_nl;
  wire[22:0] nl_AccumDotWidth_acc_2691_nl;
  wire[21:0] AccumDotWidth_acc_2692_nl;
  wire[22:0] nl_AccumDotWidth_acc_2692_nl;
  wire[21:0] MultLoop_mux_103_nl;
  wire[21:0] MultLoop_mux_104_nl;
  wire[21:0] AccumDotWidth_mux1h_1410_nl;
  wire[21:0] AccumDotWidth_acc_2693_nl;
  wire[22:0] nl_AccumDotWidth_acc_2693_nl;
  wire[21:0] AccumDotWidth_acc_2694_nl;
  wire[22:0] nl_AccumDotWidth_acc_2694_nl;
  wire[21:0] AccumDotWidth_mux1h_1411_nl;
  wire[21:0] AccumDotWidth_acc_2695_nl;
  wire[22:0] nl_AccumDotWidth_acc_2695_nl;
  wire[21:0] AccumDotWidth_acc_2696_nl;
  wire[22:0] nl_AccumDotWidth_acc_2696_nl;
  wire[21:0] MultLoop_mux_105_nl;
  wire[21:0] MultLoop_mux_106_nl;
  wire[21:0] AccumDotWidth_mux_153_nl;
  wire[21:0] AccumDotWidth_acc_2697_nl;
  wire[22:0] nl_AccumDotWidth_acc_2697_nl;
  wire[21:0] AccumDotWidth_mux_154_nl;
  wire[21:0] AccumDotWidth_acc_2698_nl;
  wire[22:0] nl_AccumDotWidth_acc_2698_nl;
  wire[21:0] AccumDotWidth_mux1h_1412_nl;
  wire[21:0] AccumDotWidth_acc_2699_nl;
  wire[22:0] nl_AccumDotWidth_acc_2699_nl;
  wire[21:0] AccumDotWidth_acc_2700_nl;
  wire[22:0] nl_AccumDotWidth_acc_2700_nl;
  wire[21:0] AccumDotWidth_acc_2701_nl;
  wire[22:0] nl_AccumDotWidth_acc_2701_nl;
  wire[21:0] AccumDotWidth_mux1h_1413_nl;
  wire[21:0] AccumDotWidth_acc_2702_nl;
  wire[22:0] nl_AccumDotWidth_acc_2702_nl;
  wire[21:0] AccumDotWidth_acc_2703_nl;
  wire[22:0] nl_AccumDotWidth_acc_2703_nl;
  wire[21:0] AccumDotWidth_acc_2704_nl;
  wire[22:0] nl_AccumDotWidth_acc_2704_nl;
  wire[21:0] MultLoop_mux_107_nl;
  wire[21:0] MultLoop_mux_108_nl;
  wire[21:0] AccumDotWidth_mux1h_1414_nl;
  wire[21:0] AccumDotWidth_acc_2705_nl;
  wire[22:0] nl_AccumDotWidth_acc_2705_nl;
  wire[21:0] AccumDotWidth_mux1h_1415_nl;
  wire[21:0] AccumDotWidth_acc_2706_nl;
  wire[22:0] nl_AccumDotWidth_acc_2706_nl;
  wire[21:0] AccumDotWidth_mux1h_1416_nl;
  wire[21:0] AccumDotWidth_acc_2707_nl;
  wire[22:0] nl_AccumDotWidth_acc_2707_nl;
  wire[21:0] AccumDotWidth_acc_2708_nl;
  wire[22:0] nl_AccumDotWidth_acc_2708_nl;
  wire[21:0] AccumDotWidth_acc_2709_nl;
  wire[22:0] nl_AccumDotWidth_acc_2709_nl;
  wire[21:0] AccumDotWidth_mux1h_1417_nl;
  wire[21:0] AccumDotWidth_acc_2710_nl;
  wire[22:0] nl_AccumDotWidth_acc_2710_nl;
  wire[21:0] AccumDotWidth_acc_2711_nl;
  wire[22:0] nl_AccumDotWidth_acc_2711_nl;
  wire[21:0] AccumDotWidth_acc_2712_nl;
  wire[22:0] nl_AccumDotWidth_acc_2712_nl;
  wire[21:0] AccumDotWidth_mux1h_1418_nl;
  wire[10:0] MultLoop_acc_1642_nl;
  wire[11:0] nl_MultLoop_acc_1642_nl;
  wire[21:0] AccumDotWidth_mux1h_1419_nl;
  wire[21:0] AccumDotWidth_mux1h_1420_nl;
  wire[21:0] AccumDotWidth_acc_2713_nl;
  wire[22:0] nl_AccumDotWidth_acc_2713_nl;
  wire[21:0] AccumDotWidth_acc_2714_nl;
  wire[22:0] nl_AccumDotWidth_acc_2714_nl;
  wire[21:0] AccumDotWidth_acc_2715_nl;
  wire[22:0] nl_AccumDotWidth_acc_2715_nl;
  wire[21:0] AccumDotWidth_mux1h_1421_nl;
  wire[21:0] AccumDotWidth_acc_2716_nl;
  wire[22:0] nl_AccumDotWidth_acc_2716_nl;
  wire[21:0] AccumDotWidth_acc_2717_nl;
  wire[22:0] nl_AccumDotWidth_acc_2717_nl;
  wire[21:0] AccumDotWidth_acc_2718_nl;
  wire[22:0] nl_AccumDotWidth_acc_2718_nl;
  wire[21:0] AccumDotWidth_mux1h_1422_nl;
  wire[21:0] AccumDotWidth_mux1h_1423_nl;
  wire[21:0] AccumDotWidth_mux1h_1424_nl;
  wire[21:0] AccumDotWidth_mux1h_1425_nl;
  wire[21:0] MultLoop_mux_109_nl;
  wire[21:0] MultLoop_acc_1643_nl;
  wire[22:0] nl_MultLoop_acc_1643_nl;
  wire[21:0] MultLoop_mux_110_nl;
  wire[21:0] AccumDotWidth_mux1h_1426_nl;
  wire[21:0] MultLoop_acc_1644_nl;
  wire[22:0] nl_MultLoop_acc_1644_nl;
  wire[21:0] MultLoop_acc_1645_nl;
  wire[22:0] nl_MultLoop_acc_1645_nl;
  wire[21:0] AccumDotWidth_mux1h_1427_nl;
  wire[21:0] AccumDotWidth_mux1h_1428_nl;
  wire[21:0] AccumDotWidth_mux1h_1429_nl;
  wire[21:0] AccumDotWidth_mux1h_1430_nl;
  wire[21:0] AccumDotWidth_mux1h_1431_nl;
  wire[21:0] MultLoop_mux_111_nl;
  wire[21:0] MultLoop_mux_112_nl;
  wire[21:0] MultLoop_acc_1646_nl;
  wire[22:0] nl_MultLoop_acc_1646_nl;
  wire[21:0] AccumDotWidth_mux1h_1432_nl;
  wire[21:0] AccumDotWidth_acc_2719_nl;
  wire[22:0] nl_AccumDotWidth_acc_2719_nl;
  wire[21:0] MultLoop_acc_1647_nl;
  wire[23:0] nl_MultLoop_acc_1647_nl;
  wire[21:0] MultLoop_acc_1649_nl;
  wire[22:0] nl_MultLoop_acc_1649_nl;
  wire[28:0] MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] MultLoop_acc_1651_nl;
  wire[22:0] nl_MultLoop_acc_1651_nl;
  wire[21:0] MultLoop_acc_1652_nl;
  wire[22:0] nl_MultLoop_acc_1652_nl;
  wire[28:0] MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire signed [29:0] nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl;
  wire[21:0] AccumDotWidth_mux1h_1433_nl;
  wire[21:0] AccumDotWidth_mux1h_1434_nl;
  wire[21:0] MultLoop_acc_1653_nl;
  wire[22:0] nl_MultLoop_acc_1653_nl;
  wire[21:0] MultLoop_acc_1654_nl;
  wire[22:0] nl_MultLoop_acc_1654_nl;
  wire[21:0] AccumDotWidth_mux1h_1435_nl;
  wire[21:0] MultLoop_acc_1655_nl;
  wire[22:0] nl_MultLoop_acc_1655_nl;
  wire[21:0] MultLoop_acc_1656_nl;
  wire[22:0] nl_MultLoop_acc_1656_nl;
  wire[21:0] MultLoop_mux_113_nl;
  wire[21:0] MultLoop_mux_114_nl;
  wire[21:0] AccumDotWidth_mux1h_1436_nl;
  wire[21:0] AccumDotWidth_mux1h_1437_nl;
  wire[21:0] MultLoop_mux_115_nl;
  wire[21:0] MultLoop_mux_116_nl;
  wire[21:0] MultLoop_mux1h_556_nl;
  wire[21:0] MultLoop_mux1h_557_nl;
  wire[21:0] MultLoop_mux1h_558_nl;
  wire[21:0] MultLoop_mux1h_559_nl;
  wire[21:0] AccumDotWidth_mux_155_nl;
  wire[21:0] MultLoop_mux1h_560_nl;
  wire[21:0] MultLoop_acc_1657_nl;
  wire[22:0] nl_MultLoop_acc_1657_nl;
  wire[21:0] MultLoop_acc_1658_nl;
  wire[22:0] nl_MultLoop_acc_1658_nl;
  wire[21:0] MultLoop_acc_1659_nl;
  wire[22:0] nl_MultLoop_acc_1659_nl;
  wire[21:0] MultLoop_acc_1660_nl;
  wire[22:0] nl_MultLoop_acc_1660_nl;
  wire[21:0] MultLoop_mux1h_561_nl;
  wire[21:0] MultLoop_mux1h_562_nl;
  wire[21:0] MultLoop_acc_1661_nl;
  wire[22:0] nl_MultLoop_acc_1661_nl;
  wire[21:0] MultLoop_acc_1662_nl;
  wire[22:0] nl_MultLoop_acc_1662_nl;
  wire[21:0] MultLoop_acc_1663_nl;
  wire[22:0] nl_MultLoop_acc_1663_nl;
  wire[21:0] MultLoop_mux1h_563_nl;
  wire[21:0] MultLoop_acc_1664_nl;
  wire[22:0] nl_MultLoop_acc_1664_nl;
  wire[21:0] MultLoop_acc_1665_nl;
  wire[22:0] nl_MultLoop_acc_1665_nl;
  wire[21:0] MultLoop_acc_1666_nl;
  wire[22:0] nl_MultLoop_acc_1666_nl;
  wire[21:0] AccumDotWidth_AccumDotWidth_mux_22_nl;
  wire[21:0] AccumDotWidth_mux1h_1438_nl;
  wire[21:0] MultLoop_mux1h_564_nl;
  wire[21:0] MultLoop_mux1h_565_nl;
  wire[21:0] MultLoop_mux_117_nl;
  wire[21:0] MultLoop_mux_118_nl;
  wire[21:0] MultLoop_mux1h_566_nl;
  wire[21:0] MultLoop_acc_1667_nl;
  wire[22:0] nl_MultLoop_acc_1667_nl;
  wire[21:0] MultLoop_mux1h_567_nl;
  wire[21:0] MultLoop_mux1h_568_nl;
  wire[21:0] MultLoop_mux1h_569_nl;
  wire[21:0] MultLoop_mux1h_570_nl;
  wire[21:0] MultLoop_mux1h_571_nl;
  wire[21:0] MultLoop_mux1h_572_nl;
  wire[21:0] MultLoop_mux1h_573_nl;
  wire[21:0] MultLoop_mux1h_574_nl;
  wire[21:0] MultLoop_mux1h_575_nl;
  wire[21:0] MultLoop_mux1h_576_nl;
  wire[21:0] MultLoop_acc_1668_nl;
  wire[22:0] nl_MultLoop_acc_1668_nl;
  wire[21:0] MultLoop_acc_1669_nl;
  wire[22:0] nl_MultLoop_acc_1669_nl;
  wire[21:0] MultLoop_mux1h_577_nl;
  wire[21:0] MultLoop_acc_1670_nl;
  wire[22:0] nl_MultLoop_acc_1670_nl;
  wire[21:0] MultLoop_mux1h_578_nl;
  wire[21:0] MultLoop_acc_1671_nl;
  wire[22:0] nl_MultLoop_acc_1671_nl;
  wire[21:0] MultLoop_acc_1672_nl;
  wire[22:0] nl_MultLoop_acc_1672_nl;
  wire[21:0] MultLoop_acc_1673_nl;
  wire[22:0] nl_MultLoop_acc_1673_nl;
  wire[21:0] MultLoop_mux1h_579_nl;
  wire[21:0] AccumDotWidth_mux1h_1439_nl;
  wire[21:0] MultLoop_acc_1674_nl;
  wire[22:0] nl_MultLoop_acc_1674_nl;
  wire[21:0] MultLoop_acc_1675_nl;
  wire[22:0] nl_MultLoop_acc_1675_nl;
  wire[21:0] AccumDotWidth_mux1h_1440_nl;
  wire[21:0] AccumDotWidth_mux1h_1441_nl;
  wire[21:0] AccumDotWidth_mux1h_1442_nl;
  wire[21:0] AccumDotWidth_mux1h_1443_nl;
  wire[21:0] AccumDotWidth_mux1h_1444_nl;
  wire[21:0] AccumDotWidth_mux1h_1445_nl;
  wire[21:0] AccumDotWidth_mux1h_1446_nl;
  wire[21:0] MultLoop_mux_119_nl;
  wire[21:0] MultLoop_mux_120_nl;
  wire[21:0] MultLoop_mux1h_580_nl;
  wire[21:0] MultLoop_mux1h_581_nl;
  wire[21:0] MultLoop_mux_121_nl;
  wire[21:0] MultLoop_mux_122_nl;
  wire[21:0] MultLoop_mux1h_582_nl;
  wire[21:0] MultLoop_acc_1676_nl;
  wire[22:0] nl_MultLoop_acc_1676_nl;
  wire[21:0] MultLoop_acc_1677_nl;
  wire[22:0] nl_MultLoop_acc_1677_nl;
  wire[21:0] MultLoop_mux1h_583_nl;
  wire[21:0] MultLoop_mux_123_nl;
  wire[21:0] MultLoop_acc_1678_nl;
  wire[22:0] nl_MultLoop_acc_1678_nl;
  wire[21:0] MultLoop_acc_1679_nl;
  wire[22:0] nl_MultLoop_acc_1679_nl;
  wire[21:0] MultLoop_acc_1680_nl;
  wire[22:0] nl_MultLoop_acc_1680_nl;
  wire[21:0] MultLoop_mux_124_nl;
  wire[21:0] AccumDotWidth_mux1h_1447_nl;
  wire[21:0] AccumDotWidth_acc_2720_nl;
  wire[23:0] nl_AccumDotWidth_acc_2720_nl;
  wire[21:0] AccumDotWidth_acc_2722_nl;
  wire[23:0] nl_AccumDotWidth_acc_2722_nl;
  wire[21:0] AccumDotWidth_mux1h_1448_nl;
  wire[21:0] MultLoop_mux1h_584_nl;
  wire[21:0] MultLoop_acc_1681_nl;
  wire[22:0] nl_MultLoop_acc_1681_nl;
  wire[21:0] MultLoop_acc_1682_nl;
  wire[22:0] nl_MultLoop_acc_1682_nl;
  wire[21:0] MultLoop_acc_1683_nl;
  wire[22:0] nl_MultLoop_acc_1683_nl;
  wire[21:0] MultLoop_mux1h_585_nl;
  wire[21:0] MultLoop_acc_1684_nl;
  wire[22:0] nl_MultLoop_acc_1684_nl;
  wire[21:0] MultLoop_acc_1685_nl;
  wire[22:0] nl_MultLoop_acc_1685_nl;
  wire[21:0] MultLoop_acc_1686_nl;
  wire[22:0] nl_MultLoop_acc_1686_nl;
  wire[21:0] MultLoop_mux1h_586_nl;
  wire[21:0] MultLoop_mux1h_587_nl;
  wire[21:0] AccumDotWidth_mux1h_1449_nl;
  wire[21:0] AccumDotWidth_mux1h_1450_nl;
  wire[21:0] AccumDotWidth_mux1h_1451_nl;
  wire[21:0] AccumDotWidth_acc_2725_nl;
  wire[22:0] nl_AccumDotWidth_acc_2725_nl;
  wire[21:0] AccumDotWidth_mux1h_1452_nl;
  wire[21:0] AccumDotWidth_mux1h_1453_nl;
  wire[21:0] AccumDotWidth_mux1h_1454_nl;
  wire[21:0] AccumDotWidth_mux1h_1455_nl;
  wire[21:0] AccumDotWidth_mux1h_1456_nl;
  wire[21:0] AccumDotWidth_mux1h_1457_nl;
  wire[21:0] AccumDotWidth_mux1h_1458_nl;
  wire[21:0] AccumDotWidth_mux1h_1459_nl;
  wire[21:0] AccumDotWidth_mux1h_1460_nl;
  wire[29:0] mul_272_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_923_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_924_nl;
  wire[29:0] mul_273_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_925_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_926_nl;
  wire[29:0] mul_274_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_927_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_928_nl;
  wire[29:0] mul_275_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_929_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_930_nl;
  wire[29:0] mul_276_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_931_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_932_nl;
  wire[29:0] mul_277_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_933_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_934_nl;
  wire[29:0] mul_278_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_935_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_936_nl;
  wire[29:0] mul_279_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_937_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_938_nl;
  wire[29:0] mul_280_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_939_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_940_nl;
  wire[29:0] mul_281_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_941_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_942_nl;
  wire[29:0] mul_282_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_943_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_944_nl;
  wire[29:0] mul_283_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_945_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_946_nl;
  wire[29:0] mul_284_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_947_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_948_nl;
  wire[29:0] mul_285_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_949_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_950_nl;
  wire[29:0] mul_286_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_951_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_952_nl;
  wire[29:0] mul_287_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_953_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_954_nl;
  wire[29:0] mul_288_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_955_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_956_nl;
  wire[29:0] mul_289_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_957_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_958_nl;
  wire[29:0] mul_290_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_959_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_960_nl;
  wire[29:0] mul_291_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_961_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_962_nl;
  wire[29:0] mul_292_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_963_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_964_nl;
  wire[29:0] mul_293_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_965_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_966_nl;
  wire[29:0] mul_294_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_967_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_40_nl;
  wire[29:0] mul_295_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_968_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_969_nl;
  wire[29:0] mul_296_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_970_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_971_nl;
  wire[29:0] mul_297_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_972_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_973_nl;
  wire[29:0] mul_298_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_974_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_975_nl;
  wire[29:0] mul_299_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_976_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_977_nl;
  wire[29:0] mul_300_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_978_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_979_nl;
  wire[29:0] mul_301_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_980_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_981_nl;
  wire[29:0] mul_302_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_982_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_983_nl;
  wire[29:0] mul_303_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_984_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_985_nl;
  wire[29:0] mul_304_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_986_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_987_nl;
  wire[29:0] mul_305_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_988_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_989_nl;
  wire[29:0] mul_306_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_990_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_991_nl;
  wire[29:0] mul_307_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_992_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_993_nl;
  wire[29:0] mul_308_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_994_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_995_nl;
  wire[29:0] mul_309_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_996_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_997_nl;
  wire[29:0] mul_310_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_998_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_999_nl;
  wire[29:0] mul_311_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1000_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1001_nl;
  wire[29:0] mul_312_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1002_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1003_nl;
  wire[29:0] mul_313_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1004_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1005_nl;
  wire[29:0] mul_314_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1006_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1007_nl;
  wire[29:0] mul_315_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1008_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1009_nl;
  wire[29:0] mul_316_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1010_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1011_nl;
  wire[29:0] mul_317_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1012_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1013_nl;
  wire[29:0] mul_318_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1014_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1015_nl;
  wire[29:0] mul_319_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1016_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1017_nl;
  wire[29:0] mul_320_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1018_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_41_nl;
  wire[29:0] mul_321_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1019_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1020_nl;
  wire[29:0] mul_322_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1021_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1022_nl;
  wire[29:0] mul_323_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1023_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_42_nl;
  wire[29:0] mul_324_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1024_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1025_nl;
  wire[29:0] mul_325_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1026_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1027_nl;
  wire[29:0] mul_326_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1028_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_43_nl;
  wire[29:0] mul_327_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1029_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1030_nl;
  wire[29:0] mul_328_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1031_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1032_nl;
  wire[29:0] mul_329_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1033_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1034_nl;
  wire[29:0] mul_330_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1035_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1036_nl;
  wire[29:0] mul_331_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1037_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1038_nl;
  wire[29:0] mul_332_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1039_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1040_nl;
  wire[29:0] mul_333_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1041_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1042_nl;
  wire[29:0] mul_334_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1043_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1044_nl;
  wire[29:0] mul_335_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1045_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1046_nl;
  wire[29:0] mul_336_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1047_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_44_nl;
  wire[29:0] mul_337_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1048_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1049_nl;
  wire[29:0] mul_338_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1050_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1051_nl;
  wire[29:0] mul_339_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1052_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1053_nl;
  wire[29:0] mul_340_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1054_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1055_nl;
  wire[29:0] mul_341_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1056_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1057_nl;
  wire[29:0] mul_342_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1058_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1059_nl;
  wire[29:0] mul_343_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1060_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1061_nl;
  wire[29:0] mul_344_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1062_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1063_nl;
  wire[29:0] mul_345_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1064_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1065_nl;
  wire[29:0] mul_346_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1066_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1067_nl;
  wire[29:0] mul_347_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1068_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1069_nl;
  wire[29:0] mul_348_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1070_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1071_nl;
  wire[29:0] mul_349_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1072_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_45_nl;
  wire[29:0] mul_350_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1073_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1074_nl;
  wire[29:0] mul_351_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1075_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1076_nl;
  wire[29:0] mul_352_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1077_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1078_nl;
  wire[29:0] mul_353_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1079_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_46_nl;
  wire[29:0] mul_354_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1080_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1081_nl;
  wire[29:0] mul_355_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1082_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1083_nl;
  wire[29:0] mul_356_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1084_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1085_nl;
  wire[29:0] mul_357_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1086_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_47_nl;
  wire[29:0] mul_358_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1087_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1088_nl;
  wire[29:0] mul_359_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1089_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1090_nl;
  wire[0:0] ConvFiltWidth_else_or_931_nl;
  wire[29:0] mul_360_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1091_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1092_nl;
  wire[29:0] mul_361_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1093_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1094_nl;
  wire[29:0] mul_362_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1095_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1096_nl;
  wire[29:0] mul_363_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1097_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1098_nl;
  wire[29:0] mul_364_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1099_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1100_nl;
  wire[29:0] mul_365_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1101_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1102_nl;
  wire[29:0] mul_366_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1103_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1104_nl;
  wire[29:0] mul_367_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1105_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1106_nl;
  wire[29:0] mul_368_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1107_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1108_nl;
  wire[29:0] mul_369_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1109_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1110_nl;
  wire[29:0] mul_370_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1111_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1112_nl;
  wire[29:0] mul_371_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1113_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1114_nl;
  wire[29:0] mul_372_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1115_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1116_nl;
  wire[29:0] mul_373_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1117_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1118_nl;
  wire[29:0] mul_374_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1119_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1120_nl;
  wire[29:0] mul_375_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1121_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1122_nl;
  wire[29:0] mul_376_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1123_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1124_nl;
  wire[29:0] mul_377_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1125_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1126_nl;
  wire[29:0] mul_378_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1127_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1128_nl;
  wire[29:0] mul_379_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1129_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1130_nl;
  wire[29:0] mul_380_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1131_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1132_nl;
  wire[29:0] mul_381_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1133_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1134_nl;
  wire[29:0] mul_382_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1135_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1136_nl;
  wire[29:0] mul_383_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1137_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1138_nl;
  wire[29:0] mul_384_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1139_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1140_nl;
  wire[29:0] mul_385_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1141_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_48_nl;
  wire[29:0] mul_386_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1142_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_49_nl;
  wire[29:0] mul_387_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1143_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1144_nl;
  wire[29:0] mul_388_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1145_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1146_nl;
  wire[29:0] mul_389_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1147_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1148_nl;
  wire[29:0] mul_390_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1149_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1150_nl;
  wire[29:0] mul_391_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1151_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1152_nl;
  wire[29:0] mul_392_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1153_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1154_nl;
  wire[29:0] mul_393_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1155_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1156_nl;
  wire[29:0] mul_394_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1157_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_50_nl;
  wire[29:0] mul_395_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1158_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1159_nl;
  wire[29:0] mul_396_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1160_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_51_nl;
  wire[29:0] mul_397_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1161_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1162_nl;
  wire[0:0] ConvFiltWidth_else_or_989_nl;
  wire[29:0] mul_398_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1163_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1164_nl;
  wire[29:0] mul_399_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1165_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1166_nl;
  wire[29:0] mul_400_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1167_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1168_nl;
  wire[29:0] mul_401_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1169_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1170_nl;
  wire[29:0] mul_402_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1171_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1172_nl;
  wire[29:0] mul_403_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1173_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1174_nl;
  wire[29:0] mul_404_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1175_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1176_nl;
  wire[29:0] mul_405_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1177_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1178_nl;
  wire[29:0] mul_406_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1179_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1180_nl;
  wire[29:0] mul_407_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1181_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1182_nl;
  wire[29:0] mul_408_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1183_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1184_nl;
  wire[29:0] mul_409_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1185_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1186_nl;
  wire[29:0] mul_410_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1187_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1188_nl;
  wire[29:0] mul_411_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1189_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1190_nl;
  wire[29:0] mul_412_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1191_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_52_nl;
  wire[29:0] mul_413_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1192_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1193_nl;
  wire[29:0] mul_414_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1194_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1195_nl;
  wire[29:0] mul_415_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1196_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1197_nl;
  wire[29:0] mul_416_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1198_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1199_nl;
  wire[29:0] mul_417_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1200_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1201_nl;
  wire[29:0] mul_418_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1202_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1203_nl;
  wire[29:0] mul_419_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1204_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1205_nl;
  wire[29:0] mul_420_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1206_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1207_nl;
  wire[29:0] mul_421_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1208_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1209_nl;
  wire[29:0] mul_422_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1210_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1211_nl;
  wire[29:0] mul_423_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1212_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1213_nl;
  wire[29:0] mul_424_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1214_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1215_nl;
  wire[29:0] mul_425_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1216_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_53_nl;
  wire[29:0] mul_426_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1217_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_54_nl;
  wire[29:0] mul_427_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1218_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1219_nl;
  wire[29:0] mul_428_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1220_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1221_nl;
  wire[29:0] mul_429_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1222_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1223_nl;
  wire[29:0] mul_430_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1224_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1225_nl;
  wire[29:0] mul_431_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1226_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1227_nl;
  wire[29:0] mul_432_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1228_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1229_nl;
  wire[29:0] mul_433_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1230_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1231_nl;
  wire[29:0] mul_434_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1232_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1233_nl;
  wire[29:0] mul_435_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1234_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1235_nl;
  wire[29:0] mul_436_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1236_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1237_nl;
  wire[29:0] mul_437_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1238_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1239_nl;
  wire[29:0] mul_438_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1240_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1241_nl;
  wire[29:0] mul_439_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1242_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1243_nl;
  wire[29:0] mul_440_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1244_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1245_nl;
  wire[29:0] mul_441_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1246_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1247_nl;
  wire[29:0] mul_442_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1248_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1249_nl;
  wire[29:0] mul_443_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1250_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1251_nl;
  wire[29:0] mul_444_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1252_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1253_nl;
  wire[29:0] mul_445_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1254_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1255_nl;
  wire[29:0] mul_446_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1256_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1257_nl;
  wire[29:0] mul_447_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1258_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_55_nl;
  wire[29:0] mul_448_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1259_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1260_nl;
  wire[29:0] mul_449_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1261_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1262_nl;
  wire[29:0] mul_450_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1263_nl;
  wire[29:0] mul_451_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1264_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_56_nl;
  wire[29:0] mul_452_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1265_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_57_nl;
  wire[29:0] mul_453_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1266_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1267_nl;
  wire[29:0] mul_454_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1268_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1269_nl;
  wire[29:0] mul_455_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1270_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1271_nl;
  wire[29:0] mul_456_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1272_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1273_nl;
  wire[29:0] mul_457_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1274_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1275_nl;
  wire[29:0] mul_458_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1276_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1277_nl;
  wire[29:0] mul_459_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1278_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1279_nl;
  wire[29:0] mul_460_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1280_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1281_nl;
  wire[29:0] mul_461_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1282_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1283_nl;
  wire[29:0] mul_462_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1284_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1285_nl;
  wire[29:0] mul_463_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1286_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1287_nl;
  wire[29:0] mul_464_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1288_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1289_nl;
  wire[29:0] mul_465_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1290_nl;
  wire[29:0] mul_466_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1291_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1292_nl;
  wire[29:0] mul_467_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1293_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1294_nl;
  wire[29:0] mul_468_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1295_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1296_nl;
  wire[29:0] mul_469_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1297_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1298_nl;
  wire[29:0] mul_470_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1299_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1300_nl;
  wire[29:0] mul_471_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1301_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1302_nl;
  wire[29:0] mul_472_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1303_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_58_nl;
  wire[29:0] mul_473_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1304_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1305_nl;
  wire[29:0] mul_474_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1306_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1307_nl;
  wire[29:0] mul_475_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1308_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1309_nl;
  wire[29:0] mul_476_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1310_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_59_nl;
  wire[29:0] mul_477_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1311_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1312_nl;
  wire[29:0] mul_478_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1313_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_60_nl;
  wire[29:0] mul_479_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1314_nl;
  wire[29:0] mul_480_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1315_nl;
  wire[29:0] mul_481_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1316_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1317_nl;
  wire[29:0] mul_482_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1318_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1319_nl;
  wire[29:0] mul_483_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1320_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1321_nl;
  wire[29:0] mul_484_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1322_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1323_nl;
  wire[29:0] mul_485_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1324_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_61_nl;
  wire[29:0] mul_486_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1325_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_62_nl;
  wire[29:0] mul_487_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1326_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1327_nl;
  wire[29:0] mul_488_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1328_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1329_nl;
  wire[29:0] mul_489_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1330_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1331_nl;
  wire[29:0] mul_490_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1332_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1333_nl;
  wire[29:0] mul_491_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1334_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1335_nl;
  wire[29:0] mul_492_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1336_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1337_nl;
  wire[29:0] mul_493_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1338_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1339_nl;
  wire[29:0] mul_494_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1340_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1341_nl;
  wire[29:0] mul_495_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1342_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1343_nl;
  wire[29:0] mul_496_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1344_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1345_nl;
  wire[29:0] mul_497_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1346_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1347_nl;
  wire[29:0] mul_498_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1348_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1349_nl;
  wire[29:0] mul_499_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1350_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1351_nl;
  wire[29:0] mul_500_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1352_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1353_nl;
  wire[29:0] mul_501_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1354_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1355_nl;
  wire[29:0] mul_502_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1356_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1357_nl;
  wire[29:0] mul_503_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1358_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1359_nl;
  wire[29:0] mul_504_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1360_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_63_nl;
  wire[29:0] mul_505_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1361_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1362_nl;
  wire[29:0] mul_506_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1363_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_64_nl;
  wire[29:0] mul_507_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1364_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1365_nl;
  wire[29:0] mul_508_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1366_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1367_nl;
  wire[29:0] mul_509_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1368_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1369_nl;
  wire[29:0] mul_510_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1370_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1371_nl;
  wire[29:0] mul_511_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1372_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1373_nl;
  wire[29:0] mul_512_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1374_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1375_nl;
  wire[29:0] mul_513_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1376_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1377_nl;
  wire[29:0] mul_514_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1378_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1379_nl;
  wire[0:0] ConvFiltWidth_else_or_1166_nl;
  wire[29:0] mul_515_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1380_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1381_nl;
  wire[29:0] mul_516_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1382_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1383_nl;
  wire[29:0] mul_517_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1384_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1385_nl;
  wire[29:0] mul_518_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1386_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1387_nl;
  wire[29:0] mul_519_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1388_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1389_nl;
  wire[29:0] mul_520_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1390_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1391_nl;
  wire[29:0] mul_521_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1392_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_65_nl;
  wire[29:0] mul_522_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1393_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1394_nl;
  wire[29:0] mul_523_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1395_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1396_nl;
  wire[29:0] mul_524_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1397_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1398_nl;
  wire[29:0] mul_525_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1399_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1400_nl;
  wire[29:0] mul_526_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1401_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1402_nl;
  wire[29:0] mul_527_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1403_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1404_nl;
  wire[29:0] mul_528_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1405_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1406_nl;
  wire[29:0] mul_529_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1407_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1408_nl;
  wire[29:0] mul_530_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1409_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1410_nl;
  wire[29:0] mul_531_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1411_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1412_nl;
  wire[29:0] mul_532_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1413_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1414_nl;
  wire[29:0] mul_533_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1415_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1416_nl;
  wire[29:0] mul_534_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1417_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1418_nl;
  wire[29:0] mul_535_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1419_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1420_nl;
  wire[29:0] mul_536_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1421_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1422_nl;
  wire[29:0] mul_537_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1423_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1424_nl;
  wire[29:0] mul_538_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1425_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1426_nl;
  wire[29:0] mul_539_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1427_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1428_nl;
  wire[29:0] mul_540_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1429_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1430_nl;
  wire[29:0] mul_541_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1431_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1432_nl;
  wire[29:0] mul_542_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1433_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1434_nl;
  wire[29:0] mul_543_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1435_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_66_nl;
  wire[29:0] mul_544_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1436_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_67_nl;
  wire[29:0] mul_545_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1437_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1438_nl;
  wire[29:0] mul_546_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1439_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1440_nl;
  wire[29:0] mul_547_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1441_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1442_nl;
  wire[29:0] mul_548_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1443_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1444_nl;
  wire[29:0] mul_549_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1445_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1446_nl;
  wire[29:0] mul_550_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1447_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1448_nl;
  wire[29:0] mul_551_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1449_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1450_nl;
  wire[29:0] mul_552_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1451_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1452_nl;
  wire[29:0] mul_553_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1453_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1454_nl;
  wire[29:0] mul_554_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1455_nl;
  wire[29:0] mul_555_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1456_nl;
  wire[29:0] mul_556_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1457_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1458_nl;
  wire[29:0] mul_557_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1459_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1460_nl;
  wire[29:0] mul_558_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1461_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1462_nl;
  wire[29:0] mul_559_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1463_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1464_nl;
  wire[29:0] mul_560_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1465_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1466_nl;
  wire[29:0] mul_561_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1467_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1468_nl;
  wire[29:0] mul_562_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1469_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1470_nl;
  wire[29:0] mul_563_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1471_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1472_nl;
  wire[29:0] mul_564_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1473_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1474_nl;
  wire[29:0] mul_565_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1475_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1476_nl;
  wire[29:0] mul_566_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1477_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1478_nl;
  wire[29:0] mul_567_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1479_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_68_nl;
  wire[29:0] mul_568_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1480_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_69_nl;
  wire[29:0] mul_569_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1481_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1482_nl;
  wire[29:0] mul_570_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1483_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1484_nl;
  wire[29:0] mul_571_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1485_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1486_nl;
  wire[29:0] mul_572_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1487_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1488_nl;
  wire[29:0] mul_573_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1489_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1490_nl;
  wire[29:0] mul_574_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1491_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1492_nl;
  wire[29:0] mul_575_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1493_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1494_nl;
  wire[29:0] mul_576_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1495_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_70_nl;
  wire[29:0] mul_577_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1496_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1497_nl;
  wire[29:0] mul_578_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1498_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1499_nl;
  wire[29:0] mul_579_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1500_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1501_nl;
  wire[29:0] mul_580_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1502_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1503_nl;
  wire[29:0] mul_581_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1504_nl;
  wire[21:0] ConvFiltWidth_else_ConvFiltWidth_else_mux_71_nl;
  wire[29:0] mul_582_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1505_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1506_nl;
  wire[29:0] mul_583_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1507_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1508_nl;
  wire[29:0] mul_584_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1509_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1510_nl;
  wire[29:0] mul_585_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1511_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1512_nl;
  wire[29:0] mul_586_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1513_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1514_nl;
  wire[29:0] mul_587_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1515_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1516_nl;
  wire[29:0] mul_588_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1517_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1518_nl;
  wire[29:0] mul_589_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1519_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1520_nl;
  wire[29:0] mul_590_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1521_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1522_nl;
  wire[29:0] mul_591_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1523_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1524_nl;
  wire[29:0] mul_592_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1525_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1526_nl;
  wire[29:0] mul_593_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1527_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1528_nl;
  wire[29:0] mul_594_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1529_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1530_nl;
  wire[29:0] mul_595_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1531_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1532_nl;
  wire[29:0] mul_596_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1533_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1534_nl;
  wire[29:0] mul_597_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1535_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1536_nl;
  wire[29:0] mul_598_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1537_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1538_nl;
  wire[29:0] mul_599_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1539_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1540_nl;
  wire[29:0] mul_600_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1541_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1542_nl;
  wire[29:0] mul_601_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1543_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1544_nl;
  wire[29:0] mul_602_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1545_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1546_nl;
  wire[29:0] mul_603_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1547_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1548_nl;
  wire[29:0] mul_604_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1549_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1550_nl;
  wire[29:0] mul_605_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1551_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1552_nl;
  wire[29:0] mul_606_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1553_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1554_nl;
  wire[29:0] mul_607_nl;
  wire[7:0] ConvFiltWidth_else_mux1h_1555_nl;
  wire[21:0] ConvFiltWidth_else_mux1h_1556_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [219:0] nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat;
  assign nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat = {1'b0 ,
      layer5_out_rsci_idat_218_198 , 1'b0 , layer5_out_rsci_idat_196_176 , 1'b0 ,
      layer5_out_rsci_idat_174_154 , 1'b0 , layer5_out_rsci_idat_152_132 , 1'b0 ,
      layer5_out_rsci_idat_130_110 , 1'b0 , layer5_out_rsci_idat_108_88 , 1'b0 ,
      layer5_out_rsci_idat_86_66 , 1'b0 , layer5_out_rsci_idat_64_44 , 1'b0 , layer5_out_rsci_idat_42_22
      , 1'b0 , layer5_out_rsci_idat_20_0};
  econ_4x4_d10_core_input_1_rsci econ_4x4_d10_core_input_1_rsci_inst (
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .input_1_rsci_idat_mxwt(input_1_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_layer5_out_rsci econ_4x4_d10_core_layer5_out_rsci_inst (
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .core_wten(core_wten),
      .layer5_out_rsci_iswt0(reg_layer5_out_rsc_triosy_obj_ld_core_psct_cse),
      .layer5_out_rsci_idat(nl_econ_4x4_d10_core_layer5_out_rsci_inst_layer5_out_rsci_idat[219:0])
    );
  econ_4x4_d10_core_const_size_in_1_rsci econ_4x4_d10_core_const_size_in_1_rsci_inst
      (
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_in_1_rsci_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_out_1_rsci econ_4x4_d10_core_const_size_out_1_rsci_inst
      (
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .core_wten(core_wten),
      .const_size_out_1_rsci_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w2_rsci econ_4x4_d10_core_w2_rsci_inst (
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .w2_rsci_idat_mxwt(w2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b2_rsci econ_4x4_d10_core_b2_rsci_inst (
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .b2_rsci_idat_mxwt(b2_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_w4_rsci econ_4x4_d10_core_w4_rsci_inst (
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .w4_rsci_idat_mxwt(w4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_b4_rsci econ_4x4_d10_core_b4_rsci_inst (
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsci_oswt(reg_b4_rsc_triosy_obj_ld_core_psct_cse),
      .b4_rsci_wen_comp(b4_rsci_wen_comp),
      .b4_rsci_idat_mxwt(b4_rsci_idat_mxwt)
    );
  econ_4x4_d10_core_input_1_rsc_triosy_obj econ_4x4_d10_core_input_1_rsc_triosy_obj_inst
      (
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .input_1_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_layer5_out_rsc_triosy_obj econ_4x4_d10_core_layer5_out_rsc_triosy_obj_inst
      (
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .core_wten(core_wten),
      .layer5_out_rsc_triosy_obj_iswt0(reg_layer5_out_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj econ_4x4_d10_core_const_size_in_1_rsc_triosy_obj_inst
      (
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_in_1_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj econ_4x4_d10_core_const_size_out_1_rsc_triosy_obj_inst
      (
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .core_wten(core_wten),
      .const_size_out_1_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w2_rsc_triosy_obj econ_4x4_d10_core_w2_rsc_triosy_obj_inst (
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .core_wten(core_wten),
      .w2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b2_rsc_triosy_obj econ_4x4_d10_core_b2_rsc_triosy_obj_inst (
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .core_wten(core_wten),
      .b2_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_w4_rsc_triosy_obj econ_4x4_d10_core_w4_rsc_triosy_obj_inst (
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .core_wten(core_wten),
      .w4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_b4_rsc_triosy_obj econ_4x4_d10_core_b4_rsc_triosy_obj_inst (
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz),
      .core_wten(core_wten),
      .b4_rsc_triosy_obj_iswt0(reg_b4_rsc_triosy_obj_ld_core_psct_cse)
    );
  econ_4x4_d10_core_staller econ_4x4_d10_core_staller_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .input_1_rsci_wen_comp(input_1_rsci_wen_comp),
      .w2_rsci_wen_comp(w2_rsci_wen_comp),
      .b2_rsci_wen_comp(b2_rsci_wen_comp),
      .w4_rsci_wen_comp(w4_rsci_wen_comp),
      .b4_rsci_wen_comp(b4_rsci_wen_comp)
    );
  econ_4x4_d10_core_core_fsm econ_4x4_d10_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign layer5_out_and_cse = core_wen & (fsm_output[8]);
  assign InitAccum_and_cse = core_wen & (fsm_output[1]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_cse = core_wen & ((fsm_output[1])
      | (fsm_output[2]) | (fsm_output[7]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse = (fsm_output[3])
      | (fsm_output[1]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_1_cse = core_wen & nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse;
  assign MultLoop_and_1_cse = core_wen & ((fsm_output[5:1]!=5'b00000));
  assign MultLoop_and_2_cse = core_wen & ((fsm_output[6:1]!=6'b000000));
  assign MultLoop_or_46_cse = (fsm_output[4:3]!=2'b00);
  assign AccumDotWidth_and_3_cse = core_wen & ((fsm_output[1]) | (fsm_output[2])
      | (fsm_output[4]));
  assign AccumDotWidth_and_5_cse = core_wen & ((fsm_output[5]) | (fsm_output[2])
      | (fsm_output[1]));
  assign AccumDotWidth_and_7_cse = core_wen & ((fsm_output[4:1]!=4'b0000));
  assign MultLoop_and_4_cse = core_wen & ((fsm_output[2:1]!=2'b00));
  assign AccumDotWidth_and_8_cse = core_wen & ((fsm_output[1]) | (fsm_output[2])
      | (fsm_output[4]) | (fsm_output[5]));
  assign AccumDotWidth_and_10_cse = core_wen & ((fsm_output[3:1]!=3'b000));
  assign MultLoop_and_11_cse = core_wen & ((fsm_output[1]) | (fsm_output[2]) | (fsm_output[4])
      | (fsm_output[5]) | (fsm_output[6]));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_10_cse = core_wen &
      (fsm_output[2]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse = (fsm_output[2])
      | (fsm_output[7]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_29_cse = core_wen
      & nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse;
  assign AccumDotWidth_or_25_cse = (fsm_output[3:2]!=2'b00);
  assign AccumDotWidth_and_25_cse = core_wen & AccumDotWidth_or_25_cse;
  assign AccumDotWidth_or_26_cse = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[6]);
  assign AccumDotWidth_and_26_cse = core_wen & AccumDotWidth_or_26_cse;
  assign AccumDotWidth_or_38_cse = (fsm_output[5:4]!=2'b00);
  assign AccumDotWidth_or_29_cse = (fsm_output[4:2]!=3'b000);
  assign MultLoop_or_17_cse = (fsm_output[5:2]!=4'b0000);
  assign MultLoop_and_35_cse = core_wen & MultLoop_or_17_cse;
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_11_cse = core_wen &
      (fsm_output[3]);
  assign MultLoop_or_22_cse = (fsm_output[7]) | (fsm_output[3]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse = (fsm_output[5:3]!=3'b000);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_32_cse = core_wen
      & nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse;
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse = (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_34_cse = core_wen
      & nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse;
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_31_cse = core_wen &
      (fsm_output[4]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_47_cse = core_wen &
      (fsm_output[5]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_59_cse = core_wen &
      (fsm_output[6]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_267[20:0]), z_out_8_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_227[20:0]), z_out_12_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_271[20:0]), z_out_15_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_228[20:0]), z_out_16_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_838[20:0]), z_out_17_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_847[20:0]), z_out_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_835[20:0]), z_out_4_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_844[20:0]), z_out_10_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_825[20:0]), z_out_11_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_269[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_756[20:0]), z_out_15_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_270[20:0]), z_out_5_22);
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(z_out_476);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_476[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_12_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_265[20:0]), z_out_9_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_538[20:0]), z_out_10_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_453[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_534[20:0]), z_out_14_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_456[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_535[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_454[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_756[20:0]), z_out_18_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_459[20:0]), z_out_3_22);
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(z_out_751);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_751[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_17_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_456[20:0]), z_out_10_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_228[20:0]), z_out_9_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_271[20:0]), z_out_11_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_267[20:0]), z_out_12_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_751[20:0]), z_out_21_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_759[20:0]), z_out_24_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_825[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_474[20:0]), z_out_8_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_466[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_270[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_756[20:0]), z_out_17_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_538[20:0]), z_out_4_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_474[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_537[20:0]), z_out_8_22);
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(z_out_759);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_759[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_18_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_755[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_533[20:0]), z_out_3_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_542[20:0]), z_out_12_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_472[20:0]), z_out_4_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_809[20:0]), z_out_4_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_563[20:0]), z_out_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_566[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_564[20:0]), z_out_8_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_565[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_812[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_813[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_475[20:0]), z_out_22_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_471[20:0]), z_out_23_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_813[20:0]), z_out_24_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_265[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_472[20:0]), z_out_22);
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(z_out_752);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_752[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_19_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_811[20:0]), z_out_13_22);
  assign nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      =  -conv_s2s_22_23(z_out_818);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl
      = nl_nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_818[20:0]), (readslicef_23_1_22((nnet_relu_layer2_t_layer3_t_relu_config3_for_21_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl))));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_271[20:0]), z_out_9_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_275[20:0]), z_out_15_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_847[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_835[20:0]), z_out_11_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_824[20:0]), z_out_12_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_825[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_836[20:0]), z_out_3_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_831[20:0]), z_out_16_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_837[20:0]), z_out_4_22);
  assign nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[2047:2040]));
  assign MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7
      = readslicef_29_22_7((MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl));
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_534[20:0]), z_out_15_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_535[20:0]), z_out_11_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_518[20:0]), z_out_10_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_530[20:0]), z_out_9_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_808[20:0]), z_out_18_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_809[20:0]), z_out_13_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_811[20:0]), z_out_22_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_759[20:0]), z_out_14_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_752[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_751[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_762[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_813[20:0]), z_out_16_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_815[20:0]), z_out_23_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_812[20:0]), z_out_24_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_470[20:0]), z_out_3_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_475[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_476[20:0]), z_out_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_534[20:0]), z_out_11_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_530[20:0]), z_out_15_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_538[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_535[20:0]), z_out_8_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_466[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_533[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_530[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_535[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_812[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_mx0w0
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_813[20:0]), z_out_8_22);
  assign nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = z_out_466 + z_out_762;
  assign AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1
      = nl_AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = z_out_823 + z_out_534;
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[21:0];
  assign nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = z_out_809 + z_out_518;
  assign nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1 = nl_nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[21:0];
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_812[20:0]), z_out_13_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_809[20:0]), z_out_23_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_535[20:0]), z_out_17_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_530[20:0]), z_out_8_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_534[20:0]), z_out_7_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_533[20:0]), z_out_6_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_475[20:0]), z_out_5_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_474[20:0]), z_out_3_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_466[20:0]), z_out_2_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_453[20:0]), z_out_1_22);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_454[20:0]), z_out_22);
  assign or_tmp_4503 = (fsm_output[2]) | (fsm_output[5]) | (fsm_output[6]);
  assign nl_MultLoop_acc_162_sdt = (z_out_1129_29_7[21:0]) + (z_out_1128_29_7[21:0]);
  assign MultLoop_acc_162_sdt = nl_MultLoop_acc_162_sdt[21:0];
  assign nl_MultLoop_acc_27_sdt = (z_out_996_29_7[21:0]) + (z_out_995_29_7[21:0]);
  assign MultLoop_acc_27_sdt = nl_MultLoop_acc_27_sdt[21:0];
  assign nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[383:376]));
  assign MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[391:384]));
  assign MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1193_sdt = (readslicef_29_22_7((MultLoop_48_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_49_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1193_sdt = nl_MultLoop_acc_1193_sdt[21:0];
  assign nl_MultLoop_acc_1201_sdt = z_out_188_28_7 + z_out_163_28_7;
  assign MultLoop_acc_1201_sdt = nl_MultLoop_acc_1201_sdt[21:0];
  assign nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[463:456]));
  assign MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[471:464]));
  assign MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1188_sdt = (readslicef_29_22_7((MultLoop_58_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_59_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1188_sdt = nl_MultLoop_acc_1188_sdt[21:0];
  assign nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[511:504]));
  assign MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[519:512]));
  assign MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl
      = nl_MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl[28:0];
  assign nl_MultLoop_acc_1185_sdt = (readslicef_29_22_7((MultLoop_64_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)))
      + (readslicef_29_22_7((MultLoop_65_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_nl)));
  assign MultLoop_acc_1185_sdt = nl_MultLoop_acc_1185_sdt[21:0];
  assign AccumDotWidth_or_132_cse_1 = (fsm_output[1]) | (fsm_output[4]);
  always @(posedge clk) begin
    if ( rst ) begin
      layer5_out_rsci_idat_218_198 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_42_22 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_64_44 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_86_66 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_108_88 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_130_110 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_152_132 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_174_154 <= 21'b000000000000000000000;
      layer5_out_rsci_idat_196_176 <= 21'b000000000000000000000;
    end
    else if ( layer5_out_and_cse ) begin
      layer5_out_rsci_idat_218_198 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_288[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_20_0 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_214[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_42_22 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_303[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_64_44 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_298[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_86_66 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_292[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_108_88 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_290[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_130_110 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_289[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
      layer5_out_rsci_idat_152_132 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_213[20:0]),
          z_out_19_22);
      layer5_out_rsci_idat_174_154 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_215[20:0]),
          z_out_20_22);
      layer5_out_rsci_idat_196_176 <= MUX_v_21_2_2(21'b000000000000000000000, (z_out_216[20:0]),
          (readslicef_23_1_22((nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl))));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      reg_layer5_out_rsc_triosy_obj_ld_core_psct_cse <= 1'b0;
      MultLoop_acc_1000_itm <= 22'b0000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      AccumDotWidth_acc_1274_itm <= 22'b0000000000000000000000;
      MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      MultLoop_acc_1284_psp <= 11'b00000000000;
      MultLoop_acc_1283_psp <= 11'b00000000000;
      MultLoop_acc_1282_psp <= 11'b00000000000;
      MultLoop_acc_1281_psp <= 11'b00000000000;
      MultLoop_acc_1280_psp <= 11'b00000000000;
    end
    else if ( core_wen ) begin
      reg_b4_rsc_triosy_obj_ld_core_psct_cse <= (fsm_output[9]) | (fsm_output[0]);
      reg_layer5_out_rsc_triosy_obj_ld_core_psct_cse <= fsm_output[8];
      MultLoop_acc_1000_itm <= MUX1HOT_v_22_5_2(z_out_779, z_out_768, z_out_800,
          z_out_789, z_out_788, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[5]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_935_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_1117_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_874_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_605_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_611_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_607_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      AccumDotWidth_acc_1274_itm <= MUX1HOT_v_22_5_2(z_out_721, z_out_762, z_out_782,
          z_out_474, z_out_779, {(fsm_output[2]) , (fsm_output[3]) , AccumDotWidth_or_38_cse
          , (fsm_output[6]) , (fsm_output[7])});
      MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_4_2(z_out_132_28_7, z_out_143_28_7, z_out_772, z_out_796,
          {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
      MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_4_2(z_out_139_28_7, z_out_135_28_7, z_out_61_28_7, z_out_185_28_7,
          {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1;
      MultLoop_acc_1284_psp <= nl_MultLoop_acc_1284_psp[10:0];
      MultLoop_acc_1283_psp <= nl_MultLoop_acc_1283_psp[10:0];
      MultLoop_acc_1282_psp <= nl_MultLoop_acc_1282_psp[10:0];
      MultLoop_acc_1281_psp <= nl_MultLoop_acc_1281_psp[10:0];
      MultLoop_acc_1280_psp <= nl_MultLoop_acc_1280_psp[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      InitAccum_io_read_b4_rsc_cse_sva <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
      MultLoop_io_read_w4_rsc_cse_sva <= {640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 640'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
      ConvFiltWidth_else_io_read_input_1_rsc_cse_sva <= {528'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 528'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
      ConvFiltWidth_else_io_read_w2_rsc_cse_sva <= {864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
          , 864'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
      nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva <=
          64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( InitAccum_and_cse ) begin
      InitAccum_io_read_b4_rsc_cse_sva <= b4_rsci_idat_mxwt;
      MultLoop_io_read_w4_rsc_cse_sva <= w4_rsci_idat_mxwt;
      ConvFiltWidth_else_io_read_input_1_rsc_cse_sva <= input_1_rsci_idat_mxwt;
      ConvFiltWidth_else_io_read_w2_rsc_cse_sva <= w2_rsci_idat_mxwt;
      nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva <=
          b2_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      AccumDotWidth_acc_1916_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1135_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          (z_out_994_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      AccumDotWidth_acc_1916_itm <= MUX1HOT_v_22_3_2(z_out_680, z_out_424, ({1'b0
          , nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0}),
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
      AccumDotWidth_acc_1135_itm <= MUX1HOT_v_22_3_2(z_out_752, z_out_766, z_out_65_28_7,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_1_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_181_itm <= 22'b0000000000000000000000;
      MultLoop_acc_243_itm <= 22'b0000000000000000000000;
    end
    else if ( MultLoop_and_1_cse ) begin
      MultLoop_acc_181_itm <= MUX1HOT_v_22_5_2(z_out_767, z_out_466, z_out_768, z_out_769,
          z_out_770, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
          , (fsm_output[5])});
      MultLoop_acc_243_itm <= MUX1HOT_v_22_5_2(z_out_781, z_out_471, z_out_753, z_out_796,
          z_out_785, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
          , (fsm_output[5])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_308_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1007_itm <= 22'b0000000000000000000000;
      MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
    end
    else if ( MultLoop_and_2_cse ) begin
      MultLoop_acc_308_itm <= MUX1HOT_v_22_5_2(z_out_771, z_out_772, z_out_773, z_out_753,
          z_out_290, {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5])
          , (fsm_output[6])});
      MultLoop_acc_1007_itm <= MUX1HOT_v_22_6_2(z_out_772, z_out_472, z_out_769,
          z_out_783, z_out_819, z_out_779, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
      MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_6_2(z_out_768, z_out_476, z_out_138_28_7, z_out_140_28_7,
          z_out_774, z_out_771, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1133_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & ((fsm_output[6]) | (fsm_output[2]) | (fsm_output[1])) )
        begin
      AccumDotWidth_acc_1133_itm <= MUX1HOT_v_22_3_2(z_out_812, z_out_534, z_out_177_28_7,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1164_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1326_itm <= 22'b0000000000000000000000;
      MultLoop_acc_105_itm <= 22'b0000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= 21'b000000000000000000000;
    end
    else if ( AccumDotWidth_and_3_cse ) begin
      AccumDotWidth_acc_1164_itm <= MUX1HOT_v_22_3_2(z_out_809, z_out_816, z_out_767,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
      AccumDotWidth_acc_1326_itm <= MUX1HOT_v_22_3_2(z_out_811, z_out_747, z_out_139_28_7,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
      MultLoop_acc_105_itm <= MUX1HOT_v_22_3_2(z_out_783, z_out_811, z_out_766, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[4])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2(z_out_978_29_9, (z_out_1119_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2((z_out_976_29_7[22:2]), (z_out_931_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1167_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & ((fsm_output[1]) | (fsm_output[2]) | (fsm_output[5]) | (fsm_output[6]))
        ) begin
      AccumDotWidth_acc_1167_itm <= MUX1HOT_v_22_4_2(z_out_474, z_out_475, z_out_776,
          z_out_777, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1169_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1181_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1184_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1186_itm <= 22'b0000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= 21'b000000000000000000000;
    end
    else if ( AccumDotWidth_and_5_cse ) begin
      AccumDotWidth_acc_1169_itm <= MUX1HOT_v_22_3_2(z_out_756, z_out_769, z_out_779,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
      AccumDotWidth_acc_1181_itm <= MUX1HOT_v_22_3_2(z_out_813, z_out_815, z_out_809,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
      AccumDotWidth_acc_1184_itm <= MUX1HOT_v_22_3_2(z_out_808, z_out_818, z_out_281,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
      AccumDotWidth_acc_1186_itm <= MUX1HOT_v_22_3_2(z_out_815, z_out_775, z_out_283,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2((z_out_974_29_7[22:2]), (z_out_1118_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2((z_out_970_29_7[22:2]), (z_out_933_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1201_itm <= 22'b0000000000000000000000;
      MultLoop_acc_229_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1203_itm <= 22'b0000000000000000000000;
      ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
    end
    else if ( AccumDotWidth_and_7_cse ) begin
      AccumDotWidth_acc_1201_itm <= MUX1HOT_v_22_4_2(z_out_751, z_out_470, z_out_815,
          z_out_779, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      MultLoop_acc_229_itm <= MUX1HOT_v_22_4_2(z_out_774, z_out_773, z_out_770, z_out_440,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      AccumDotWidth_acc_1203_itm <= MUX1HOT_v_22_4_2(z_out_466, z_out_781, z_out_689,
          z_out_757, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_4_2((z_out_969_29_7[22:2]), (z_out_1120_29_7[22:2]), (z_out_1021_29_7[22:2]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_slc_29_9_itm
          <= MUX1HOT_v_21_4_2((z_out_973_29_7[22:2]), (z_out_1121_29_7[22:2]), (z_out_1130_29_7[22:2]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_4_2((z_out_971_29_7[22:2]), (z_out_1110_29_7[22:2]), (z_out_618_29_7[22:2]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= MUX1HOT_v_21_4_2((z_out_968_29_7[22:2]), (z_out_896_29_7[22:2]), z_out_978_29_9,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_4_2(z_out_979_29_9, (z_out_929_29_7[22:2]), (z_out_1174_29_7[22:2]),
          nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_102_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & ((fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
        | (fsm_output[7])) ) begin
      MultLoop_acc_102_itm <= MUX1HOT_v_22_4_2(z_out_776, z_out_473, z_out_781, z_out_783,
          {nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse , (fsm_output[2])
          , (fsm_output[4]) , (fsm_output[7])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_1095_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1012_itm <= 22'b0000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm
          <= 21'b000000000000000000000;
    end
    else if ( MultLoop_and_4_cse ) begin
      MultLoop_acc_1095_itm <= MUX_v_22_2_2(z_out_770, z_out_786, fsm_output[2]);
      MultLoop_acc_1012_itm <= MUX_v_22_2_2(z_out_788, z_out_223, fsm_output[2]);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm
          <= MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
          nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
          fsm_output[2]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1300_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1010_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1018_itm <= 22'b0000000000000000000000;
    end
    else if ( AccumDotWidth_and_8_cse ) begin
      AccumDotWidth_acc_1300_itm <= MUX1HOT_v_22_4_2(z_out_467, z_out_382, z_out_816,
          z_out_761, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_1010_itm <= MUX1HOT_v_22_4_2(z_out_790, z_out_484, z_out_775,
          z_out_824, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_1018_itm <= MUX1HOT_v_22_4_2(z_out_782, z_out_774, z_out_798,
          z_out_783, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1352_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1218_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1220_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1235_itm <= 22'b0000000000000000000000;
      MultLoop_acc_215_itm <= 22'b0000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= 21'b000000000000000000000;
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= 21'b000000000000000000000;
    end
    else if ( AccumDotWidth_and_10_cse ) begin
      AccumDotWidth_acc_1352_itm <= MUX1HOT_v_22_3_2(z_out_816, z_out_741, z_out_771,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      AccumDotWidth_acc_1218_itm <= MUX1HOT_v_22_3_2(z_out_759, z_out_820, z_out_796,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      AccumDotWidth_acc_1220_itm <= MUX1HOT_v_22_3_2(z_out_472, z_out_765, z_out_215,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      AccumDotWidth_acc_1235_itm <= MUX1HOT_v_22_3_2(z_out_755, z_out_823, z_out_779,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      MultLoop_acc_215_itm <= MUX1HOT_v_22_3_2(z_out_796, z_out_808, z_out_772, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[3])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_609_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
          (z_out_617_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2((z_out_972_29_7[22:2]), (z_out_1112_29_7[22:2]), nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm
          <= MUX1HOT_v_21_3_2((z_out_1041_29_7[22:2]), (z_out_936_29_7[22:2]), (nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_nl),
          {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_1089_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1121_itm <= 22'b0000000000000000000000;
      MultLoop_acc_113_itm <= 22'b0000000000000000000000;
    end
    else if ( MultLoop_and_11_cse ) begin
      MultLoop_acc_1089_itm <= MUX1HOT_v_22_5_2(z_out_785, z_out_762, z_out_787,
          z_out_775, z_out_200, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[5]) , (fsm_output[6])});
      MultLoop_acc_1121_itm <= MUX1HOT_v_22_5_2(z_out_775, z_out_481, z_out_785,
          z_out_790, z_out_796, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])
          , (fsm_output[5]) , (fsm_output[6])});
      MultLoop_acc_113_itm <= MUX1HOT_v_22_5_2(z_out_787, z_out_469, z_out_789, z_out_781,
          z_out_767, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_128_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & ((fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
        | (fsm_output[6])) ) begin
      MultLoop_acc_128_itm <= MUX1HOT_v_22_5_2(z_out_789, z_out_474, z_out_765, z_out_803,
          z_out_783, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
          , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_1222_itm <= 22'b0000000000000000000000;
      MultLoop_acc_1266_itm <= 22'b0000000000000000000000;
      MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_1139_itm <= 22'b0000000000000000000000;
      MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_841_itm <= 22'b0000000000000000000000;
      MultLoop_acc_885_itm <= 22'b0000000000000000000000;
      MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_714_itm <= 22'b0000000000000000000000;
      MultLoop_acc_758_itm <= 22'b0000000000000000000000;
      MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_587_itm <= 22'b0000000000000000000000;
      MultLoop_acc_631_itm <= 22'b0000000000000000000000;
      MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_460_itm <= 22'b0000000000000000000000;
      MultLoop_acc_504_itm <= 22'b0000000000000000000000;
      MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_333_itm <= 22'b0000000000000000000000;
      MultLoop_acc_377_itm <= 22'b0000000000000000000000;
      MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_206_itm <= 22'b0000000000000000000000;
      MultLoop_acc_250_itm <= 22'b0000000000000000000000;
      MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_79_itm <= 22'b0000000000000000000000;
      MultLoop_acc_123_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_10_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_144_28_7;
      MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_143_28_7;
      MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_72_28_7;
      MultLoop_acc_1222_itm <= z_out_213;
      MultLoop_acc_1266_itm <= z_out_783;
      MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_139_28_7;
      MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_136_28_7;
      MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_71_28_7;
      MultLoop_acc_1139_itm <= z_out_231;
      MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_135_28_7;
      MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_68_28_7;
      MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_67_28_7;
      MultLoop_acc_841_itm <= z_out_214;
      MultLoop_acc_885_itm <= z_out_292;
      MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_129_28_7;
      MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_66_28_7;
      MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_65_28_7;
      MultLoop_acc_714_itm <= z_out_788;
      MultLoop_acc_758_itm <= z_out_288;
      MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_133_28_7;
      MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_64_28_7;
      MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_63_28_7;
      MultLoop_acc_587_itm <= z_out_767;
      MultLoop_acc_631_itm <= z_out_796;
      MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_130_28_7;
      MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_62_28_7;
      MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_61_28_7;
      MultLoop_acc_460_itm <= z_out_777;
      MultLoop_acc_504_itm <= z_out_212;
      MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_118_28_7;
      MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_69_28_7;
      MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_70_28_7;
      MultLoop_acc_333_itm <= z_out_771;
      MultLoop_acc_377_itm <= z_out_289;
      MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_122_28_7;
      MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_140_28_7;
      MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_138_28_7;
      MultLoop_acc_206_itm <= z_out_215;
      MultLoop_acc_250_itm <= z_out_290;
      MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_134_28_7;
      MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_142_28_7;
      MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_121_28_7;
      MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= z_out_73_28_7;
      MultLoop_acc_79_itm <= z_out_216;
      MultLoop_acc_123_itm <= z_out_779;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_968_itm <= 22'b0000000000000000000000;
      MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1932_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1937_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1945_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1877_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1871_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1837_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1845_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1426_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_29_cse )
        begin
      MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX_v_22_2_2(z_out_76_28_7, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      MultLoop_acc_968_itm <= MUX_v_22_2_2(z_out_776, z_out_767, fsm_output[7]);
      MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX_v_22_2_2(z_out_75_28_7, z_out_121_28_7, fsm_output[7]);
      MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX_v_22_2_2(z_out_77_28_7, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      AccumDotWidth_acc_1932_itm <= MUX_v_22_2_2(z_out_712, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      AccumDotWidth_acc_1937_itm <= MUX_v_22_2_2(z_out_364, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      AccumDotWidth_acc_1945_itm <= MUX_v_22_2_2(z_out_822, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      AccumDotWidth_acc_1877_itm <= MUX_v_22_2_2(z_out_542, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0}),
          fsm_output[7]);
      AccumDotWidth_acc_1871_itm <= MUX_v_22_2_2(z_out_360, ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1}),
          fsm_output[7]);
      AccumDotWidth_acc_1837_itm <= MUX_v_22_2_2(z_out_357, z_out_64_28_7, fsm_output[7]);
      AccumDotWidth_acc_1845_itm <= MUX_v_22_2_2(z_out_821, z_out_63_28_7, fsm_output[7]);
      AccumDotWidth_acc_1426_itm <= MUX_v_22_2_2(z_out_795, z_out_62_28_7, fsm_output[7]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1392_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1397_itm <= 22'b0000000000000000000000;
      AccumDotWidth_acc_1371_itm <= 22'b0000000000000000000000;
    end
    else if ( AccumDotWidth_and_25_cse ) begin
      AccumDotWidth_acc_1392_itm <= MUX_v_22_2_2(z_out_538, z_out_214, fsm_output[3]);
      AccumDotWidth_acc_1397_itm <= MUX_v_22_2_2(z_out_535, z_out_767, fsm_output[3]);
      AccumDotWidth_acc_1371_itm <= MUX_v_22_2_2(z_out_536, z_out_216, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1378_itm <= 22'b0000000000000000000000;
      MultLoop_acc_372_itm <= 22'b0000000000000000000000;
    end
    else if ( AccumDotWidth_and_26_cse ) begin
      AccumDotWidth_acc_1378_itm <= MUX1HOT_v_22_4_2(z_out_358, z_out_682, z_out_770,
          z_out_772, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
      MultLoop_acc_372_itm <= MUX1HOT_v_22_4_2(z_out_518, z_out_800, z_out_774, z_out_776,
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      AccumDotWidth_acc_1198_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & AccumDotWidth_or_29_cse ) begin
      AccumDotWidth_acc_1198_itm <= MUX1HOT_v_22_3_2(z_out_524, z_out_808, z_out_784,
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_435_itm <= 22'b0000000000000000000000;
      MultLoop_acc_356_itm <= 22'b0000000000000000000000;
      MultLoop_acc_483_itm <= 22'b0000000000000000000000;
    end
    else if ( MultLoop_and_35_cse ) begin
      MultLoop_acc_435_itm <= MUX1HOT_v_22_4_2(z_out_784, z_out_757, z_out_761, z_out_787,
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_356_itm <= MUX1HOT_v_22_4_2(z_out_540, z_out_774, z_out_792, z_out_765,
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_483_itm <= MUX1HOT_v_22_4_2(z_out_770, z_out_775, z_out_790, z_out_784,
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_36_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & ((fsm_output[2]) | (fsm_output[3]) | (fsm_output[6])) )
        begin
      MultLoop_acc_36_itm <= MUX1HOT_v_22_3_2(z_out_782, z_out_781, z_out_788, {(fsm_output[2])
          , (fsm_output[3]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      MultLoop_acc_629_itm <= 22'b0000000000000000000000;
      MultLoop_acc_597_itm <= 22'b0000000000000000000000;
      MultLoop_acc_596_itm <= 22'b0000000000000000000000;
      MultLoop_acc_502_itm <= 22'b0000000000000000000000;
      MultLoop_acc_470_itm <= 22'b0000000000000000000000;
      MultLoop_acc_89_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_11_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_809[20:0]), z_out_19_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_820[20:0]), z_out_20_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      MultLoop_acc_629_itm <= z_out_783;
      MultLoop_acc_597_itm <= z_out_231;
      MultLoop_acc_596_itm <= z_out_213;
      MultLoop_acc_502_itm <= z_out_788;
      MultLoop_acc_470_itm <= z_out_223;
      MultLoop_acc_89_itm <= z_out_212;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_acc_88_itm <= 22'b0000000000000000000000;
    end
    else if ( core_wen & MultLoop_or_22_cse ) begin
      MultLoop_acc_88_itm <= MUX_v_22_2_2(z_out_786, MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7,
          fsm_output[7]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_54_itm <= 22'b0000000000000000000000;
      MultLoop_acc_562_itm <= 22'b0000000000000000000000;
      MultLoop_acc_689_itm <= 22'b0000000000000000000000;
      MultLoop_acc_628_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_32_cse )
        begin
      MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_3_2(z_out_126_28_7, z_out_125_28_7, z_out_278, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_3_2(z_out_125_28_7, z_out_134_28_7, z_out_286, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_54_itm <= MUX1HOT_v_22_3_2(z_out_798, z_out_768, z_out_771, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_562_itm <= MUX1HOT_v_22_3_2(z_out_803, z_out_753, z_out_767, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_689_itm <= MUX1HOT_v_22_3_2(z_out_761, z_out_765, z_out_796, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
      MultLoop_acc_628_itm <= MUX1HOT_v_22_3_2(z_out_766, z_out_776, z_out_788, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[5])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= 22'b0000000000000000000000;
      MultLoop_acc_499_itm <= 22'b0000000000000000000000;
      MultLoop_acc_626_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_product_layer3_t_config4_weight_t_config4_accum_t_and_34_cse )
        begin
      MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
          <= MUX1HOT_v_22_3_2(z_out_121_28_7, z_out_130_28_7, z_out_118_28_7, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[6])});
      MultLoop_acc_499_itm <= MUX1HOT_v_22_3_2(z_out_777, z_out_771, z_out_786, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[6])});
      MultLoop_acc_626_itm <= MUX1HOT_v_22_3_2(z_out_792, z_out_772, z_out_794, {(fsm_output[3])
          , (fsm_output[4]) , (fsm_output[6])});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      MultLoop_acc_867_itm <= 22'b0000000000000000000000;
      MultLoop_acc_883_itm <= 22'b0000000000000000000000;
      MultLoop_acc_740_itm <= 22'b0000000000000000000000;
      MultLoop_acc_756_itm <= 22'b0000000000000000000000;
      MultLoop_acc_724_itm <= 22'b0000000000000000000000;
      MultLoop_acc_613_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_31_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_818[20:0]), z_out_21_22);
      MultLoop_acc_867_itm <= z_out_777;
      MultLoop_acc_883_itm <= nl_MultLoop_acc_883_itm[21:0];
      MultLoop_acc_740_itm <= z_out_786;
      MultLoop_acc_756_itm <= z_out_280;
      MultLoop_acc_724_itm <= nl_MultLoop_acc_724_itm[21:0];
      MultLoop_acc_613_itm <= z_out_788;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      MultLoop_acc_994_itm <= 22'b0000000000000000000000;
      MultLoop_acc_861_itm <= 22'b0000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_47_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_812[20:0]), z_out_9_22);
      MultLoop_acc_994_itm <= z_out_757;
      MultLoop_acc_861_itm <= z_out_766;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm <=
          21'b000000000000000000000;
    end
    else if ( nnet_relu_layer2_t_layer3_t_relu_config3_for_if_and_59_cse ) begin
      nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_227[20:0]), z_out_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_228[20:0]), z_out_3_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_229[20:0]), z_out_10_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_445[20:0]), z_out_16_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1[20:0]),
          z_out_11_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1[20:0]),
          z_out_12_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_480[20:0]), z_out_15_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_476[20:0]), z_out_17_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_475[20:0]), z_out_21_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_206[20:0]), z_out_1_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (z_out_444[20:0]), z_out_2_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm <=
          MUX_v_21_2_2(21'b000000000000000000000, (AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1[20:0]),
          z_out_4_22);
      nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
      nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm <=
          nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_mx0w0;
    end
  end
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_288);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_10_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_214);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_1_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_303);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_2_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_298);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_3_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_292);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_4_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_290);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_5_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_289);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_6_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      =  -conv_s2s_22_23(z_out_216);
  assign nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl
      = nl_nnet_relu_layer4_t_result_t_relu_config5_for_9_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign nl_MultLoop_acc_1284_psp  = (z_out_63_28_7[21:11]) + conv_s2u_8_11(InitAccum_io_read_b4_rsc_cse_sva[47:40]);
  assign nl_MultLoop_acc_1283_psp  = (z_out_64_28_7[21:11]) + conv_s2u_8_11(InitAccum_io_read_b4_rsc_cse_sva[39:32]);
  assign nl_MultLoop_acc_1282_psp  = (z_out_62_28_7[21:11]) + conv_s2u_8_11(InitAccum_io_read_b4_rsc_cse_sva[31:24]);
  assign nl_MultLoop_acc_1281_psp  = (z_out_65_28_7[21:11]) + conv_s2u_8_11(InitAccum_io_read_b4_rsc_cse_sva[23:16]);
  assign nl_MultLoop_acc_1280_psp  = (MultLoop_256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_itm_28_7[21:11])
      + conv_s2u_8_11(InitAccum_io_read_b4_rsc_cse_sva[15:8]);
  assign nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_nl
      = MUX_v_21_2_2(21'b000000000000000000000, (z_out_755[20:0]), z_out_21_22);
  assign nl_MultLoop_acc_883_itm  = z_out_455 + z_out_448;
  assign nl_MultLoop_acc_724_itm  = z_out_827 + z_out_842;
  assign operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse = (fsm_output[2]) | (fsm_output[4]);
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_21_nl = MUX1HOT_v_22_6_2((~ z_out_227),
      (~ z_out_847), (~ z_out_563), (~ z_out_472), (~ z_out_476), (~ z_out_454),
      {(fsm_output[6]) , (fsm_output[1]) , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_21_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_nl[22:0];
  assign z_out_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_22_nl = MUX1HOT_v_22_7_2((~ z_out_206),
      (~ z_out_456), (~ z_out_270), (~ z_out_812), (~ z_out_265), (~ z_out_475),
      (~ z_out_453), {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_22_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl[22:0];
  assign z_out_1_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_1_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_23_nl = MUX1HOT_v_22_7_2((~ z_out_444),
      (~ z_out_454), (~ z_out_474), (~ z_out_755), (~ z_out_813), (~ z_out_847),
      (~ z_out_466), {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_23_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl[22:0];
  assign z_out_2_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_2_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_24_nl = MUX1HOT_v_22_6_2((~ z_out_228),
      (~ z_out_459), (~ z_out_533), (~ z_out_836), (~ z_out_470), (~ z_out_474),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_24_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl[22:0];
  assign z_out_3_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_3_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse = (fsm_output[5]) | (fsm_output[7]);
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_25_nl = MUX1HOT_v_22_6_2((~ AccumOutHeight_3_AccumOutWidth_3_AccumFilt_2_AccumDotWidth_acc_ncse_sva_1),
      (~ z_out_835), (~ z_out_538), (~ z_out_472), (~ z_out_809), (~ z_out_837),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[2]) , (fsm_output[3])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_25_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl[22:0];
  assign z_out_4_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_4_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_26_nl = MUX1HOT_v_22_7_2((~ z_out_270),
      (~ z_out_535), (~ z_out_825), (~ z_out_752), (~ z_out_466), (~ z_out_812),
      (~ z_out_475), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_26_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl[22:0];
  assign z_out_5_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_5_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_27_nl = MUX1HOT_v_22_7_2((~ z_out_453),
      (~ z_out_565), (~ z_out_825), (~ z_out_751), (~ z_out_538), (~ z_out_535),
      (~ z_out_533), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_27_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl[22:0];
  assign z_out_6_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_6_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_28_nl = MUX1HOT_v_22_7_2((~ z_out_269),
      (~ z_out_466), (~ z_out_566), (~ z_out_762), (~ z_out_533), (~ z_out_530),
      (~ z_out_534), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_28_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl[22:0];
  assign z_out_7_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_7_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_29_nl = MUX1HOT_v_22_7_2((~ z_out_267),
      (~ z_out_474), (~ z_out_537), (~ z_out_564), (~ z_out_535), (~ z_out_813),
      (~ z_out_530), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_29_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl[22:0];
  assign z_out_8_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_8_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_30_nl = MUX1HOT_v_22_5_2((~ z_out_812),
      (~ z_out_265), (~ z_out_228), (~ z_out_271), (~ z_out_530), {(fsm_output[5])
      , (fsm_output[1]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_30_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl[22:0];
  assign z_out_9_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_9_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_31_nl = MUX1HOT_v_22_5_2((~ z_out_229),
      (~ z_out_844), (~ z_out_538), (~ z_out_456), (~ z_out_518), {(fsm_output[6])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) , AccumDotWidth_or_38_cse});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_31_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl[22:0];
  assign z_out_10_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_10_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_32_nl = MUX1HOT_v_22_6_2((~ nnet_conv_2d_input_t_layer2_t_config2_acc_59_sva_1),
      (~ z_out_825), (~ z_out_271), (~ z_out_835), (~ z_out_535), (~ z_out_534),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_32_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl[22:0];
  assign z_out_11_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_11_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_33_nl = MUX1HOT_v_22_5_2((~ nnet_conv_2d_input_t_layer2_t_config2_acc_60_sva_1),
      (~ z_out_227), (~ z_out_267), (~ z_out_542), (~ z_out_824), {(fsm_output[6])
      , (fsm_output[1]) , (fsm_output[7]) , AccumDotWidth_or_38_cse , (fsm_output[3])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_33_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl[22:0];
  assign z_out_12_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_12_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_34_nl = MUX1HOT_v_22_3_2((~ z_out_811),
      (~ z_out_809), (~ z_out_812), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_34_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl[22:0];
  assign z_out_13_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_13_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux_2_nl = MUX_v_22_2_2((~ z_out_534),
      (~ z_out_759), fsm_output[4]);
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux_2_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl[22:0];
  assign z_out_14_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_14_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_35_nl = MUX1HOT_v_22_6_2((~ z_out_480),
      (~ z_out_271), (~ z_out_756), (~ z_out_275), (~ z_out_534), (~ z_out_530),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_35_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl[22:0];
  assign z_out_15_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_15_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse = (fsm_output[4]) | (fsm_output[7]);
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_36_nl = MUX1HOT_v_22_4_2((~ z_out_445),
      (~ z_out_228), (~ z_out_831), (~ z_out_813), {(fsm_output[6]) , (fsm_output[1])
      , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_36_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl[22:0];
  assign z_out_16_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_16_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_37_nl = MUX1HOT_v_22_4_2((~ z_out_476),
      (~ z_out_838), (~ z_out_756), (~ z_out_535), {(fsm_output[6]) , nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse
      , (fsm_output[4]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_37_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl[22:0];
  assign z_out_17_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_17_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux_3_nl = MUX_v_22_2_2((~ z_out_756),
      (~ z_out_808), fsm_output[4]);
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux_3_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl[22:0];
  assign z_out_18_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_18_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_1_mux_2_nl = MUX_v_22_2_2((~ z_out_213),
      (~ z_out_809), fsm_output[3]);
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_1_mux_2_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl[22:0];
  assign z_out_19_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_1_acc_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_1_mux_3_nl = MUX_v_22_2_2((~ z_out_215),
      (~ z_out_820), fsm_output[3]);
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_1_mux_3_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl[22:0];
  assign z_out_20_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_1_acc_1_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_38_nl = MUX1HOT_v_22_4_2((~ z_out_755),
      (~ z_out_818), (~ z_out_475), (~ z_out_751), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_38_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl[22:0];
  assign z_out_21_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_19_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_operator_22_4_true_AC_TRN_AC_WRAP_mux_1_nl
      = MUX_v_22_2_2((~ z_out_475), (~ z_out_811), operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse);
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_operator_22_4_true_AC_TRN_AC_WRAP_mux_1_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl[22:0];
  assign z_out_22_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_20_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_39_nl = MUX1HOT_v_22_3_2((~ z_out_471),
      (~ z_out_815), (~ z_out_809), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[7])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_39_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl[22:0];
  assign z_out_23_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_21_nl));
  assign operator_22_4_true_AC_TRN_AC_WRAP_mux1h_40_nl = MUX1HOT_v_22_3_2((~ z_out_759),
      (~ z_out_813), (~ z_out_812), {(fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl = conv_s2u_22_23(operator_22_4_true_AC_TRN_AC_WRAP_mux1h_40_nl)
      + 23'b00000000000000000000001;
  assign operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl = nl_operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl[22:0];
  assign z_out_24_22 = readslicef_23_1_22((operator_22_4_true_AC_TRN_AC_WRAP_acc_22_nl));
  assign AccumDotWidth_mux1h_752_nl = MUX1HOT_v_10_3_2((z_out_628_29_7[22:13]), (nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm[20:11]),
      (z_out_627_29_7[22:13]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign AccumDotWidth_mux1h_753_nl = MUX1HOT_v_8_3_2((b2_rsci_idat_mxwt[55:48]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_25 = (AccumDotWidth_mux1h_752_nl) + conv_s2u_8_10(AccumDotWidth_mux1h_753_nl);
  assign z_out_25 = nl_z_out_25[9:0];
  assign AccumDotWidth_or_138_cse = (fsm_output[6:4]!=3'b000);
  assign AccumDotWidth_mux1h_755_nl = MUX1HOT_v_10_6_2((z_out_623_29_7[22:13]), (z_out_1033_29_9[20:11]),
      (z_out_1040_29_7[22:13]), (z_out_590_29_7[22:13]), (z_out_1108_29_7[22:13]),
      (z_out_1018_29_9[20:11]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_756_nl = MUX1HOT_v_8_3_2((b2_rsci_idat_mxwt[39:32]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]),
      {(fsm_output[1]) , MultLoop_or_22_cse , AccumDotWidth_or_138_cse});
  assign nl_z_out_27 = (AccumDotWidth_mux1h_755_nl) + conv_s2u_8_10(AccumDotWidth_mux1h_756_nl);
  assign z_out_27 = nl_z_out_27[9:0];
  assign AccumDotWidth_mux1h_757_nl = MUX1HOT_v_10_3_2((z_out_630_29_7[22:13]), (z_out_622_29_7[22:13]),
      (z_out_629_29_7[22:13]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign AccumDotWidth_mux1h_758_nl = MUX1HOT_v_8_3_2((b2_rsci_idat_mxwt[31:24]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_28 = (AccumDotWidth_mux1h_757_nl) + conv_s2u_8_10(AccumDotWidth_mux1h_758_nl);
  assign z_out_28 = nl_z_out_28[9:0];
  assign AccumDotWidth_or_140_cse = (fsm_output[7:6]!=2'b00);
  assign AccumDotWidth_or_139_cse = (fsm_output[3]) | (fsm_output[5]);
  assign AccumDotWidth_mux1h_759_nl = MUX1HOT_v_10_6_2((z_out_1156_29_7[22:13]),
      (z_out_1028_29_7[22:13]), (z_out_618_29_7[22:13]), (z_out_908_29_7[22:13]),
      (z_out_588_29_7[22:13]), (z_out_929_29_7[22:13]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_760_nl = MUX1HOT_v_8_4_2((b2_rsci_idat_mxwt[31:24]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , (fsm_output[4]) , AccumDotWidth_or_140_cse});
  assign nl_z_out_30 = (AccumDotWidth_mux1h_759_nl) + conv_s2u_8_10(AccumDotWidth_mux1h_760_nl);
  assign z_out_30 = nl_z_out_30[9:0];
  assign AccumDotWidth_mux_81_nl = MUX_v_10_2_2((nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm[20:11]),
      (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11]),
      fsm_output[5]);
  assign nl_z_out_31 = (AccumDotWidth_mux_81_nl) + conv_s2u_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign z_out_31 = nl_z_out_31[9:0];
  assign AccumDotWidth_AccumDotWidth_mux_18_nl = MUX_v_10_2_2((z_out_621_29_7[22:13]),
      (z_out_1133_29_9[20:11]), AccumDotWidth_or_140_cse);
  assign AccumDotWidth_AccumDotWidth_mux_19_nl = MUX_v_8_2_2((nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]),
      fsm_output[7]);
  assign nl_z_out_32 = (AccumDotWidth_AccumDotWidth_mux_18_nl) + conv_s2u_8_10(AccumDotWidth_AccumDotWidth_mux_19_nl);
  assign z_out_32 = nl_z_out_32[9:0];
  assign AccumDotWidth_or_142_cse = (fsm_output[7:5]!=3'b000);
  assign AccumDotWidth_mux1h_761_nl = MUX1HOT_v_10_4_2((z_out_628_29_7[22:13]), (z_out_989_29_9[20:11]),
      (z_out_609_29_7[22:13]), (z_out_883_29_7[22:13]), {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_AccumDotWidth_mux_20_nl = MUX_v_8_2_2((nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]),
      AccumDotWidth_or_142_cse);
  assign nl_z_out_33 = (AccumDotWidth_mux1h_761_nl) + conv_s2u_8_10(AccumDotWidth_AccumDotWidth_mux_20_nl);
  assign z_out_33 = nl_z_out_33[9:0];
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_332_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[6383:6376]),
      (w4_rsci_idat_mxwt[7095:7088]), (MultLoop_io_read_w4_rsc_cse_sva[4135:4128]),
      (MultLoop_io_read_w4_rsc_cse_sva[4471:4464]), (MultLoop_io_read_w4_rsc_cse_sva[6007:6000]),
      (MultLoop_io_read_w4_rsc_cse_sva[8967:8960]), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_333_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[2])
      , (fsm_output[7])});
  assign nl_mul_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_332_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_333_nl));
  assign mul_nl = nl_mul_nl[28:0];
  assign z_out_34_28_7 = readslicef_29_22_7((mul_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_334_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[3111:3104]),
      (w4_rsci_idat_mxwt[7087:7080]), (MultLoop_io_read_w4_rsc_cse_sva[5999:5992]),
      (MultLoop_io_read_w4_rsc_cse_sva[7543:7536]), (MultLoop_io_read_w4_rsc_cse_sva[8975:8968]),
      (MultLoop_io_read_w4_rsc_cse_sva[3247:3240]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_335_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[4])});
  assign nl_mul_1_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_334_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_335_nl));
  assign mul_1_nl = nl_mul_1_nl[28:0];
  assign z_out_35_28_7 = readslicef_29_22_7((mul_1_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_336_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1463:1456]),
      (w4_rsci_idat_mxwt[919:912]), (MultLoop_io_read_w4_rsc_cse_sva[4327:4320]),
      (MultLoop_io_read_w4_rsc_cse_sva[3103:3096]), (MultLoop_io_read_w4_rsc_cse_sva[5991:5984]),
      (MultLoop_io_read_w4_rsc_cse_sva[8999:8992]), {(fsm_output[5]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_337_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2])
      , (fsm_output[7])});
  assign nl_mul_2_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_336_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_337_nl));
  assign mul_2_nl = nl_mul_2_nl[28:0];
  assign z_out_36_28_7 = readslicef_29_22_7((mul_2_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_338_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[3991:3984]),
      (MultLoop_io_read_w4_rsc_cse_sva[4335:4328]), (MultLoop_io_read_w4_rsc_cse_sva[4455:4448]),
      (MultLoop_io_read_w4_rsc_cse_sva[3191:3184]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_339_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_3_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_338_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_339_nl));
  assign mul_3_nl = nl_mul_3_nl[28:0];
  assign z_out_37_28_7 = readslicef_29_22_7((mul_3_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_340_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[3999:3992]),
      (MultLoop_io_read_w4_rsc_cse_sva[2255:2248]), (MultLoop_io_read_w4_rsc_cse_sva[4447:4440]),
      (MultLoop_io_read_w4_rsc_cse_sva[1639:1632]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_341_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_4_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_340_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_341_nl));
  assign mul_4_nl = nl_mul_4_nl[28:0];
  assign z_out_38_28_7 = readslicef_29_22_7((mul_4_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_342_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[4007:4000]),
      (MultLoop_io_read_w4_rsc_cse_sva[2263:2256]), (MultLoop_io_read_w4_rsc_cse_sva[4439:4432]),
      (MultLoop_io_read_w4_rsc_cse_sva[1631:1624]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_343_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_5_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_342_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_343_nl));
  assign mul_5_nl = nl_mul_5_nl[28:0];
  assign z_out_39_28_7 = readslicef_29_22_7((mul_5_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_344_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[4015:4008]),
      (MultLoop_io_read_w4_rsc_cse_sva[2079:2072]), (MultLoop_io_read_w4_rsc_cse_sva[2279:2272]),
      (MultLoop_io_read_w4_rsc_cse_sva[2479:2472]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_345_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_6_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_344_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_345_nl));
  assign mul_6_nl = nl_mul_6_nl[28:0];
  assign z_out_40_28_7 = readslicef_29_22_7((mul_6_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_346_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[4023:4016]),
      (MultLoop_io_read_w4_rsc_cse_sva[2295:2288]), (MultLoop_io_read_w4_rsc_cse_sva[7535:7528]),
      (MultLoop_io_read_w4_rsc_cse_sva[4159:4152]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_347_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_7_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_346_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_347_nl));
  assign mul_7_nl = nl_mul_7_nl[28:0];
  assign z_out_41_28_7 = readslicef_29_22_7((mul_7_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_348_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[3311:3304]),
      (w4_rsci_idat_mxwt[7055:7048]), (MultLoop_io_read_w4_rsc_cse_sva[4463:4456]),
      (MultLoop_io_read_w4_rsc_cse_sva[5983:5976]), (MultLoop_io_read_w4_rsc_cse_sva[3175:3168]),
      (MultLoop_io_read_w4_rsc_cse_sva[9007:9000]), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_349_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[7])});
  assign nl_mul_8_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_348_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_349_nl));
  assign mul_8_nl = nl_mul_8_nl[28:0];
  assign z_out_42_28_7 = readslicef_29_22_7((mul_8_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_350_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[2087:2080]),
      (MultLoop_io_read_w4_rsc_cse_sva[5367:5360]), (w4_rsci_idat_mxwt[7047:7040]),
      (MultLoop_io_read_w4_rsc_cse_sva[2487:2480]), (MultLoop_io_read_w4_rsc_cse_sva[7031:7024]),
      (MultLoop_io_read_w4_rsc_cse_sva[9015:9008]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_351_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[2])
      , (fsm_output[7])});
  assign nl_mul_9_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_350_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_351_nl));
  assign mul_9_nl = nl_mul_9_nl[28:0];
  assign z_out_43_28_7 = readslicef_29_22_7((mul_9_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_352_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[3319:3312]),
      (MultLoop_io_read_w4_rsc_cse_sva[3447:3440]), (w4_rsci_idat_mxwt[7039:7032]),
      (MultLoop_io_read_w4_rsc_cse_sva[4127:4120]), (MultLoop_io_read_w4_rsc_cse_sva[7023:7016]),
      (MultLoop_io_read_w4_rsc_cse_sva[9023:9016]), {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_353_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[2])
      , (fsm_output[7])});
  assign nl_mul_10_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_352_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_353_nl));
  assign mul_10_nl = nl_mul_10_nl[28:0];
  assign z_out_44_28_7 = readslicef_29_22_7((mul_10_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_354_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[895:888]),
      (MultLoop_io_read_w4_rsc_cse_sva[5359:5352]), (MultLoop_io_read_w4_rsc_cse_sva[2471:2464]),
      (MultLoop_io_read_w4_rsc_cse_sva[7015:7008]), (MultLoop_io_read_w4_rsc_cse_sva[3143:3136]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_355_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_11_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_354_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_355_nl));
  assign mul_11_nl = nl_mul_11_nl[28:0];
  assign z_out_45_28_7 = readslicef_29_22_7((mul_11_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_356_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[6399:6392]),
      (MultLoop_io_read_w4_rsc_cse_sva[3183:3176]), (MultLoop_io_read_w4_rsc_cse_sva[3463:3456]),
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_357_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_12_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_356_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_357_nl));
  assign mul_12_nl = nl_mul_12_nl[28:0];
  assign z_out_46_28_7 = readslicef_29_22_7((mul_12_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_358_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2271:2264]),
      (MultLoop_io_read_w4_rsc_cse_sva[7007:7000]), (MultLoop_io_read_w4_rsc_cse_sva[3151:3144]),
      (MultLoop_io_read_w4_rsc_cse_sva[3487:3480]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_359_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_13_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_358_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_359_nl));
  assign mul_13_nl = nl_mul_13_nl[28:0];
  assign z_out_47_28_7 = readslicef_29_22_7((mul_13_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_360_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[903:896]),
      (MultLoop_io_read_w4_rsc_cse_sva[2303:2296]), (MultLoop_io_read_w4_rsc_cse_sva[2455:2448]),
      (MultLoop_io_read_w4_rsc_cse_sva[8055:8048]), (MultLoop_io_read_w4_rsc_cse_sva[3159:3152]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_361_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_14_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_360_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_361_nl));
  assign mul_14_nl = nl_mul_14_nl[28:0];
  assign z_out_48_28_7 = readslicef_29_22_7((mul_14_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_362_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[911:904]),
      (MultLoop_io_read_w4_rsc_cse_sva[1279:1272]), (MultLoop_io_read_w4_rsc_cse_sva[1095:1088]),
      (MultLoop_io_read_w4_rsc_cse_sva[2463:2456]), (MultLoop_io_read_w4_rsc_cse_sva[8047:8040]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[2])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_363_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[2])});
  assign nl_mul_15_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_362_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_363_nl));
  assign mul_15_nl = nl_mul_15_nl[28:0];
  assign z_out_49_28_7 = readslicef_29_22_7((mul_15_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_364_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1103:1096]),
      (MultLoop_io_read_w4_rsc_cse_sva[5351:5344]), (w4_rsci_idat_mxwt[7063:7056]),
      (MultLoop_io_read_w4_rsc_cse_sva[8039:8032]), (MultLoop_io_read_w4_rsc_cse_sva[7527:7520]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_365_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_16_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_364_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_365_nl));
  assign mul_16_nl = nl_mul_16_nl[28:0];
  assign z_out_50_28_7 = readslicef_29_22_7((mul_16_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_366_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1111:1104]),
      (MultLoop_io_read_w4_rsc_cse_sva[2287:2280]), (w4_rsci_idat_mxwt[7071:7064]),
      (MultLoop_io_read_w4_rsc_cse_sva[8031:8024]), (MultLoop_io_read_w4_rsc_cse_sva[7519:7512]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_367_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_17_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_366_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_367_nl));
  assign mul_17_nl = nl_mul_17_nl[28:0];
  assign z_out_51_28_7 = readslicef_29_22_7((mul_17_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_368_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1119:1112]),
      (MultLoop_io_read_w4_rsc_cse_sva[3303:3296]), (MultLoop_io_read_w4_rsc_cse_sva[4959:4952]),
      (MultLoop_io_read_w4_rsc_cse_sva[7511:7504]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_369_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_18_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_368_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_369_nl));
  assign mul_18_nl = nl_mul_18_nl[28:0];
  assign z_out_52_28_7 = readslicef_29_22_7((mul_18_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_370_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1127:1120]),
      (MultLoop_io_read_w4_rsc_cse_sva[6375:6368]), (MultLoop_io_read_w4_rsc_cse_sva[2447:2440]),
      (MultLoop_io_read_w4_rsc_cse_sva[4967:4960]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[2])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_371_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2])});
  assign nl_mul_19_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_370_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_371_nl));
  assign mul_19_nl = nl_mul_19_nl[28:0];
  assign z_out_53_28_7 = readslicef_29_22_7((mul_19_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_372_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2247:2240]),
      (MultLoop_io_read_w4_rsc_cse_sva[2439:2432]), (MultLoop_io_read_w4_rsc_cse_sva[4975:4968]),
      (MultLoop_io_read_w4_rsc_cse_sva[3167:3160]), {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_373_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_20_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_372_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_373_nl));
  assign mul_20_nl = nl_mul_20_nl[28:0];
  assign z_out_54_28_7 = readslicef_29_22_7((mul_20_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_374_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[927:920]),
      (MultLoop_io_read_w4_rsc_cse_sva[3455:3448]), (MultLoop_io_read_w4_rsc_cse_sva[4271:4264]),
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_375_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_21_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_374_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_375_nl));
  assign mul_21_nl = nl_mul_21_nl[28:0];
  assign z_out_55_28_7 = readslicef_29_22_7((mul_21_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_376_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[3287:3280]),
      (w4_rsci_idat_mxwt[7079:7072]), (MultLoop_io_read_w4_rsc_cse_sva[3479:3472]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_377_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_mul_22_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_376_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_377_nl));
  assign mul_22_nl = nl_mul_22_nl[28:0];
  assign z_out_56_28_7 = readslicef_29_22_7((mul_22_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_89_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[951:944]),
      (MultLoop_io_read_w4_rsc_cse_sva[3295:3288]), fsm_output[4]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_90_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      fsm_output[4]);
  assign nl_mul_23_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_89_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_90_nl));
  assign mul_23_nl = nl_mul_23_nl[28:0];
  assign z_out_57_28_7 = readslicef_29_22_7((mul_23_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_91_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[943:936]),
      (MultLoop_io_read_w4_rsc_cse_sva[6391:6384]), fsm_output[4]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_92_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[4]);
  assign nl_mul_24_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_91_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_92_nl));
  assign mul_24_nl = nl_mul_24_nl[28:0];
  assign z_out_58_28_7 = readslicef_29_22_7((mul_24_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_378_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[935:928]),
      (MultLoop_io_read_w4_rsc_cse_sva[4343:4336]), (MultLoop_io_read_w4_rsc_cse_sva[2431:2424]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_379_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_25_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_378_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_379_nl));
  assign mul_25_nl = nl_mul_25_nl[28:0];
  assign z_out_59_28_7 = readslicef_29_22_7((mul_25_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_380_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[3279:3272]),
      (w4_rsci_idat_mxwt[2999:2992]), (MultLoop_io_read_w4_rsc_cse_sva[3471:3464]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_381_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_mul_26_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_380_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_381_nl));
  assign mul_26_nl = nl_mul_26_nl[28:0];
  assign z_out_60_28_7 = readslicef_29_22_7((mul_26_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_382_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1159:1152]),
      (w4_rsci_idat_mxwt[4991:4984]), (MultLoop_io_read_w4_rsc_cse_sva[4895:4888]),
      (MultLoop_io_read_w4_rsc_cse_sva[8863:8856]), (MultLoop_io_read_w4_rsc_cse_sva[4407:4400]),
      (MultLoop_io_read_w4_rsc_cse_sva[6583:6576]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_383_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_mul_27_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_382_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_383_nl));
  assign mul_27_nl = nl_mul_27_nl[28:0];
  assign z_out_61_28_7 = readslicef_29_22_7((mul_27_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_384_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1167:1160]),
      (w4_rsci_idat_mxwt[3007:3000]), (MultLoop_io_read_w4_rsc_cse_sva[4887:4880]),
      (MultLoop_io_read_w4_rsc_cse_sva[4367:4360]), (MultLoop_io_read_w4_rsc_cse_sva[6575:6568]),
      (MultLoop_io_read_w4_rsc_cse_sva[4095:4088]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_385_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7])});
  assign nl_mul_28_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_384_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_385_nl));
  assign mul_28_nl = nl_mul_28_nl[28:0];
  assign z_out_62_28_7 = readslicef_29_22_7((mul_28_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_386_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[9167:9160]),
      (MultLoop_io_read_w4_rsc_cse_sva[5919:5912]), (MultLoop_io_read_w4_rsc_cse_sva[6455:6448]),
      (MultLoop_io_read_w4_rsc_cse_sva[4247:4240]), (MultLoop_io_read_w4_rsc_cse_sva[6567:6560]),
      (MultLoop_io_read_w4_rsc_cse_sva[6143:6136]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_387_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[7])});
  assign nl_mul_29_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_386_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_387_nl));
  assign mul_29_nl = nl_mul_29_nl[28:0];
  assign z_out_63_28_7 = readslicef_29_22_7((mul_29_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_388_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1175:1168]),
      (w4_rsci_idat_mxwt[5047:5040]), (MultLoop_io_read_w4_rsc_cse_sva[5911:5904]),
      (MultLoop_io_read_w4_rsc_cse_sva[4279:4272]), (MultLoop_io_read_w4_rsc_cse_sva[5511:5504]),
      (MultLoop_io_read_w4_rsc_cse_sva[5119:5112]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_389_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7])});
  assign nl_mul_30_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_388_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_389_nl));
  assign mul_30_nl = nl_mul_30_nl[28:0];
  assign z_out_64_28_7 = readslicef_29_22_7((mul_30_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_390_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[2175:2168]),
      (w4_rsci_idat_mxwt[5055:5048]), (MultLoop_io_read_w4_rsc_cse_sva[6943:6936]),
      (MultLoop_io_read_w4_rsc_cse_sva[6447:6440]), (MultLoop_io_read_w4_rsc_cse_sva[5527:5520]),
      (MultLoop_io_read_w4_rsc_cse_sva[3071:3064]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_391_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7])});
  assign nl_mul_31_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_390_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_391_nl));
  assign mul_31_nl = nl_mul_31_nl[28:0];
  assign z_out_65_28_7 = readslicef_29_22_7((mul_31_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_392_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[959:952]),
      (MultLoop_io_read_w4_rsc_cse_sva[6935:6928]), (MultLoop_io_read_w4_rsc_cse_sva[4239:4232]),
      (MultLoop_io_read_w4_rsc_cse_sva[3335:3328]), (MultLoop_io_read_w4_rsc_cse_sva[9039:9032]),
      (MultLoop_io_read_w4_rsc_cse_sva[5503:5496]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_393_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[5])});
  assign nl_mul_32_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_392_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_393_nl));
  assign mul_32_nl = nl_mul_32_nl[28:0];
  assign z_out_66_28_7 = readslicef_29_22_7((mul_32_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_394_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[6039:6032]),
      (MultLoop_io_read_w4_rsc_cse_sva[3263:3256]), (MultLoop_io_read_w4_rsc_cse_sva[7967:7960]),
      (MultLoop_io_read_w4_rsc_cse_sva[4223:4216]), (MultLoop_io_read_w4_rsc_cse_sva[9031:9024]),
      (MultLoop_io_read_w4_rsc_cse_sva[6559:6552]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_395_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[5])});
  assign nl_mul_33_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_394_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_395_nl));
  assign mul_33_nl = nl_mul_33_nl[28:0];
  assign z_out_67_28_7 = readslicef_29_22_7((mul_33_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_396_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[6023:6016]),
      (MultLoop_io_read_w4_rsc_cse_sva[7959:7952]), (MultLoop_io_read_w4_rsc_cse_sva[8959:8952]),
      (MultLoop_io_read_w4_rsc_cse_sva[3223:3216]), (MultLoop_io_read_w4_rsc_cse_sva[3255:3248]),
      (MultLoop_io_read_w4_rsc_cse_sva[6551:6544]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_397_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_mul_34_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_396_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_397_nl));
  assign mul_34_nl = nl_mul_34_nl[28:0];
  assign z_out_68_28_7 = readslicef_29_22_7((mul_34_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_398_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[6047:6040]),
      (MultLoop_io_read_w4_rsc_cse_sva[3863:3856]), (MultLoop_io_read_w4_rsc_cse_sva[6431:6424]),
      (MultLoop_io_read_w4_rsc_cse_sva[5159:5152]), (MultLoop_io_read_w4_rsc_cse_sva[4495:4488]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_399_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_35_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_398_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_399_nl));
  assign mul_35_nl = nl_mul_35_nl[28:0];
  assign z_out_69_28_7 = readslicef_29_22_7((mul_35_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_400_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[4031:4024]),
      (MultLoop_io_read_w4_rsc_cse_sva[3871:3864]), (MultLoop_io_read_w4_rsc_cse_sva[6415:6408]),
      (MultLoop_io_read_w4_rsc_cse_sva[4503:4496]), (MultLoop_io_read_w4_rsc_cse_sva[1063:1056]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_401_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_36_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_400_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_401_nl));
  assign mul_36_nl = nl_mul_36_nl[28:0];
  assign z_out_70_28_7 = readslicef_29_22_7((mul_36_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_402_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[6071:6064]),
      (MultLoop_io_read_w4_rsc_cse_sva[10071:10064]), (MultLoop_io_read_w4_rsc_cse_sva[7583:7576]),
      (MultLoop_io_read_w4_rsc_cse_sva[5423:5416]), (MultLoop_io_read_w4_rsc_cse_sva[1055:1048]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_403_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_37_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_402_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_403_nl));
  assign mul_37_nl = nl_mul_37_nl[28:0];
  assign z_out_71_28_7 = readslicef_29_22_7((mul_37_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_404_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[6031:6024]),
      (MultLoop_io_read_w4_rsc_cse_sva[855:848]), (MultLoop_io_read_w4_rsc_cse_sva[6407:6400]),
      (MultLoop_io_read_w4_rsc_cse_sva[7591:7584]), (MultLoop_io_read_w4_rsc_cse_sva[6183:6176]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_405_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_38_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_404_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_405_nl));
  assign mul_38_nl = nl_mul_38_nl[28:0];
  assign z_out_72_28_7 = readslicef_29_22_7((mul_38_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_406_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[6063:6056]),
      (MultLoop_io_read_w4_rsc_cse_sva[1879:1872]), (MultLoop_io_read_w4_rsc_cse_sva[4511:4504]),
      (MultLoop_io_read_w4_rsc_cse_sva[6175:6168]), (MultLoop_io_read_w4_rsc_cse_sva[5431:5424]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_407_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_39_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_406_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_407_nl));
  assign mul_39_nl = nl_mul_39_nl[28:0];
  assign z_out_73_28_7 = readslicef_29_22_7((mul_39_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_408_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[9175:9168]),
      (MultLoop_io_read_w4_rsc_cse_sva[4231:4224]), (MultLoop_io_read_w4_rsc_cse_sva[4519:4512]),
      (MultLoop_io_read_w4_rsc_cse_sva[4359:4352]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_409_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_40_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_408_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_409_nl));
  assign mul_40_nl = nl_mul_40_nl[28:0];
  assign z_out_74_28_7 = readslicef_29_22_7((mul_40_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_410_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[6055:6048]),
      (MultLoop_io_read_w4_rsc_cse_sva[8983:8976]), (MultLoop_io_read_w4_rsc_cse_sva[6423:6416]),
      (MultLoop_io_read_w4_rsc_cse_sva[5151:5144]), (MultLoop_io_read_w4_rsc_cse_sva[4535:4528]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_411_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_41_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_410_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_411_nl));
  assign mul_41_nl = nl_mul_41_nl[28:0];
  assign z_out_75_28_7 = readslicef_29_22_7((mul_41_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_412_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[8087:8080]),
      (MultLoop_io_read_w4_rsc_cse_sva[9047:9040]), (MultLoop_io_read_w4_rsc_cse_sva[5447:5440]),
      (MultLoop_io_read_w4_rsc_cse_sva[5519:5512]), (MultLoop_io_read_w4_rsc_cse_sva[6207:6200]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_413_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_42_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_412_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_413_nl));
  assign mul_42_nl = nl_mul_42_nl[28:0];
  assign z_out_76_28_7 = readslicef_29_22_7((mul_42_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_414_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1151:1144]),
      (MultLoop_io_read_w4_rsc_cse_sva[1207:1200]), (w4_rsci_idat_mxwt[5071:5064]),
      (MultLoop_io_read_w4_rsc_cse_sva[8991:8984]), (MultLoop_io_read_w4_rsc_cse_sva[5535:5528]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_415_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_43_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_414_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_415_nl));
  assign mul_43_nl = nl_mul_43_nl[28:0];
  assign z_out_77_28_7 = readslicef_29_22_7((mul_43_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_416_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[5039:5032]),
      (MultLoop_io_read_w4_rsc_cse_sva[3207:3200]), (MultLoop_io_read_w4_rsc_cse_sva[5415:5408]),
      (MultLoop_io_read_w4_rsc_cse_sva[6543:6536]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_417_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_44_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_416_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_417_nl));
  assign mul_44_nl = nl_mul_44_nl[28:0];
  assign z_out_78_28_7 = readslicef_29_22_7((mul_44_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_418_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[5031:5024]),
      (MultLoop_io_read_w4_rsc_cse_sva[3215:3208]), (MultLoop_io_read_w4_rsc_cse_sva[4527:4520]),
      (MultLoop_io_read_w4_rsc_cse_sva[5407:5400]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_419_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_45_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_418_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_419_nl));
  assign mul_45_nl = nl_mul_45_nl[28:0];
  assign z_out_79_28_7 = readslicef_29_22_7((mul_45_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_420_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[2599:2592]),
      (w4_rsci_idat_mxwt[2023:2016]), (MultLoop_io_read_w4_rsc_cse_sva[6439:6432]),
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_421_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4])});
  assign nl_mul_46_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_420_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_421_nl));
  assign mul_46_nl = nl_mul_46_nl[28:0];
  assign z_out_80_28_7 = readslicef_29_22_7((mul_46_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_422_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7351:7344]),
      (MultLoop_io_read_w4_rsc_cse_sva[3647:3640]), (w4_rsci_idat_mxwt[2031:2024]),
      (MultLoop_io_read_w4_rsc_cse_sva[7599:7592]), {(fsm_output[4]) , (fsm_output[3])
      , (fsm_output[1]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_423_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_mul_47_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_422_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_423_nl));
  assign mul_47_nl = nl_mul_47_nl[28:0];
  assign z_out_81_28_7 = readslicef_29_22_7((mul_47_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_424_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2199:2192]),
      (w4_rsci_idat_mxwt[4999:4992]), (MultLoop_io_read_w4_rsc_cse_sva[4487:4480]),
      (MultLoop_io_read_w4_rsc_cse_sva[4399:4392]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_425_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_48_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_424_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_425_nl));
  assign mul_48_nl = nl_mul_48_nl[28:0];
  assign z_out_82_28_7 = readslicef_29_22_7((mul_48_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_426_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[6095:6088]),
      (MultLoop_io_read_w4_rsc_cse_sva[1599:1592]), (MultLoop_io_read_w4_rsc_cse_sva[7607:7600]),
      (MultLoop_io_read_w4_rsc_cse_sva[5303:5296]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_427_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_49_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_426_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_427_nl));
  assign mul_49_nl = nl_mul_49_nl[28:0];
  assign z_out_83_28_7 = readslicef_29_22_7((mul_49_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_428_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2191:2184]),
      (w4_rsci_idat_mxwt[5007:5000]), (MultLoop_io_read_w4_rsc_cse_sva[4391:4384]),
      (MultLoop_io_read_w4_rsc_cse_sva[6527:6520]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_429_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_50_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_428_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_429_nl));
  assign mul_50_nl = nl_mul_50_nl[28:0];
  assign z_out_84_28_7 = readslicef_29_22_7((mul_50_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_93_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[6079:6072]),
      (MultLoop_io_read_w4_rsc_cse_sva[5383:5376]), fsm_output[4]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_94_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[4]);
  assign nl_mul_51_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_93_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_94_nl));
  assign mul_51_nl = nl_mul_51_nl[28:0];
  assign z_out_85_28_7 = readslicef_29_22_7((mul_51_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_95_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[9191:9184]),
      (MultLoop_io_read_w4_rsc_cse_sva[5391:5384]), fsm_output[4]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_96_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[4]);
  assign nl_mul_52_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_95_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_96_nl));
  assign mul_52_nl = nl_mul_52_nl[28:0];
  assign z_out_86_28_7 = readslicef_29_22_7((mul_52_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_430_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2183:2176]),
      (w4_rsci_idat_mxwt[5015:5008]), (MultLoop_io_read_w4_rsc_cse_sva[4479:4472]),
      (MultLoop_io_read_w4_rsc_cse_sva[4383:4376]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_431_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_53_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_430_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_431_nl));
  assign mul_53_nl = nl_mul_53_nl[28:0];
  assign z_out_87_28_7 = readslicef_29_22_7((mul_53_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_432_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[6111:6104]),
      (MultLoop_io_read_w4_rsc_cse_sva[4671:4664]), (MultLoop_io_read_w4_rsc_cse_sva[5399:5392]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_433_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_54_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_432_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_433_nl));
  assign mul_54_nl = nl_mul_54_nl[28:0];
  assign z_out_88_28_7 = readslicef_29_22_7((mul_54_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_434_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[5023:5016]),
      (MultLoop_io_read_w4_rsc_cse_sva[3199:3192]), (MultLoop_io_read_w4_rsc_cse_sva[4375:4368]),
      (MultLoop_io_read_w4_rsc_cse_sva[6535:6528]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_435_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_55_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_434_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_435_nl));
  assign mul_55_nl = nl_mul_55_nl[28:0];
  assign z_out_89_28_7 = readslicef_29_22_7((mul_55_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_436_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1423:1416]),
      (w4_rsci_idat_mxwt[5095:5088]), (MultLoop_io_read_w4_rsc_cse_sva[887:880]),
      (MultLoop_io_read_w4_rsc_cse_sva[3327:3320]), (MultLoop_io_read_w4_rsc_cse_sva[5207:5200]),
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_437_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_56_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_436_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_437_nl));
  assign mul_56_nl = nl_mul_56_nl[28:0];
  assign z_out_90_28_7 = readslicef_29_22_7((mul_56_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_438_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1431:1424]),
      (w4_rsci_idat_mxwt[9183:9176]), (MultLoop_io_read_w4_rsc_cse_sva[3271:3264]),
      (MultLoop_io_read_w4_rsc_cse_sva[879:872]), (MultLoop_io_read_w4_rsc_cse_sva[5215:5208]),
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_439_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_57_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_438_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_439_nl));
  assign mul_57_nl = nl_mul_57_nl[28:0];
  assign z_out_91_28_7 = readslicef_29_22_7((mul_57_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_440_nl = MUX1HOT_v_8_7_2((MultLoop_io_read_w4_rsc_cse_sva[8951:8944]),
      (w4_rsci_idat_mxwt[5079:5072]), (MultLoop_io_read_w4_rsc_cse_sva[1375:1368]),
      (MultLoop_io_read_w4_rsc_cse_sva[6335:6328]), (MultLoop_io_read_w4_rsc_cse_sva[1655:1648]),
      (MultLoop_io_read_w4_rsc_cse_sva[2911:2904]), (MultLoop_io_read_w4_rsc_cse_sva[5191:5184]),
      {(fsm_output[7]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_441_nl = MUX1HOT_v_21_7_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[7]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_58_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_440_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_441_nl));
  assign mul_58_nl = nl_mul_58_nl[28:0];
  assign z_out_92_28_7 = readslicef_29_22_7((mul_58_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_442_nl = MUX1HOT_v_8_7_2((MultLoop_io_read_w4_rsc_cse_sva[8551:8544]),
      (MultLoop_io_read_w4_rsc_cse_sva[8943:8936]), (w4_rsci_idat_mxwt[5111:5104]),
      (MultLoop_io_read_w4_rsc_cse_sva[1647:1640]), (MultLoop_io_read_w4_rsc_cse_sva[2919:2912]),
      (MultLoop_io_read_w4_rsc_cse_sva[5199:5192]), (MultLoop_io_read_w4_rsc_cse_sva[5295:5288]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_443_nl = MUX1HOT_v_21_7_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_59_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_442_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_443_nl));
  assign mul_59_nl = nl_mul_59_nl[28:0];
  assign z_out_93_28_7 = readslicef_29_22_7((mul_59_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_444_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1303:1296]),
      (MultLoop_io_read_w4_rsc_cse_sva[8543:8536]), (w4_rsci_idat_mxwt[5103:5096]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_445_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_mul_60_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_444_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_445_nl));
  assign mul_60_nl = nl_mul_60_nl[28:0];
  assign z_out_94_28_7 = readslicef_29_22_7((mul_60_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_446_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1287:1280]),
      (MultLoop_io_read_w4_rsc_cse_sva[8535:8528]), (w4_rsci_idat_mxwt[2983:2976]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_447_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_mul_61_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_446_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_447_nl));
  assign mul_61_nl = nl_mul_61_nl[28:0];
  assign z_out_95_28_7 = readslicef_29_22_7((mul_61_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_448_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[1447:1440]),
      (w4_rsci_idat_mxwt[9199:9192]), (MultLoop_io_read_w4_rsc_cse_sva[2351:2344]),
      (MultLoop_io_read_w4_rsc_cse_sva[871:864]), (MultLoop_io_read_w4_rsc_cse_sva[5223:5216]),
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_449_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_62_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_448_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_449_nl));
  assign mul_62_nl = nl_mul_62_nl[28:0];
  assign z_out_96_28_7 = readslicef_29_22_7((mul_62_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_450_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[3423:3416]),
      (MultLoop_io_read_w4_rsc_cse_sva[863:856]), (MultLoop_io_read_w4_rsc_cse_sva[5231:5224]),
      (MultLoop_io_read_w4_rsc_cse_sva[5375:5368]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_451_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_63_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_450_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_451_nl));
  assign mul_63_nl = nl_mul_63_nl[28:0];
  assign z_out_97_28_7 = readslicef_29_22_7((mul_63_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_452_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2391:2384]),
      (MultLoop_io_read_w4_rsc_cse_sva[2359:2352]), (MultLoop_io_read_w4_rsc_cse_sva[2927:2920]),
      (MultLoop_io_read_w4_rsc_cse_sva[5239:5232]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_453_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_64_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_452_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_453_nl));
  assign mul_64_nl = nl_mul_64_nl[28:0];
  assign z_out_98_28_7 = readslicef_29_22_7((mul_64_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_454_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1439:1432]),
      (MultLoop_io_read_w4_rsc_cse_sva[2231:2224]), (MultLoop_io_read_w4_rsc_cse_sva[2935:2928]),
      (MultLoop_io_read_w4_rsc_cse_sva[4167:4160]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_455_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_65_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_454_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_455_nl));
  assign mul_65_nl = nl_mul_65_nl[28:0];
  assign z_out_99_28_7 = readslicef_29_22_7((mul_65_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_456_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1367:1360]),
      (MultLoop_io_read_w4_rsc_cse_sva[1887:1880]), (MultLoop_io_read_w4_rsc_cse_sva[4175:4168]),
      (MultLoop_io_read_w4_rsc_cse_sva[4351:4344]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_457_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_66_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_456_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_457_nl));
  assign mul_66_nl = nl_mul_66_nl[28:0];
  assign z_out_100_28_7 = readslicef_29_22_7((mul_66_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_458_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2399:2392]),
      (MultLoop_io_read_w4_rsc_cse_sva[2319:2312]), (MultLoop_io_read_w4_rsc_cse_sva[1895:1888]),
      (MultLoop_io_read_w4_rsc_cse_sva[4183:4176]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_459_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_67_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_458_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_459_nl));
  assign mul_67_nl = nl_mul_67_nl[28:0];
  assign z_out_101_28_7 = readslicef_29_22_7((mul_67_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_460_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1407:1400]),
      (MultLoop_io_read_w4_rsc_cse_sva[1295:1288]), (MultLoop_io_read_w4_rsc_cse_sva[2143:2136]),
      (w4_rsci_idat_mxwt[5063:5056]), {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])
      , (fsm_output[1])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_461_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[1])});
  assign nl_mul_68_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_460_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_461_nl));
  assign mul_68_nl = nl_mul_68_nl[28:0];
  assign z_out_102_28_7 = readslicef_29_22_7((mul_68_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_462_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[1415:1408]),
      (MultLoop_io_read_w4_rsc_cse_sva[1319:1312]), (w4_rsci_idat_mxwt[9207:9200]),
      (MultLoop_io_read_w4_rsc_cse_sva[2135:2128]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_463_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_69_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_462_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_463_nl));
  assign mul_69_nl = nl_mul_69_nl[28:0];
  assign z_out_103_28_7 = readslicef_29_22_7((mul_69_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_464_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1311:1304]),
      (MultLoop_io_read_w4_rsc_cse_sva[1383:1376]), (w4_rsci_idat_mxwt[2975:2968]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_465_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_mul_70_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_464_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_465_nl));
  assign mul_70_nl = nl_mul_70_nl[28:0];
  assign z_out_104_28_7 = readslicef_29_22_7((mul_70_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_466_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2151:2144]),
      (MultLoop_io_read_w4_rsc_cse_sva[1215:1208]), (MultLoop_io_read_w4_rsc_cse_sva[1391:1384]),
      (w4_rsci_idat_mxwt[7103:7096]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[1])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_467_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_mul_71_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_466_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_467_nl));
  assign mul_71_nl = nl_mul_71_nl[28:0];
  assign z_out_105_28_7 = readslicef_29_22_7((mul_71_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_468_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2127:2120]),
      (w4_rsci_idat_mxwt[5087:5080]), (MultLoop_io_read_w4_rsc_cse_sva[5311:5304]),
      (MultLoop_io_read_w4_rsc_cse_sva[3439:3432]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_469_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_72_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_468_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_469_nl));
  assign mul_72_nl = nl_mul_72_nl[28:0];
  assign z_out_106_28_7 = readslicef_29_22_7((mul_72_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_470_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2159:2152]),
      (MultLoop_io_read_w4_rsc_cse_sva[8559:8552]), (w4_rsci_idat_mxwt[2991:2984]),
      (MultLoop_io_read_w4_rsc_cse_sva[2343:2336]), {(fsm_output[3]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_471_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[4])});
  assign nl_mul_73_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_470_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_471_nl));
  assign mul_73_nl = nl_mul_73_nl[28:0];
  assign z_out_107_28_7 = readslicef_29_22_7((mul_73_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_472_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1455:1448]),
      (MultLoop_io_read_w4_rsc_cse_sva[1335:1328]), (MultLoop_io_read_w4_rsc_cse_sva[1143:1136]),
      (MultLoop_io_read_w4_rsc_cse_sva[8911:8904]), (w4_rsci_idat_mxwt[2967:2960]),
      (MultLoop_io_read_w4_rsc_cse_sva[3951:3944]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[2])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_473_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_90_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[1])
      , (fsm_output[2])});
  assign nl_mul_74_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_472_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_473_nl));
  assign mul_74_nl = nl_mul_74_nl[28:0];
  assign z_out_108_28_7 = readslicef_29_22_7((mul_74_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_474_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[3431:3424]),
      (MultLoop_io_read_w4_rsc_cse_sva[2335:2328]), (MultLoop_io_read_w4_rsc_cse_sva[1903:1896]),
      (MultLoop_io_read_w4_rsc_cse_sva[4191:4184]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_475_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_12_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_75_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_474_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_475_nl));
  assign mul_75_nl = nl_mul_75_nl[28:0];
  assign z_out_109_28_7 = readslicef_29_22_7((mul_75_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_476_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2407:2400]),
      (MultLoop_io_read_w4_rsc_cse_sva[2327:2320]), (MultLoop_io_read_w4_rsc_cse_sva[1911:1904]),
      (MultLoop_io_read_w4_rsc_cse_sva[4199:4192]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_477_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_13_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_76_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_476_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_477_nl));
  assign mul_76_nl = nl_mul_76_nl[28:0];
  assign z_out_110_28_7 = readslicef_29_22_7((mul_76_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_478_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1327:1320]),
      (MultLoop_io_read_w4_rsc_cse_sva[8935:8928]), (MultLoop_io_read_w4_rsc_cse_sva[2423:2416]),
      (w4_rsci_idat_mxwt[2959:2952]), (MultLoop_io_read_w4_rsc_cse_sva[4983:4976]),
      (MultLoop_io_read_w4_rsc_cse_sva[4207:4200]), {(fsm_output[4]) , (fsm_output[7])
      , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_479_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[4]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3])});
  assign nl_mul_77_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_478_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_479_nl));
  assign mul_77_nl = nl_mul_77_nl[28:0];
  assign z_out_111_28_7 = readslicef_29_22_7((mul_77_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_480_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[8567:8560]),
      (MultLoop_io_read_w4_rsc_cse_sva[8927:8920]), (MultLoop_io_read_w4_rsc_cse_sva[4287:4280]),
      (w4_rsci_idat_mxwt[2951:2944]), (MultLoop_io_read_w4_rsc_cse_sva[3935:3928]),
      (MultLoop_io_read_w4_rsc_cse_sva[4215:4208]), {(fsm_output[5]) , (fsm_output[7])
      , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_481_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_92_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3])});
  assign nl_mul_78_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_480_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_481_nl));
  assign mul_78_nl = nl_mul_78_nl[28:0];
  assign z_out_112_28_7 = readslicef_29_22_7((mul_78_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_482_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[1135:1128]),
      (MultLoop_io_read_w4_rsc_cse_sva[8903:8896]), (MultLoop_io_read_w4_rsc_cse_sva[3415:3408]),
      (w4_rsci_idat_mxwt[2943:2936]), (MultLoop_io_read_w4_rsc_cse_sva[3959:3952]),
      (MultLoop_io_read_w4_rsc_cse_sva[6327:6320]), {(fsm_output[3]) , (fsm_output[7])
      , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_483_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_14_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_89_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_23_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[3]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_mul_79_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_482_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_483_nl));
  assign mul_79_nl = nl_mul_79_nl[28:0];
  assign z_out_113_28_7 = readslicef_29_22_7((mul_79_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_484_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1087:1080]),
      (w4_rsci_idat_mxwt[2007:2000]), (MultLoop_io_read_w4_rsc_cse_sva[9303:9296]),
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_485_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6])});
  assign nl_mul_80_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_484_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_485_nl));
  assign mul_80_nl = nl_mul_80_nl[28:0];
  assign z_out_114_28_7 = readslicef_29_22_7((mul_80_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_486_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[7343:7336]),
      (MultLoop_io_read_w4_rsc_cse_sva[2119:2112]), (MultLoop_io_read_w4_rsc_cse_sva[8919:8912]),
      (MultLoop_io_read_w4_rsc_cse_sva[1399:1392]), (w4_rsci_idat_mxwt[8127:8120]),
      (MultLoop_io_read_w4_rsc_cse_sva[3943:3936]), {(fsm_output[4]) , (fsm_output[3])
      , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_487_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_91_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[2])});
  assign nl_mul_81_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_486_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_487_nl));
  assign mul_81_nl = nl_mul_81_nl[28:0];
  assign z_out_115_28_7 = readslicef_29_22_7((mul_81_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_488_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2167:2160]),
      (w4_rsci_idat_mxwt[1983:1976]), (MultLoop_io_read_w4_rsc_cse_sva[2415:2408]),
      (MultLoop_io_read_w4_rsc_cse_sva[2311:2304]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_489_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_15_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_120_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_82_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_488_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_489_nl));
  assign mul_82_nl = nl_mul_82_nl[28:0];
  assign z_out_116_28_7 = readslicef_29_22_7((mul_82_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_97_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7495:7488]),
      (MultLoop_io_read_w4_rsc_cse_sva[9543:9536]), fsm_output[8]);
  assign nl_mul_83_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_97_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_83_nl = nl_mul_83_nl[28:0];
  assign z_out_117_28_7 = readslicef_29_22_7((mul_83_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_490_nl = MUX1HOT_v_8_7_2((w4_rsci_idat_mxwt[3967:3960]),
      (MultLoop_io_read_w4_rsc_cse_sva[2207:2200]), (MultLoop_io_read_w4_rsc_cse_sva[8895:8888]),
      (MultLoop_io_read_w4_rsc_cse_sva[3591:3584]), (MultLoop_io_read_w4_rsc_cse_sva[4423:4416]),
      (MultLoop_io_read_w4_rsc_cse_sva[8855:8848]), (MultLoop_io_read_w4_rsc_cse_sva[7551:7544]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_491_nl = MUX1HOT_v_21_7_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_88_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[5])});
  assign nl_mul_84_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_490_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_491_nl));
  assign mul_84_nl = nl_mul_84_nl[28:0];
  assign z_out_118_28_7 = readslicef_29_22_7((mul_84_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_492_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[3975:3968]),
      (MultLoop_io_read_w4_rsc_cse_sva[3343:3336]), (MultLoop_io_read_w4_rsc_cse_sva[6503:6496]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_493_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_85_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_492_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_493_nl));
  assign mul_85_nl = nl_mul_85_nl[28:0];
  assign z_out_119_28_7 = readslicef_29_22_7((mul_85_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_494_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[3983:3976]),
      (MultLoop_io_read_w4_rsc_cse_sva[3495:3488]), (MultLoop_io_read_w4_rsc_cse_sva[3351:3344]),
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_495_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_86_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_494_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_495_nl));
  assign mul_86_nl = nl_mul_86_nl[28:0];
  assign z_out_120_28_7 = readslicef_29_22_7((mul_86_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_496_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[5495:5488]),
      (w4_rsci_idat_mxwt[1967:1960]), (MultLoop_io_read_w4_rsc_cse_sva[1823:1816]),
      (MultLoop_io_read_w4_rsc_cse_sva[10239:10232]), (MultLoop_io_read_w4_rsc_cse_sva[1343:1336]),
      (MultLoop_io_read_w4_rsc_cse_sva[1079:1072]), {(fsm_output[5]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_497_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_128_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4])
      , (fsm_output[3])});
  assign nl_mul_87_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_496_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_497_nl));
  assign mul_87_nl = nl_mul_87_nl[28:0];
  assign z_out_121_28_7 = readslicef_29_22_7((mul_87_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_498_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[2215:2208]),
      (MultLoop_io_read_w4_rsc_cse_sva[5463:5456]), (w4_rsci_idat_mxwt[1959:1952]),
      (MultLoop_io_read_w4_rsc_cse_sva[2239:2232]), (MultLoop_io_read_w4_rsc_cse_sva[2567:2560]),
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_499_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2])});
  assign nl_mul_88_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_498_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_499_nl));
  assign mul_88_nl = nl_mul_88_nl[28:0];
  assign z_out_122_28_7 = readslicef_29_22_7((mul_88_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_500_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2367:2360]),
      (w4_rsci_idat_mxwt[8063:8056]), (MultLoop_io_read_w4_rsc_cse_sva[5487:5480]),
      (MultLoop_io_read_w4_rsc_cse_sva[4255:4248]), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_501_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_89_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_500_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_501_nl));
  assign mul_89_nl = nl_mul_89_nl[28:0];
  assign z_out_123_28_7 = readslicef_29_22_7((mul_89_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_502_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[2375:2368]),
      (w4_rsci_idat_mxwt[1975:1968]), (MultLoop_io_read_w4_rsc_cse_sva[5279:5272]),
      (MultLoop_io_read_w4_rsc_cse_sva[5559:5552]), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_503_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_90_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_502_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_503_nl));
  assign mul_90_nl = nl_mul_90_nl[28:0];
  assign z_out_124_28_7 = readslicef_29_22_7((mul_90_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_504_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[1927:1920]),
      (MultLoop_io_read_w4_rsc_cse_sva[5455:5448]), (MultLoop_io_read_w4_rsc_cse_sva[4151:4144]),
      (MultLoop_io_read_w4_rsc_cse_sva[5551:5544]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_505_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_91_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_504_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_505_nl));
  assign mul_91_nl = nl_mul_91_nl[28:0];
  assign z_out_125_28_7 = readslicef_29_22_7((mul_91_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_506_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[8071:8064]),
      (MultLoop_io_read_w4_rsc_cse_sva[3391:3384]), (MultLoop_io_read_w4_rsc_cse_sva[6511:6504]),
      (MultLoop_io_read_w4_rsc_cse_sva[5175:5168]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_507_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_113_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_92_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_506_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_507_nl));
  assign mul_92_nl = nl_mul_92_nl[28:0];
  assign z_out_126_28_7 = readslicef_29_22_7((mul_92_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_98_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[8079:8072]),
      (MultLoop_io_read_w4_rsc_cse_sva[5439:5432]), fsm_output[4]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_99_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[4]);
  assign nl_mul_93_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_98_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_99_nl));
  assign mul_93_nl = nl_mul_93_nl[28:0];
  assign z_out_127_28_7 = readslicef_29_22_7((mul_93_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_100_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8511:8504]),
      (MultLoop_io_read_w4_rsc_cse_sva[9535:9528]), fsm_output[8]);
  assign nl_mul_94_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_100_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_94_nl = nl_mul_94_nl[28:0];
  assign z_out_128_28_7 = readslicef_29_22_7((mul_94_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_508_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[8095:8088]),
      (MultLoop_io_read_w4_rsc_cse_sva[6663:6656]), (MultLoop_io_read_w4_rsc_cse_sva[8879:8872]),
      (MultLoop_io_read_w4_rsc_cse_sva[6487:6480]), (MultLoop_io_read_w4_rsc_cse_sva[5287:5280]),
      (MultLoop_io_read_w4_rsc_cse_sva[1351:1344]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_509_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_43_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[4])});
  assign nl_mul_95_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_508_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_509_nl));
  assign mul_95_nl = nl_mul_95_nl[28:0];
  assign z_out_129_28_7 = readslicef_29_22_7((mul_95_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_510_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[8103:8096]),
      (MultLoop_io_read_w4_rsc_cse_sva[4615:4608]), (MultLoop_io_read_w4_rsc_cse_sva[8887:8880]),
      (MultLoop_io_read_w4_rsc_cse_sva[6519:6512]), (MultLoop_io_read_w4_rsc_cse_sva[1191:1184]),
      (MultLoop_io_read_w4_rsc_cse_sva[2383:2376]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_511_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_117_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[4])});
  assign nl_mul_96_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_510_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_511_nl));
  assign mul_96_nl = nl_mul_96_nl[28:0];
  assign z_out_130_28_7 = readslicef_29_22_7((mul_96_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_512_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[8111:8104]),
      (MultLoop_io_read_w4_rsc_cse_sva[4263:4256]), (MultLoop_io_read_w4_rsc_cse_sva[3503:3496]),
      (MultLoop_io_read_w4_rsc_cse_sva[3367:3360]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_513_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_118_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_97_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_512_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_513_nl));
  assign mul_97_nl = nl_mul_97_nl[28:0];
  assign z_out_131_28_7 = readslicef_29_22_7((mul_97_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_514_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[8119:8112]),
      (MultLoop_io_read_w4_rsc_cse_sva[3511:3504]), (MultLoop_io_read_w4_rsc_cse_sva[3359:3352]),
      (MultLoop_io_read_w4_rsc_cse_sva[6199:6192]), {(fsm_output[1]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_515_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_119_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_98_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_514_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_515_nl));
  assign mul_98_nl = nl_mul_98_nl[28:0];
  assign z_out_132_28_7 = readslicef_29_22_7((mul_98_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_516_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[3231:3224]),
      (MultLoop_io_read_w4_rsc_cse_sva[5471:5464]), (w4_rsci_idat_mxwt[1919:1912]),
      (MultLoop_io_read_w4_rsc_cse_sva[5639:5632]), (MultLoop_io_read_w4_rsc_cse_sva[3383:3376]),
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_517_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
  assign nl_mul_99_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_516_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_517_nl));
  assign mul_99_nl = nl_mul_99_nl[28:0];
  assign z_out_133_28_7 = readslicef_29_22_7((mul_99_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_518_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[3239:3232]),
      (MultLoop_io_read_w4_rsc_cse_sva[1543:1536]), (MultLoop_io_read_w4_rsc_cse_sva[8591:8584]),
      (MultLoop_io_read_w4_rsc_cse_sva[4431:4424]), {(fsm_output[3]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_519_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[3]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_mul_100_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_518_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_519_nl));
  assign mul_100_nl = nl_mul_100_nl[28:0];
  assign z_out_134_28_7 = readslicef_29_22_7((mul_100_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_520_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[1951:1944]),
      (MultLoop_io_read_w4_rsc_cse_sva[7687:7680]), (MultLoop_io_read_w4_rsc_cse_sva[8871:8864]),
      (MultLoop_io_read_w4_rsc_cse_sva[1359:1352]), (MultLoop_io_read_w4_rsc_cse_sva[1183:1176]),
      (MultLoop_io_read_w4_rsc_cse_sva[5543:5536]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_521_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_116_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_85_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[3])
      , (fsm_output[5])});
  assign nl_mul_101_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_520_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_521_nl));
  assign mul_101_nl = nl_mul_101_nl[28:0];
  assign z_out_135_28_7 = readslicef_29_22_7((mul_101_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_522_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[3399:3392]),
      (MultLoop_io_read_w4_rsc_cse_sva[5479:5472]), (w4_rsci_idat_mxwt[1935:1928]),
      (MultLoop_io_read_w4_rsc_cse_sva[10015:10008]), (MultLoop_io_read_w4_rsc_cse_sva[6215:6208]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_523_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_114_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_mul_102_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_522_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_523_nl));
  assign mul_102_nl = nl_mul_102_nl[28:0];
  assign z_out_136_28_7 = readslicef_29_22_7((mul_102_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_524_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[6015:6008]),
      (MultLoop_io_read_w4_rsc_cse_sva[3375:3368]), (MultLoop_io_read_w4_rsc_cse_sva[6495:6488]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_525_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_112_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_44_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_103_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_524_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_525_nl));
  assign mul_103_nl = nl_mul_103_nl[28:0];
  assign z_out_137_28_7 = readslicef_29_22_7((mul_103_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_526_nl = MUX1HOT_v_8_6_2((w4_rsci_idat_mxwt[6087:6080]),
      (MultLoop_io_read_w4_rsc_cse_sva[3127:3120]), (MultLoop_io_read_w4_rsc_cse_sva[9311:9304]),
      (MultLoop_io_read_w4_rsc_cse_sva[2847:2840]), (MultLoop_io_read_w4_rsc_cse_sva[4415:4408]),
      (MultLoop_io_read_w4_rsc_cse_sva[7567:7560]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_527_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_mul_104_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_526_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_527_nl));
  assign mul_104_nl = nl_mul_104_nl[28:0];
  assign z_out_138_28_7 = readslicef_29_22_7((mul_104_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_528_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[7359:7352]),
      (w4_rsci_idat_mxwt[6127:6120]), (MultLoop_io_read_w4_rsc_cse_sva[9327:9320]),
      (MultLoop_io_read_w4_rsc_cse_sva[10007:10000]), (MultLoop_io_read_w4_rsc_cse_sva[2103:2096]),
      (MultLoop_io_read_w4_rsc_cse_sva[7575:7568]), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_529_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_24_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[5])});
  assign nl_mul_105_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_528_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_529_nl));
  assign mul_105_nl = nl_mul_105_nl[28:0];
  assign z_out_139_28_7 = readslicef_29_22_7((mul_105_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_530_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[3407:3400]),
      (MultLoop_io_read_w4_rsc_cse_sva[2839:2832]), (MultLoop_io_read_w4_rsc_cse_sva[8583:8576]),
      (MultLoop_io_read_w4_rsc_cse_sva[5271:5264]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_531_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_106_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_530_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_531_nl));
  assign mul_106_nl = nl_mul_106_nl[28:0];
  assign z_out_140_28_7 = readslicef_29_22_7((mul_106_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_532_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[2111:2104]),
      (w4_rsci_idat_mxwt[1999:1992]), (MultLoop_io_read_w4_rsc_cse_sva[9319:9312]),
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_533_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6])});
  assign nl_mul_107_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_532_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_533_nl));
  assign mul_107_nl = nl_mul_107_nl[28:0];
  assign z_out_141_28_7 = readslicef_29_22_7((mul_107_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_534_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[1943:1936]),
      (MultLoop_io_read_w4_rsc_cse_sva[1815:1808]), (MultLoop_io_read_w4_rsc_cse_sva[6463:6456]),
      (MultLoop_io_read_w4_rsc_cse_sva[7559:7552]), (MultLoop_io_read_w4_rsc_cse_sva[5247:5240]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_535_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_115_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_16_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_mul_108_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_534_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_535_nl));
  assign mul_108_nl = nl_mul_108_nl[28:0];
  assign z_out_142_28_7 = readslicef_29_22_7((mul_108_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_536_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[799:792]),
      (MultLoop_io_read_w4_rsc_cse_sva[8599:8592]), (MultLoop_io_read_w4_rsc_cse_sva[6479:6472]),
      (MultLoop_io_read_w4_rsc_cse_sva[5263:5256]), {(fsm_output[2]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_537_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_100_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_18_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_109_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_536_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_537_nl));
  assign mul_109_nl = nl_mul_109_nl[28:0];
  assign z_out_143_28_7 = readslicef_29_22_7((mul_109_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_538_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[791:784]),
      (MultLoop_io_read_w4_rsc_cse_sva[8575:8568]), (MultLoop_io_read_w4_rsc_cse_sva[6471:6464]),
      (MultLoop_io_read_w4_rsc_cse_sva[5255:5248]), {(fsm_output[2]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_539_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_99_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_17_if_exu_pmx_20_0_lpi_1_dfm_mx0w1,
      {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_110_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_538_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_539_nl));
  assign mul_110_nl = nl_mul_110_nl[28:0];
  assign z_out_144_28_7 = readslicef_29_22_7((mul_110_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_101_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[2039:2032]),
      (MultLoop_io_read_w4_rsc_cse_sva[3623:3616]), fsm_output[3]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_102_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[3]);
  assign nl_mul_111_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_101_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_102_nl));
  assign mul_111_nl = nl_mul_111_nl[28:0];
  assign z_out_145_28_7 = readslicef_29_22_7((mul_111_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_103_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[10151:10144]),
      (MultLoop_io_read_w4_rsc_cse_sva[847:840]), fsm_output[8]);
  assign nl_mul_112_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_103_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_112_nl = nl_mul_112_nl[28:0];
  assign z_out_146_28_7 = readslicef_29_22_7((mul_112_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_104_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[10143:10136]),
      (MultLoop_io_read_w4_rsc_cse_sva[839:832]), fsm_output[8]);
  assign nl_mul_113_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_104_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_113_nl = nl_mul_113_nl[28:0];
  assign z_out_147_28_7 = readslicef_29_22_7((mul_113_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_105_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[10135:10128]),
      (MultLoop_io_read_w4_rsc_cse_sva[831:824]), fsm_output[8]);
  assign nl_mul_114_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_105_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_114_nl = nl_mul_114_nl[28:0];
  assign z_out_148_28_7 = readslicef_29_22_7((mul_114_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse = (fsm_output[5])
      | (fsm_output[8]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_540_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[7463:7456]),
      (MultLoop_io_read_w4_rsc_cse_sva[9367:9360]), (MultLoop_io_read_w4_rsc_cse_sva[10199:10192]),
      (MultLoop_io_read_w4_rsc_cse_sva[7271:7264]), (MultLoop_io_read_w4_rsc_cse_sva[295:288]),
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_541_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm,
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse , (fsm_output[6])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse});
  assign nl_mul_115_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_540_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_541_nl));
  assign mul_115_nl = nl_mul_115_nl[28:0];
  assign z_out_149_28_7 = readslicef_29_22_7((mul_115_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_542_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[7471:7464]),
      (MultLoop_io_read_w4_rsc_cse_sva[9375:9368]), (MultLoop_io_read_w4_rsc_cse_sva[10207:10200]),
      (MultLoop_io_read_w4_rsc_cse_sva[7279:7272]), (MultLoop_io_read_w4_rsc_cse_sva[9519:9512]),
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_543_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm,
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse , (fsm_output[6])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse});
  assign nl_mul_116_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_542_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_543_nl));
  assign mul_116_nl = nl_mul_116_nl[28:0];
  assign z_out_150_28_7 = readslicef_29_22_7((mul_116_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_544_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[7295:7288]),
      (MultLoop_io_read_w4_rsc_cse_sva[9343:9336]), (MultLoop_io_read_w4_rsc_cse_sva[8319:8312]),
      (MultLoop_io_read_w4_rsc_cse_sva[10223:10216]), (MultLoop_io_read_w4_rsc_cse_sva[783:776]),
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_106_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[8]);
  assign nl_mul_117_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_544_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_106_nl));
  assign mul_117_nl = nl_mul_117_nl[28:0];
  assign z_out_151_28_7 = readslicef_29_22_7((mul_117_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_545_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[7303:7296]),
      (MultLoop_io_read_w4_rsc_cse_sva[9351:9344]), (MultLoop_io_read_w4_rsc_cse_sva[8327:8320]),
      (MultLoop_io_read_w4_rsc_cse_sva[10231:10224]), (MultLoop_io_read_w4_rsc_cse_sva[775:768]),
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_107_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[8]);
  assign nl_mul_118_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_545_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_107_nl));
  assign mul_118_nl = nl_mul_118_nl[28:0];
  assign z_out_152_28_7 = readslicef_29_22_7((mul_118_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_108_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[10127:10120]),
      (MultLoop_io_read_w4_rsc_cse_sva[823:816]), fsm_output[8]);
  assign nl_mul_119_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_108_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_119_nl = nl_mul_119_nl[28:0];
  assign z_out_153_28_7 = readslicef_29_22_7((mul_119_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_109_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8527:8520]),
      (MultLoop_io_read_w4_rsc_cse_sva[9551:9544]), fsm_output[8]);
  assign nl_mul_120_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_109_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_120_nl = nl_mul_120_nl[28:0];
  assign z_out_154_28_7 = readslicef_29_22_7((mul_120_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_110_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[2607:2600]),
      (w4_rsci_idat_mxwt[2015:2008]), fsm_output[1]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_111_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[1]);
  assign nl_mul_121_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_110_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_111_nl));
  assign mul_121_nl = nl_mul_121_nl[28:0];
  assign z_out_155_28_7 = readslicef_29_22_7((mul_121_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_546_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[8303:8296]),
      (MultLoop_io_read_w4_rsc_cse_sva[6255:6248]), (MultLoop_io_read_w4_rsc_cse_sva[111:104]),
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_122_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_546_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_122_nl = nl_mul_122_nl[28:0];
  assign z_out_156_28_7 = readslicef_29_22_7((mul_122_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_112_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[6279:6272]),
      (MultLoop_io_read_w4_rsc_cse_sva[135:128]), fsm_output[8]);
  assign nl_mul_123_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_112_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_123_nl = nl_mul_123_nl[28:0];
  assign z_out_157_28_7 = readslicef_29_22_7((mul_123_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_42_cse = (fsm_output[5])
      | (fsm_output[4]) | (fsm_output[8]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_547_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9383:9376]),
      (MultLoop_io_read_w4_rsc_cse_sva[8287:8280]), (MultLoop_io_read_w4_rsc_cse_sva[6239:6232]),
      (MultLoop_io_read_w4_rsc_cse_sva[95:88]), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_113_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_42_cse);
  assign nl_mul_124_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_547_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_113_nl));
  assign mul_124_nl = nl_mul_124_nl[28:0];
  assign z_out_158_28_7 = readslicef_29_22_7((mul_124_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_548_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9439:9432]),
      (MultLoop_io_read_w4_rsc_cse_sva[8295:8288]), (MultLoop_io_read_w4_rsc_cse_sva[6247:6240]),
      (MultLoop_io_read_w4_rsc_cse_sva[103:96]), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_114_nl = MUX_v_21_2_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_42_cse);
  assign nl_mul_125_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_548_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_114_nl));
  assign mul_125_nl = nl_mul_125_nl[28:0];
  assign z_out_159_28_7 = readslicef_29_22_7((mul_125_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_549_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[9447:9440]),
      (MultLoop_io_read_w4_rsc_cse_sva[8423:8416]), (MultLoop_io_read_w4_rsc_cse_sva[10167:10160]),
      (MultLoop_io_read_w4_rsc_cse_sva[6223:6216]), (MultLoop_io_read_w4_rsc_cse_sva[231:224]),
      {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_115_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm,
      operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse);
  assign nl_mul_126_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_549_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_115_nl));
  assign mul_126_nl = nl_mul_126_nl[28:0];
  assign z_out_160_28_7 = readslicef_29_22_7((mul_126_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_550_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[9455:9448]),
      (MultLoop_io_read_w4_rsc_cse_sva[8431:8424]), (MultLoop_io_read_w4_rsc_cse_sva[10175:10168]),
      (MultLoop_io_read_w4_rsc_cse_sva[6231:6224]), (MultLoop_io_read_w4_rsc_cse_sva[239:232]),
      {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_116_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm,
      operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse);
  assign nl_mul_127_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_550_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_116_nl));
  assign mul_127_nl = nl_mul_127_nl[28:0];
  assign z_out_161_28_7 = readslicef_29_22_7((mul_127_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_551_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[9463:9456]),
      (MultLoop_io_read_w4_rsc_cse_sva[8439:8432]), (MultLoop_io_read_w4_rsc_cse_sva[10191:10184]),
      (MultLoop_io_read_w4_rsc_cse_sva[7263:7256]), (MultLoop_io_read_w4_rsc_cse_sva[247:240]),
      {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_117_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm,
      operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse);
  assign nl_mul_128_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_551_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_117_nl));
  assign mul_128_nl = nl_mul_128_nl[28:0];
  assign z_out_162_28_7 = readslicef_29_22_7((mul_128_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_118_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8455:8448]),
      (MultLoop_io_read_w4_rsc_cse_sva[263:256]), fsm_output[8]);
  assign nl_mul_129_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_118_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_129_nl = nl_mul_129_nl[28:0];
  assign z_out_163_28_7 = readslicef_29_22_7((mul_129_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_119_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8487:8480]),
      (MultLoop_io_read_w4_rsc_cse_sva[9511:9504]), fsm_output[8]);
  assign nl_mul_130_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_119_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_37_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_130_nl = nl_mul_130_nl[28:0];
  assign z_out_164_28_7 = readslicef_29_22_7((mul_130_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_120_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8495:8488]),
      (MultLoop_io_read_w4_rsc_cse_sva[303:296]), fsm_output[8]);
  assign nl_mul_131_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_120_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_38_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_131_nl = nl_mul_131_nl[28:0];
  assign z_out_165_28_7 = readslicef_29_22_7((mul_131_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_552_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8271:8264]),
      (MultLoop_io_read_w4_rsc_cse_sva[9143:9136]), (MultLoop_io_read_w4_rsc_cse_sva[7247:7240]),
      (MultLoop_io_read_w4_rsc_cse_sva[79:72]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_132_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_552_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_132_nl = nl_mul_132_nl[28:0];
  assign z_out_166_28_7 = readslicef_29_22_7((mul_132_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_553_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8279:8272]),
      (MultLoop_io_read_w4_rsc_cse_sva[9151:9144]), (MultLoop_io_read_w4_rsc_cse_sva[7255:7248]),
      (MultLoop_io_read_w4_rsc_cse_sva[87:80]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_133_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_553_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_133_nl = nl_mul_133_nl[28:0];
  assign z_out_167_28_7 = readslicef_29_22_7((mul_133_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_121_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[6271:6264]),
      (MultLoop_io_read_w4_rsc_cse_sva[127:120]), fsm_output[8]);
  assign nl_mul_134_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_121_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_134_nl = nl_mul_134_nl[28:0];
  assign z_out_168_28_7 = readslicef_29_22_7((mul_134_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_554_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[7423:7416]),
      (MultLoop_io_read_w4_rsc_cse_sva[2095:2088]), (MultLoop_io_read_w4_rsc_cse_sva[9471:9464]),
      (w4_rsci_idat_mxwt[6103:6096]), (MultLoop_io_read_w4_rsc_cse_sva[9295:9288]),
      (MultLoop_io_read_w4_rsc_cse_sva[3135:3128]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_555_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[3])});
  assign nl_mul_135_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_554_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_555_nl));
  assign mul_135_nl = nl_mul_135_nl[28:0];
  assign z_out_169_28_7 = readslicef_29_22_7((mul_135_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_556_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[6743:6736]),
      (MultLoop_io_read_w4_rsc_cse_sva[7767:7760]), (MultLoop_io_read_w4_rsc_cse_sva[599:592]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_136_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_556_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_136_nl = nl_mul_136_nl[28:0];
  assign z_out_170_28_7 = readslicef_29_22_7((mul_136_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse = (fsm_output[4])
      | (fsm_output[8]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_557_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7439:7432]),
      (MultLoop_io_read_w4_rsc_cse_sva[9487:9480]), (MultLoop_io_read_w4_rsc_cse_sva[6719:6712]),
      (MultLoop_io_read_w4_rsc_cse_sva[575:568]), {(fsm_output[5]) , (fsm_output[7])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_122_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse);
  assign nl_mul_137_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_557_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_122_nl));
  assign mul_137_nl = nl_mul_137_nl[28:0];
  assign z_out_171_28_7 = readslicef_29_22_7((mul_137_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_558_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[6735:6728]),
      (MultLoop_io_read_w4_rsc_cse_sva[7759:7752]), (MultLoop_io_read_w4_rsc_cse_sva[591:584]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_138_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_558_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_138_nl = nl_mul_138_nl[28:0];
  assign z_out_172_28_7 = readslicef_29_22_7((mul_138_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_559_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[6727:6720]),
      (MultLoop_io_read_w4_rsc_cse_sva[7751:7744]), (MultLoop_io_read_w4_rsc_cse_sva[583:576]),
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_139_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_559_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_139_nl = nl_mul_139_nl[28:0];
  assign z_out_173_28_7 = readslicef_29_22_7((mul_139_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_560_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8263:8256]),
      (MultLoop_io_read_w4_rsc_cse_sva[9287:9280]), (MultLoop_io_read_w4_rsc_cse_sva[6703:6696]),
      (MultLoop_io_read_w4_rsc_cse_sva[559:552]), {(fsm_output[5]) , (fsm_output[6])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_123_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse);
  assign nl_mul_140_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_560_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_123_nl));
  assign mul_140_nl = nl_mul_140_nl[28:0];
  assign z_out_174_28_7 = readslicef_29_22_7((mul_140_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_561_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[7735:7728]),
      (MultLoop_io_read_w4_rsc_cse_sva[6711:6704]), (MultLoop_io_read_w4_rsc_cse_sva[567:560]),
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_141_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_561_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_141_nl = nl_mul_141_nl[28:0];
  assign z_out_175_28_7 = readslicef_29_22_7((mul_141_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_562_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7479:7472]),
      (MultLoop_io_read_w4_rsc_cse_sva[9479:9472]), (MultLoop_io_read_w4_rsc_cse_sva[10159:10152]),
      (MultLoop_io_read_w4_rsc_cse_sva[311:304]), {(fsm_output[5]) , (fsm_output[7])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_563_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm,
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse , (fsm_output[7])
      , (fsm_output[2])});
  assign nl_mul_142_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_562_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_563_nl));
  assign mul_142_nl = nl_mul_142_nl[28:0];
  assign z_out_176_28_7 = readslicef_29_22_7((mul_142_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_564_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9223:9216]),
      (w4_rsci_idat_mxwt[1991:1984]), (MultLoop_io_read_w4_rsc_cse_sva[5183:5176]),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_565_nl = MUX1HOT_v_21_3_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_143_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_564_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_565_nl));
  assign mul_143_nl = nl_mul_143_nl[28:0];
  assign z_out_177_28_7 = readslicef_29_22_7((mul_143_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_566_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8255:8248]),
      (MultLoop_io_read_w4_rsc_cse_sva[9279:9272]), (MultLoop_io_read_w4_rsc_cse_sva[6695:6688]),
      (MultLoop_io_read_w4_rsc_cse_sva[551:544]), {(fsm_output[5]) , (fsm_output[6])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_124_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse);
  assign nl_mul_144_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_566_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_124_nl));
  assign mul_144_nl = nl_mul_144_nl[28:0];
  assign z_out_178_28_7 = readslicef_29_22_7((mul_144_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_125_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8503:8496]),
      (MultLoop_io_read_w4_rsc_cse_sva[9527:9520]), fsm_output[8]);
  assign nl_mul_145_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_125_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_39_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_145_nl = nl_mul_145_nl[28:0];
  assign z_out_179_28_7 = readslicef_29_22_7((mul_145_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_567_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[7711:7704]),
      (MultLoop_io_read_w4_rsc_cse_sva[6687:6680]), (MultLoop_io_read_w4_rsc_cse_sva[543:536]),
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_146_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_567_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_146_nl = nl_mul_146_nl[28:0];
  assign z_out_180_28_7 = readslicef_29_22_7((mul_146_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_126_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7503:7496]),
      (MultLoop_io_read_w4_rsc_cse_sva[335:328]), fsm_output[8]);
  assign nl_mul_147_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_126_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_42_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_147_nl = nl_mul_147_nl[28:0];
  assign z_out_181_28_7 = readslicef_29_22_7((mul_147_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_127_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8519:8512]),
      (MultLoop_io_read_w4_rsc_cse_sva[327:320]), fsm_output[8]);
  assign nl_mul_148_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_127_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_41_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_148_nl = nl_mul_148_nl[28:0];
  assign z_out_182_28_7 = readslicef_29_22_7((mul_148_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_128_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7487:7480]),
      (MultLoop_io_read_w4_rsc_cse_sva[319:312]), fsm_output[8]);
  assign nl_mul_149_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_128_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_40_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_149_nl = nl_mul_149_nl[28:0];
  assign z_out_183_28_7 = readslicef_29_22_7((mul_149_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_129_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[6119:6112]),
      (MultLoop_io_read_w4_rsc_cse_sva[3631:3624]), fsm_output[3]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_130_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[3]);
  assign nl_mul_150_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_129_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_130_nl));
  assign mul_150_nl = nl_mul_150_nl[28:0];
  assign z_out_184_28_7 = readslicef_29_22_7((mul_150_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_568_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[8479:8472]),
      (MultLoop_io_read_w4_rsc_cse_sva[9503:9496]), (MultLoop_io_read_w4_rsc_cse_sva[287:280]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_mul_151_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_568_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_151_nl = nl_mul_151_nl[28:0];
  assign z_out_185_28_7 = readslicef_29_22_7((mul_151_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_569_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9495:9488]),
      (MultLoop_io_read_w4_rsc_cse_sva[8471:8464]), (MultLoop_io_read_w4_rsc_cse_sva[279:272]),
      {(fsm_output[7]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_152_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_569_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_152_nl = nl_mul_152_nl[28:0];
  assign z_out_186_28_7 = readslicef_29_22_7((mul_152_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_131_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8463:8456]),
      (MultLoop_io_read_w4_rsc_cse_sva[271:264]), fsm_output[8]);
  assign nl_mul_153_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_131_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_34_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_153_nl = nl_mul_153_nl[28:0];
  assign z_out_187_28_7 = readslicef_29_22_7((mul_153_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_132_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[8447:8440]),
      (MultLoop_io_read_w4_rsc_cse_sva[255:248]), fsm_output[8]);
  assign nl_mul_154_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_132_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_32_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_154_nl = nl_mul_154_nl[28:0];
  assign z_out_188_28_7 = readslicef_29_22_7((mul_154_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_570_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9271:9264]),
      (MultLoop_io_read_w4_rsc_cse_sva[7223:7216]), (MultLoop_io_read_w4_rsc_cse_sva[55:48]),
      {(fsm_output[6]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_155_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_570_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_155_nl = nl_mul_155_nl[28:0];
  assign z_out_189_28_7 = readslicef_29_22_7((mul_155_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_133_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[9263:9256]),
      (MultLoop_io_read_w4_rsc_cse_sva[47:40]), fsm_output[8]);
  assign nl_mul_156_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_133_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_156_nl = nl_mul_156_nl[28:0];
  assign z_out_190_28_7 = readslicef_29_22_7((mul_156_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_571_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9255:9248]),
      (MultLoop_io_read_w4_rsc_cse_sva[7207:7200]), (MultLoop_io_read_w4_rsc_cse_sva[39:32]),
      {(fsm_output[6]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_157_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_571_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_157_nl = nl_mul_157_nl[28:0];
  assign z_out_191_28_7 = readslicef_29_22_7((mul_157_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_572_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9247:9240]),
      (MultLoop_io_read_w4_rsc_cse_sva[7199:7192]), (MultLoop_io_read_w4_rsc_cse_sva[31:24]),
      {(fsm_output[6]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_mul_158_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_572_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_158_nl = nl_mul_158_nl[28:0];
  assign z_out_192_28_7 = readslicef_29_22_7((mul_158_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_573_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8311:8304]),
      (MultLoop_io_read_w4_rsc_cse_sva[9335:9328]), (MultLoop_io_read_w4_rsc_cse_sva[10215:10208]),
      (MultLoop_io_read_w4_rsc_cse_sva[9815:9808]), {(fsm_output[5]) , (fsm_output[6])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_134_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[8]);
  assign nl_mul_159_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_573_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_134_nl));
  assign mul_159_nl = nl_mul_159_nl[28:0];
  assign z_out_193_28_7 = readslicef_29_22_7((mul_159_nl));
  assign MultLoop_mux1h_310_nl = MUX1HOT_v_22_4_2(z_out_42_28_7, z_out_105_28_7,
      z_out_44_28_7, z_out_643_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[3])});
  assign MultLoop_mux1h_311_nl = MUX1HOT_v_22_4_2(z_out_44_28_7, z_out_115_28_7,
      z_out_43_28_7, z_out_644_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[3])});
  assign nl_z_out_194 = (MultLoop_mux1h_310_nl) + (MultLoop_mux1h_311_nl);
  assign z_out_194 = nl_z_out_194[21:0];
  assign MultLoop_mux1h_312_nl = MUX1HOT_v_22_3_2(z_out_155_28_7, z_out_57_28_7,
      z_out_810, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1290_nl = z_out_466 + MultLoop_acc_504_itm;
  assign MultLoop_acc_1290_nl = nl_MultLoop_acc_1290_nl[21:0];
  assign MultLoop_mux1h_313_nl = MUX1HOT_v_22_3_2(z_out_80_28_7, z_out_52_28_7, (MultLoop_acc_1290_nl),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_195 = (MultLoop_mux1h_312_nl) + (MultLoop_mux1h_313_nl);
  assign z_out_195 = nl_z_out_195[21:0];
  assign MultLoop_mux1h_314_nl = MUX1HOT_v_22_4_2(z_out_102_28_7, z_out_60_28_7,
      z_out_663_28_7, z_out_54_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3])});
  assign MultLoop_mux1h_315_nl = MUX1HOT_v_22_4_2(z_out_103_28_7, z_out_56_28_7,
      z_out_662_28_7, z_out_42_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3])});
  assign nl_z_out_196 = (MultLoop_mux1h_314_nl) + (MultLoop_mux1h_315_nl);
  assign z_out_196 = nl_z_out_196[21:0];
  assign MultLoop_mux1h_316_nl = MUX1HOT_v_22_5_2(z_out_107_28_7, z_out_85_28_7,
      z_out_37_28_7, z_out_42_28_7, z_out_181_28_7, {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])});
  assign MultLoop_mux1h_317_nl = MUX1HOT_v_22_5_2(z_out_116_28_7, z_out_138_28_7,
      z_out_59_28_7, z_out_36_28_7, z_out_52_28_7, {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_z_out_197 = (MultLoop_mux1h_316_nl) + (MultLoop_mux1h_317_nl);
  assign z_out_197 = nl_z_out_197[21:0];
  assign MultLoop_mux1h_318_nl = MUX1HOT_v_22_4_2(z_out_92_28_7, z_out_656_28_7,
      z_out_111_28_7, z_out_47_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3])});
  assign MultLoop_mux1h_319_nl = MUX1HOT_v_22_4_2(z_out_104_28_7, z_out_655_28_7,
      z_out_108_28_7, z_out_48_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3])});
  assign nl_z_out_198 = (MultLoop_mux1h_318_nl) + (MultLoop_mux1h_319_nl);
  assign z_out_198 = nl_z_out_198[21:0];
  assign MultLoop_mux1h_320_nl = MUX1HOT_v_22_6_2(z_out_90_28_7, z_out_643_28_7,
      z_out_638_28_7, z_out_98_28_7, z_out_46_28_7, z_out_68_28_7, {(fsm_output[5])
      , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])});
  assign MultLoop_mux1h_321_nl = MUX1HOT_v_22_6_2(z_out_91_28_7, z_out_36_28_7, z_out_631_28_7,
      z_out_99_28_7, z_out_37_28_7, z_out_34_28_7, {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])});
  assign nl_z_out_199 = (MultLoop_mux1h_320_nl) + (MultLoop_mux1h_321_nl);
  assign z_out_199 = nl_z_out_199[21:0];
  assign MultLoop_mux1h_322_nl = MUX1HOT_v_22_7_2(z_out_99_28_7, z_out_116_28_7,
      z_out_658_28_7, z_out_631_28_7, z_out_109_28_7, z_out_42_28_7, z_out_645_28_7,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[3])});
  assign MultLoop_mux1h_323_nl = MUX1HOT_v_22_7_2(z_out_96_28_7, z_out_177_28_7,
      z_out_657_28_7, z_out_633_28_7, z_out_110_28_7, z_out_43_28_7, z_out_646_28_7,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[3])});
  assign nl_z_out_200 = (MultLoop_mux1h_322_nl) + (MultLoop_mux1h_323_nl);
  assign z_out_200 = nl_z_out_200[21:0];
  assign MultLoop_mux1h_324_nl = MUX1HOT_v_22_6_2(z_out_108_28_7, z_out_141_28_7,
      z_out_662_28_7, z_out_93_28_7, z_out_100_28_7, z_out_169_28_7, {(fsm_output[5])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[2]) , (fsm_output[3])});
  assign MultLoop_mux1h_325_nl = MUX1HOT_v_22_6_2(z_out_36_28_7, z_out_114_28_7,
      z_out_637_28_7, z_out_92_28_7, z_out_101_28_7, z_out_45_28_7, {(fsm_output[5])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_z_out_201 = (MultLoop_mux1h_324_nl) + (MultLoop_mux1h_325_nl);
  assign z_out_201 = nl_z_out_201[21:0];
  assign MultLoop_mux1h_326_nl = MUX1HOT_v_22_5_2(z_out_659_28_7, z_out_116_28_7,
      z_out_115_28_7, z_out_92_28_7, z_out_651_28_7, {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign MultLoop_mux1h_327_nl = MUX1HOT_v_22_5_2(z_out_645_28_7, z_out_111_28_7,
      z_out_648_28_7, z_out_93_28_7, z_out_652_28_7, {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_z_out_202 = (MultLoop_mux1h_326_nl) + (MultLoop_mux1h_327_nl);
  assign z_out_202 = nl_z_out_202[21:0];
  assign MultLoop_mux1h_328_nl = MUX1HOT_v_22_4_2(z_out_102_28_7, z_out_646_28_7,
      z_out_104_28_7, z_out_38_28_7, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5])});
  assign MultLoop_mux1h_329_nl = MUX1HOT_v_22_4_2(z_out_105_28_7, z_out_651_28_7,
      z_out_95_28_7, z_out_37_28_7, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5])});
  assign nl_z_out_203 = (MultLoop_mux1h_328_nl) + (MultLoop_mux1h_329_nl);
  assign z_out_203 = nl_z_out_203[21:0];
  assign MultLoop_mux1h_330_nl = MUX1HOT_v_22_3_2(z_out_657_28_7, z_out_642_28_7,
      z_out_811, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_331_nl = MUX1HOT_v_22_3_2(z_out_642_28_7, z_out_53_28_7,
      z_out_821, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_204 = (MultLoop_mux1h_330_nl) + (MultLoop_mux1h_331_nl);
  assign z_out_204 = nl_z_out_204[21:0];
  assign MultLoop_mux1h_332_nl = MUX1HOT_v_22_3_2(z_out_51_28_7, z_out_655_28_7,
      z_out_41_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0))
      * $signed((w4_rsci_idat_mxwt[8151:8144]));
  assign MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign MultLoop_mux1h_333_nl = MUX1HOT_v_22_3_2(z_out_41_28_7, (readslicef_29_22_7((MultLoop_1019_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      z_out_35_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_205 = (MultLoop_mux1h_332_nl) + (MultLoop_mux1h_333_nl);
  assign z_out_205 = nl_z_out_205[21:0];
  assign nl_MultLoop_acc_1291_nl = MultLoop_100_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_667_28_7;
  assign MultLoop_acc_1291_nl = nl_MultLoop_acc_1291_nl[21:0];
  assign AccumDotWidth_mux_82_nl = MUX_v_22_2_2(z_out_821, (MultLoop_acc_1291_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1292_nl = z_out_668_28_7 + z_out_153_28_7;
  assign MultLoop_acc_1292_nl = nl_MultLoop_acc_1292_nl[21:0];
  assign AccumDotWidth_mux_83_nl = MUX_v_22_2_2(z_out_758, (MultLoop_acc_1292_nl),
      fsm_output[8]);
  assign nl_z_out_206 = (AccumDotWidth_mux_82_nl) + (AccumDotWidth_mux_83_nl);
  assign z_out_206 = nl_z_out_206[21:0];
  assign MultLoop_mux1h_334_nl = MUX1HOT_v_22_3_2(z_out_101_28_7, z_out_34_28_7,
      z_out_107_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])});
  assign MultLoop_mux1h_335_nl = MUX1HOT_v_22_3_2(z_out_110_28_7, z_out_58_28_7,
      z_out_60_28_7, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])});
  assign nl_z_out_207 = (MultLoop_mux1h_334_nl) + (MultLoop_mux1h_335_nl);
  assign z_out_207 = nl_z_out_207[21:0];
  assign MultLoop_mux1h_336_nl = MUX1HOT_v_22_4_2(z_out_652_28_7, z_out_113_28_7,
      z_out_51_28_7, z_out_659_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])
      , (fsm_output[3])});
  assign MultLoop_mux1h_337_nl = MUX1HOT_v_22_4_2(z_out_647_28_7, z_out_112_28_7,
      z_out_50_28_7, z_out_662_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])
      , (fsm_output[3])});
  assign nl_z_out_208 = (MultLoop_mux1h_336_nl) + (MultLoop_mux1h_337_nl);
  assign z_out_208 = nl_z_out_208[21:0];
  assign nl_MultLoop_acc_1304_nl = (z_out_1150_29_7[21:0]) + (z_out_934_29_7[21:0]);
  assign MultLoop_acc_1304_nl = nl_MultLoop_acc_1304_nl[21:0];
  assign nl_MultLoop_acc_1305_nl = (z_out_1040_29_7[21:0]) + (z_out_1041_29_7[21:0]);
  assign MultLoop_acc_1305_nl = nl_MultLoop_acc_1305_nl[21:0];
  assign nl_MultLoop_acc_1297_nl = (z_out_1152_29_7[21:0]) + (z_out_1154_29_7[21:0]);
  assign MultLoop_acc_1297_nl = nl_MultLoop_acc_1297_nl[21:0];
  assign nl_MultLoop_acc_1298_nl = (z_out_1153_29_7[21:0]) + (z_out_1151_29_7[21:0]);
  assign MultLoop_acc_1298_nl = nl_MultLoop_acc_1298_nl[21:0];
  assign nl_MultLoop_acc_1300_nl = (z_out_1145_29_7[21:0]) + (z_out_1147_29_7[21:0]);
  assign MultLoop_acc_1300_nl = nl_MultLoop_acc_1300_nl[21:0];
  assign nl_MultLoop_acc_1301_nl = (z_out_1148_29_7[21:0]) + (z_out_1149_29_7[21:0]);
  assign MultLoop_acc_1301_nl = nl_MultLoop_acc_1301_nl[21:0];
  assign nl_MultLoop_acc_1307_nl = (z_out_1043_29_7[21:0]) + (z_out_1036_29_7[21:0]);
  assign MultLoop_acc_1307_nl = nl_MultLoop_acc_1307_nl[21:0];
  assign nl_MultLoop_acc_1308_nl = (z_out_1044_29_7[21:0]) + (z_out_1039_29_7[21:0]);
  assign MultLoop_acc_1308_nl = nl_MultLoop_acc_1308_nl[21:0];
  assign nl_MultLoop_acc_1294_nl = (MultLoop_acc_1304_nl) + (MultLoop_acc_1305_nl)
      + (MultLoop_acc_1297_nl) + (MultLoop_acc_1298_nl) + (MultLoop_acc_1300_nl)
      + (MultLoop_acc_1301_nl) + (MultLoop_acc_1307_nl) + (MultLoop_acc_1308_nl);
  assign MultLoop_acc_1294_nl = nl_MultLoop_acc_1294_nl[21:0];
  assign nl_MultLoop_acc_1293_nl = z_out_475 + (MultLoop_acc_1294_nl);
  assign MultLoop_acc_1293_nl = nl_MultLoop_acc_1293_nl[21:0];
  assign MultLoop_mux1h_338_nl = MUX1HOT_v_22_5_2(z_out_104_28_7, z_out_636_28_7,
      z_out_97_28_7, z_out_100_28_7, (MultLoop_acc_1293_nl), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[8])});
  assign MultLoop_mux1h_339_nl = MUX1HOT_v_22_5_2(z_out_103_28_7, z_out_659_28_7,
      z_out_109_28_7, z_out_101_28_7, z_out_760, {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_209 = (MultLoop_mux1h_338_nl) + (MultLoop_mux1h_339_nl);
  assign z_out_209 = nl_z_out_209[21:0];
  assign MultLoop_mux1h_340_nl = MUX1HOT_v_22_3_2(z_out_81_28_7, z_out_45_28_7, z_out_42_28_7,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_341_nl = MUX1HOT_v_22_3_2(z_out_145_28_7, z_out_43_28_7,
      z_out_34_28_7, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_210 = (MultLoop_mux1h_340_nl) + (MultLoop_mux1h_341_nl);
  assign z_out_210 = nl_z_out_210[21:0];
  assign MultLoop_mux1h_342_nl = MUX1HOT_v_22_3_2(z_out_652_28_7, z_out_649_28_7,
      z_out_819, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_343_nl = MUX1HOT_v_22_3_2(z_out_640_28_7, z_out_50_28_7,
      z_out_846, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_211 = (MultLoop_mux1h_342_nl) + (MultLoop_mux1h_343_nl);
  assign z_out_211 = nl_z_out_211[21:0];
  assign MultLoop_mux1h_344_nl = MUX1HOT_v_22_5_2(z_out_268, z_out_272, MultLoop_acc_215_itm,
      z_out_441, z_out_479, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[3])});
  assign MultLoop_mux1h_345_nl = MUX1HOT_v_22_5_2(z_out_205, z_out_305, MultLoop_acc_105_itm,
      z_out_438, z_out_506, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nl_z_out_212 = (MultLoop_mux1h_344_nl) + (MultLoop_mux1h_345_nl);
  assign z_out_212 = nl_z_out_212[21:0];
  assign MultLoop_mux1h_346_nl = MUX1HOT_v_22_7_2(z_out_196, z_out_268, z_out_506,
      z_out_199, z_out_287, z_out_477, z_out_485, {(fsm_output[5]) , (fsm_output[7])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1312_nl = z_out_243 + MultLoop_acc_724_itm;
  assign MultLoop_acc_1312_nl = nl_MultLoop_acc_1312_nl[21:0];
  assign nl_MultLoop_acc_1311_nl = (MultLoop_acc_1312_nl) + z_out_825;
  assign MultLoop_acc_1311_nl = nl_MultLoop_acc_1311_nl[21:0];
  assign nl_MultLoop_acc_1310_nl = (MultLoop_acc_1311_nl) + z_out_472;
  assign MultLoop_acc_1310_nl = nl_MultLoop_acc_1310_nl[21:0];
  assign nl_MultLoop_acc_1315_nl = z_out_238 + z_out_237;
  assign MultLoop_acc_1315_nl = nl_MultLoop_acc_1315_nl[21:0];
  assign nl_MultLoop_acc_1316_nl = z_out_246 + MultLoop_acc_714_itm;
  assign MultLoop_acc_1316_nl = nl_MultLoop_acc_1316_nl[21:0];
  assign nl_MultLoop_acc_1309_nl = (MultLoop_acc_1310_nl) + MultLoop_acc_758_itm
      + (MultLoop_acc_1315_nl) + (MultLoop_acc_1316_nl);
  assign MultLoop_acc_1309_nl = nl_MultLoop_acc_1309_nl[21:0];
  assign MultLoop_mux1h_347_nl = MUX1HOT_v_22_7_2(z_out_199, z_out_279, z_out_301,
      z_out_197, z_out_276, z_out_507, (MultLoop_acc_1309_nl), {(fsm_output[5]) ,
      (fsm_output[7]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[8])});
  assign nl_z_out_213 = (MultLoop_mux1h_346_nl) + (MultLoop_mux1h_347_nl);
  assign z_out_213 = nl_z_out_213[21:0];
  assign MultLoop_or_81_cse = (fsm_output[5]) | (fsm_output[1]);
  assign MultLoop_mux1h_348_nl = MUX1HOT_v_22_7_2(z_out_200, z_out_201, MultLoop_acc_36_itm,
      z_out_268, z_out_451, z_out_457, z_out_482, {MultLoop_or_81_cse , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[8])});
  assign MultLoop_mux1h_349_nl = MUX1HOT_v_22_6_2(z_out_201, z_out_200, z_out_268,
      z_out_279, z_out_478, z_out_233, {MultLoop_or_81_cse , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_214 = (MultLoop_mux1h_348_nl) + (MultLoop_mux1h_349_nl);
  assign z_out_214 = nl_z_out_214[21:0];
  assign MultLoop_mux1h_350_nl = MUX1HOT_v_22_6_2(z_out_447, z_out_209, z_out_204,
      z_out_202, z_out_268, z_out_505, {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1317_nl = z_out_155_28_7 + z_out_654_28_7;
  assign MultLoop_acc_1317_nl = nl_MultLoop_acc_1317_nl[21:0];
  assign nl_MultLoop_acc_1318_nl = z_out_60_28_7 + z_out_56_28_7;
  assign MultLoop_acc_1318_nl = nl_MultLoop_acc_1318_nl[21:0];
  assign MultLoop_mux1h_351_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1317_nl), z_out_282,
      z_out_207, z_out_199, (MultLoop_acc_1318_nl), z_out_220, {(fsm_output[3]) ,
      (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_215 = (MultLoop_mux1h_350_nl) + (MultLoop_mux1h_351_nl);
  assign z_out_215 = nl_z_out_215[21:0];
  assign nl_MultLoop_acc_1319_nl = z_out_123_28_7 + z_out_126_28_7;
  assign MultLoop_acc_1319_nl = nl_MultLoop_acc_1319_nl[21:0];
  assign nl_MultLoop_acc_1320_nl = z_out_90_28_7 + z_out_66_28_7;
  assign MultLoop_acc_1320_nl = nl_MultLoop_acc_1320_nl[21:0];
  assign MultLoop_mux1h_352_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1319_nl), z_out_201,
      z_out_441, (MultLoop_acc_1320_nl), z_out_301, z_out_496, {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1321_nl = z_out_127_28_7 + z_out_76_28_7;
  assign MultLoop_acc_1321_nl = nl_MultLoop_acc_1321_nl[21:0];
  assign nl_MultLoop_acc_1322_nl = z_out_184_28_7 + z_out_634_28_7;
  assign MultLoop_acc_1322_nl = nl_MultLoop_acc_1322_nl[21:0];
  assign nl_MultLoop_acc_1323_nl = z_out_119_28_7 + z_out_120_28_7;
  assign MultLoop_acc_1323_nl = nl_MultLoop_acc_1323_nl[21:0];
  assign MultLoop_mux1h_353_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1321_nl), z_out_200,
      (MultLoop_acc_1322_nl), (MultLoop_acc_1323_nl), z_out_287, z_out_211, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_216 = (MultLoop_mux1h_352_nl) + (MultLoop_mux1h_353_nl);
  assign z_out_216 = nl_z_out_216[21:0];
  assign MultLoop_mux1h_354_nl = MUX1HOT_v_22_3_2(z_out_438, z_out_195, z_out_451,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_355_nl = MUX1HOT_v_22_3_2(z_out_442, z_out_194, z_out_452,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_217 = (MultLoop_mux1h_354_nl) + (MultLoop_mux1h_355_nl);
  assign z_out_217 = nl_z_out_217[21:0];
  assign MultLoop_mux1h_356_nl = MUX1HOT_v_22_3_2(z_out_831, z_out_220, z_out_477,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_MultLoop_mux_10_nl = MUX_v_22_2_2(z_out_479, z_out_211, fsm_output[1]);
  assign nl_z_out_218 = (MultLoop_mux1h_356_nl) + (MultLoop_MultLoop_mux_10_nl);
  assign z_out_218 = nl_z_out_218[21:0];
  assign MultLoop_mux1h_357_nl = MUX1HOT_v_22_3_2(z_out_507, z_out_442, z_out_468,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_MultLoop_mux_11_nl = MUX_v_22_2_2(z_out_451, z_out_478, fsm_output[5]);
  assign nl_z_out_219 = (MultLoop_mux1h_357_nl) + (MultLoop_MultLoop_mux_11_nl);
  assign z_out_219 = nl_z_out_219[21:0];
  assign nl_MultLoop_acc_1325_nl = z_out_263 + z_out_283;
  assign MultLoop_acc_1325_nl = nl_MultLoop_acc_1325_nl[21:0];
  assign nl_MultLoop_acc_1324_nl = (MultLoop_acc_1325_nl) + z_out_473;
  assign MultLoop_acc_1324_nl = nl_MultLoop_acc_1324_nl[21:0];
  assign MultLoop_mux1h_358_nl = MUX1HOT_v_22_6_2(z_out_65_28_7, z_out_107_28_7,
      z_out_632_28_7, z_out_109_28_7, MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      (MultLoop_acc_1324_nl), {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1326_nl = z_out_476 + MultLoop_acc_885_itm;
  assign MultLoop_acc_1326_nl = nl_MultLoop_acc_1326_nl[21:0];
  assign MultLoop_mux1h_359_nl = MUX1HOT_v_22_6_2(z_out_87_28_7, z_out_112_28_7,
      z_out_660_28_7, z_out_107_28_7, z_out_135_28_7, (MultLoop_acc_1326_nl), {(fsm_output[3])
      , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_220 = (MultLoop_mux1h_358_nl) + (MultLoop_mux1h_359_nl);
  assign z_out_220 = nl_z_out_220[21:0];
  assign MultLoop_mux1h_360_nl = MUX1HOT_v_22_5_2(z_out_111_28_7, z_out_77_28_7,
      z_out_53_28_7, z_out_142_28_7, z_out_535, {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1335_nl = z_out_128_28_7 + z_out_117_28_7;
  assign MultLoop_acc_1335_nl = nl_MultLoop_acc_1335_nl[21:0];
  assign nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9559:9552]));
  assign MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1336_nl = z_out_154_28_7 + (readslicef_29_22_7((MultLoop_1195_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1336_nl = nl_MultLoop_acc_1336_nl[21:0];
  assign nl_MultLoop_acc_1331_nl = MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_164_28_7;
  assign MultLoop_acc_1331_nl = nl_MultLoop_acc_1331_nl[21:0];
  assign nl_MultLoop_acc_1332_nl = z_out_150_28_7 + z_out_179_28_7;
  assign MultLoop_acc_1332_nl = nl_MultLoop_acc_1332_nl[21:0];
  assign nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9567:9560]));
  assign MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9575:9568]));
  assign MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1338_nl = (readslicef_29_22_7((MultLoop_1196_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1197_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1338_nl = nl_MultLoop_acc_1338_nl[21:0];
  assign nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9583:9576]));
  assign MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9591:9584]));
  assign MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1339_nl = (readslicef_29_22_7((MultLoop_1198_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1199_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1339_nl = nl_MultLoop_acc_1339_nl[21:0];
  assign nl_MultLoop_acc_1328_nl = MultLoop_acc_102_itm + (MultLoop_acc_1335_nl)
      + (MultLoop_acc_1336_nl) + (MultLoop_acc_1331_nl) + (MultLoop_acc_1332_nl)
      + (MultLoop_acc_1338_nl) + (MultLoop_acc_1339_nl);
  assign MultLoop_acc_1328_nl = nl_MultLoop_acc_1328_nl[21:0];
  assign nl_MultLoop_acc_1327_nl = (MultLoop_acc_1328_nl) + z_out_543;
  assign MultLoop_acc_1327_nl = nl_MultLoop_acc_1327_nl[21:0];
  assign MultLoop_mux1h_361_nl = MUX1HOT_v_22_5_2(z_out_108_28_7, z_out_92_28_7,
      z_out_48_28_7, z_out_144_28_7, (MultLoop_acc_1327_nl), {(fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_221 = (MultLoop_mux1h_360_nl) + (MultLoop_mux1h_361_nl);
  assign z_out_221 = nl_z_out_221[21:0];
  assign MultLoop_mux1h_362_nl = MUX1HOT_v_22_3_2(z_out_441, z_out_506, z_out_457,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_363_nl = MUX1HOT_v_22_3_2(z_out_447, z_out_507, z_out_482,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_222 = (MultLoop_mux1h_362_nl) + (MultLoop_mux1h_363_nl);
  assign z_out_222 = nl_z_out_222[21:0];
  assign MultLoop_mux_78_nl = MUX_v_22_2_2(z_out_303, z_out_202, fsm_output[3]);
  assign MultLoop_mux_79_nl = MUX_v_22_2_2(z_out_298, z_out_208, fsm_output[3]);
  assign nl_z_out_223 = (MultLoop_mux_78_nl) + (MultLoop_mux_79_nl);
  assign z_out_223 = nl_z_out_223[21:0];
  assign MultLoop_MultLoop_mux_12_nl = MUX_v_22_2_2(z_out_497, z_out_468, fsm_output[4]);
  assign MultLoop_MultLoop_mux_13_nl = MUX_v_22_2_2(z_out_495, z_out_452, fsm_output[4]);
  assign nl_z_out_224 = (MultLoop_MultLoop_mux_12_nl) + (MultLoop_MultLoop_mux_13_nl);
  assign z_out_224 = nl_z_out_224[21:0];
  assign MultLoop_mux1h_364_nl = MUX1HOT_v_22_3_2(z_out_233, z_out_194, z_out_507,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4])});
  assign MultLoop_mux1h_365_nl = MUX1HOT_v_22_3_2(z_out_279, z_out_468, z_out_495,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[4])});
  assign nl_z_out_225 = (MultLoop_mux1h_364_nl) + (MultLoop_mux1h_365_nl);
  assign z_out_225 = nl_z_out_225[21:0];
  assign nl_MultLoop_acc_1340_nl = z_out_133_28_7 + z_out_125_28_7;
  assign MultLoop_acc_1340_nl = nl_MultLoop_acc_1340_nl[21:0];
  assign MultLoop_mux1h_366_nl = MUX1HOT_v_22_3_2((MultLoop_acc_1340_nl), z_out_211,
      MultLoop_acc_689_itm, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_367_nl = MUX1HOT_v_22_3_2(z_out_446, z_out_210, z_out_447,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_226 = (MultLoop_mux1h_366_nl) + (MultLoop_mux1h_367_nl);
  assign z_out_226 = nl_z_out_226[21:0];
  assign AccumDotWidth_mux1h_762_nl = MUX1HOT_v_22_4_2(z_out_740, z_out_539, z_out_755,
      z_out_325, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_763_nl = MUX1HOT_v_22_4_2(z_out_396, z_out_529, z_out_759,
      MultLoop_acc_470_itm, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_227 = (AccumDotWidth_mux1h_762_nl) + (AccumDotWidth_mux1h_763_nl);
  assign z_out_227 = nl_z_out_227[21:0];
  assign AccumDotWidth_mux1h_764_nl = MUX1HOT_v_22_5_2(z_out_734, z_out_543, z_out_756,
      z_out_330, z_out_512, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_765_nl = MUX1HOT_v_22_5_2(z_out_739, z_out_508, z_out_538,
      z_out_531, z_out_239, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_228 = (AccumDotWidth_mux1h_764_nl) + (AccumDotWidth_mux1h_765_nl);
  assign z_out_228 = nl_z_out_228[21:0];
  assign nl_MultLoop_acc_1341_nl = (z_out_1105_29_7[21:0]) + (z_out_1102_29_7[21:0]);
  assign MultLoop_acc_1341_nl = nl_MultLoop_acc_1341_nl[21:0];
  assign AccumDotWidth_mux1h_766_nl = MUX1HOT_v_22_7_2(z_out_264, z_out_850, z_out_844,
      AccumDotWidth_acc_1300_itm, z_out_754, z_out_307, (MultLoop_acc_1341_nl), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_767_nl = MUX1HOT_v_22_7_2(z_out_263, z_out_778, z_out_835,
      z_out_256, z_out_536, z_out_283, z_out_314, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_229 = (AccumDotWidth_mux1h_766_nl) + (AccumDotWidth_mux1h_767_nl);
  assign z_out_229 = nl_z_out_229[21:0];
  assign MultLoop_mux_80_nl = MUX_v_22_2_2(z_out_452, z_out_478, fsm_output[4]);
  assign MultLoop_mux_81_nl = MUX_v_22_2_2(z_out_233, z_out_477, fsm_output[4]);
  assign nl_z_out_230 = (MultLoop_mux_80_nl) + (MultLoop_mux_81_nl);
  assign z_out_230 = nl_z_out_230[21:0];
  assign MultLoop_mux_82_nl = MUX_v_22_2_2(z_out_291, z_out_194, fsm_output[3]);
  assign MultLoop_mux_83_nl = MUX_v_22_2_2(z_out_293, z_out_200, fsm_output[3]);
  assign nl_z_out_231 = (MultLoop_mux_82_nl) + (MultLoop_mux_83_nl);
  assign z_out_231 = nl_z_out_231[21:0];
  assign MultLoop_mux1h_368_nl = MUX1HOT_v_22_3_2(z_out_306, z_out_465, z_out_506,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_369_nl = MUX1HOT_v_22_3_2(z_out_279, z_out_485, z_out_497,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_232 = (MultLoop_mux1h_368_nl) + (MultLoop_mux1h_369_nl);
  assign z_out_232 = nl_z_out_232[21:0];
  assign nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1932_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[703:696]));
  assign MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1937_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[711:704]));
  assign MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1346_nl = (readslicef_29_22_7((MultLoop_88_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_89_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1346_nl = nl_MultLoop_acc_1346_nl[21:0];
  assign nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1945_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[719:712]));
  assign MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0]))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[727:720]));
  assign MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1347_nl = (readslicef_29_22_7((MultLoop_90_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_91_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1347_nl = nl_MultLoop_acc_1347_nl[21:0];
  assign nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0]))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[735:728]));
  assign MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[743:736]));
  assign MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1349_nl = (readslicef_29_22_7((MultLoop_92_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_93_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1349_nl = nl_MultLoop_acc_1349_nl[21:0];
  assign nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[751:744]));
  assign MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[759:752]));
  assign MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1350_nl = (readslicef_29_22_7((MultLoop_94_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_95_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1350_nl = nl_MultLoop_acc_1350_nl[21:0];
  assign nl_MultLoop_acc_1344_nl = (MultLoop_acc_1346_nl) + (MultLoop_acc_1347_nl)
      + (MultLoop_acc_1349_nl) + (MultLoop_acc_1350_nl);
  assign MultLoop_acc_1344_nl = nl_MultLoop_acc_1344_nl[21:0];
  assign nl_MultLoop_acc_1343_nl = z_out_454 + (MultLoop_acc_1344_nl);
  assign MultLoop_acc_1343_nl = nl_MultLoop_acc_1343_nl[21:0];
  assign nl_MultLoop_acc_1342_nl = z_out_538 + (MultLoop_acc_1343_nl);
  assign MultLoop_acc_1342_nl = nl_MultLoop_acc_1342_nl[21:0];
  assign MultLoop_mux1h_370_nl = MUX1HOT_v_22_5_2(z_out_133_28_7, z_out_102_28_7,
      z_out_643_28_7, z_out_143_28_7, (MultLoop_acc_1342_nl), {(fsm_output[5]) ,
      (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0))
      * $signed((w4_rsci_idat_mxwt[4055:4048]));
  assign MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1355_nl = z_out_151_28_7 + MultLoop_99_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1355_nl = nl_MultLoop_acc_1355_nl[21:0];
  assign nl_MultLoop_acc_1354_nl = z_out_561 + (MultLoop_acc_1355_nl);
  assign MultLoop_acc_1354_nl = nl_MultLoop_acc_1354_nl[21:0];
  assign nl_MultLoop_acc_1353_nl = (MultLoop_acc_1354_nl) + z_out_206;
  assign MultLoop_acc_1353_nl = nl_MultLoop_acc_1353_nl[21:0];
  assign nl_MultLoop_acc_1351_nl = MultLoop_acc_1266_itm + (MultLoop_acc_1353_nl)
      + z_out_460;
  assign MultLoop_acc_1351_nl = nl_MultLoop_acc_1351_nl[21:0];
  assign MultLoop_mux1h_371_nl = MUX1HOT_v_22_5_2(z_out_136_28_7, z_out_94_28_7,
      (readslicef_29_22_7((MultLoop_507_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      z_out_140_28_7, (MultLoop_acc_1351_nl), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_233 = (MultLoop_mux1h_370_nl) + (MultLoop_mux1h_371_nl);
  assign z_out_233 = nl_z_out_233[21:0];
  assign AccumDotWidth_mux1h_768_nl = MUX1HOT_v_22_7_2(z_out_314, z_out_849, z_out_851,
      z_out_311, z_out_370, z_out_850, MultLoop_868_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_769_nl = MUX1HOT_v_22_6_2(z_out_315, z_out_848, z_out_778,
      z_out_245, z_out_366, (z_out_939_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_234 = (AccumDotWidth_mux1h_768_nl) + (AccumDotWidth_mux1h_769_nl);
  assign z_out_234 = nl_z_out_234[21:0];
  assign AccumDotWidth_mux1h_770_nl = MUX1HOT_v_22_7_2(z_out_308, z_out_849, z_out_503,
      z_out_316, z_out_365, z_out_311, (z_out_935_29_7[21:0]), {(fsm_output[1]) ,
      operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_771_nl = MUX1HOT_v_22_8_2(z_out_316, AccumDotWidth_acc_1220_itm,
      AccumDotWidth_acc_1218_itm, z_out_850, z_out_849, z_out_352, z_out_244, MultLoop_483_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_235 = (AccumDotWidth_mux1h_770_nl) + (AccumDotWidth_mux1h_771_nl);
  assign z_out_235 = nl_z_out_235[21:0];
  assign nl_AccumDotWidth_acc_2401_nl = z_out_545 + z_out_346;
  assign AccumDotWidth_acc_2401_nl = nl_AccumDotWidth_acc_2401_nl[21:0];
  assign AccumDotWidth_mux1h_772_nl = MUX1HOT_v_22_8_2(z_out_310, z_out_377, z_out_807,
      z_out_557, (AccumDotWidth_acc_2401_nl), z_out_362, z_out_316, z_out_253, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_773_nl = MUX1HOT_v_22_8_2(z_out_850, z_out_380, z_out_687,
      z_out_556, z_out_315, z_out_367, z_out_308, z_out_244, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_236 = (AccumDotWidth_mux1h_772_nl) + (AccumDotWidth_mux1h_773_nl);
  assign z_out_236 = nl_z_out_236[21:0];
  assign AccumDotWidth_or_145_cse = (fsm_output[4]) | (fsm_output[6]);
  assign AccumDotWidth_mux1h_774_nl = MUX1HOT_v_22_7_2(z_out_412, z_out_842, z_out_491,
      z_out_267, z_out_531, z_out_245, z_out_234, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1356_nl = (z_out_947_29_7[21:0]) + (z_out_948_29_7[21:0]);
  assign MultLoop_acc_1356_nl = nl_MultLoop_acc_1356_nl[21:0];
  assign AccumDotWidth_mux1h_775_nl = MUX1HOT_v_22_8_2(z_out_413, z_out_836, AccumDotWidth_acc_1235_itm,
      z_out_271, z_out_265, z_out_795, z_out_266, (MultLoop_acc_1356_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_237 = (AccumDotWidth_mux1h_774_nl) + (AccumDotWidth_mux1h_775_nl);
  assign z_out_237 = nl_z_out_237[21:0];
  assign nl_MultLoop_acc_1357_nl = (z_out_1186_29_7[21:0]) + (z_out_952_29_7[21:0]);
  assign MultLoop_acc_1357_nl = nl_MultLoop_acc_1357_nl[21:0];
  assign AccumDotWidth_mux1h_776_nl = MUX1HOT_v_22_4_2(z_out_315, z_out_314, z_out_816,
      (MultLoop_acc_1357_nl), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_777_nl = MUX1HOT_v_22_4_2(z_out_313, z_out_310, z_out_852,
      z_out_254, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_238 = (AccumDotWidth_mux1h_776_nl) + (AccumDotWidth_mux1h_777_nl);
  assign z_out_238 = nl_z_out_238[21:0];
  assign nl_MultLoop_acc_1358_nl = (z_out_1095_29_7[21:0]) + (z_out_1092_29_7[21:0]);
  assign MultLoop_acc_1358_nl = nl_MultLoop_acc_1358_nl[21:0];
  assign AccumDotWidth_mux_84_nl = MUX_v_22_2_2(z_out_528, (MultLoop_acc_1358_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1359_nl = (z_out_1080_29_7[21:0]) + (z_out_1131_29_7[21:0]);
  assign MultLoop_acc_1359_nl = nl_MultLoop_acc_1359_nl[21:0];
  assign AccumDotWidth_mux_85_nl = MUX_v_22_2_2(z_out_307, (MultLoop_acc_1359_nl),
      fsm_output[8]);
  assign nl_z_out_239 = (AccumDotWidth_mux_84_nl) + (AccumDotWidth_mux_85_nl);
  assign z_out_239 = nl_z_out_239[21:0];
  assign nl_MultLoop_acc_1360_nl = (z_out_983_29_7[21:0]) + (z_out_982_29_7[21:0]);
  assign MultLoop_acc_1360_nl = nl_MultLoop_acc_1360_nl[21:0];
  assign AccumDotWidth_mux1h_778_nl = MUX1HOT_v_22_3_2(z_out_526, z_out_274, (MultLoop_acc_1360_nl),
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1361_nl = (z_out_981_29_7[21:0]) + (z_out_980_29_7[21:0]);
  assign MultLoop_acc_1361_nl = nl_MultLoop_acc_1361_nl[21:0];
  assign AccumDotWidth_mux1h_779_nl = MUX1HOT_v_22_3_2(z_out_274, z_out_806, (MultLoop_acc_1361_nl),
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_240 = (AccumDotWidth_mux1h_778_nl) + (AccumDotWidth_mux1h_779_nl);
  assign z_out_240 = nl_z_out_240[21:0];
  assign nl_MultLoop_acc_1362_nl = (z_out_1103_29_7[21:0]) + (z_out_1101_29_7[21:0]);
  assign MultLoop_acc_1362_nl = nl_MultLoop_acc_1362_nl[21:0];
  assign AccumDotWidth_mux1h_780_nl = MUX1HOT_v_22_6_2(z_out_804, z_out_274, z_out_529,
      z_out_737, z_out_826, (MultLoop_acc_1362_nl), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1363_nl = (z_out_1099_29_7[21:0]) + (z_out_1027_29_7[21:0]);
  assign MultLoop_acc_1363_nl = nl_MultLoop_acc_1363_nl[21:0];
  assign AccumDotWidth_mux1h_781_nl = MUX1HOT_v_22_6_2(z_out_806, z_out_307, z_out_273,
      z_out_739, z_out_851, (MultLoop_acc_1363_nl), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_241 = (AccumDotWidth_mux1h_780_nl) + (AccumDotWidth_mux1h_781_nl);
  assign z_out_241 = nl_z_out_241[21:0];
  assign AccumDotWidth_mux1h_782_nl = MUX1HOT_v_22_4_2(z_out_804, z_out_802, z_out_736,
      z_out_314, {AccumDotWidth_or_132_cse_1 , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_783_nl = MUX1HOT_v_22_5_2(z_out_802, z_out_680, z_out_805,
      z_out_734, z_out_312, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_242 = (AccumDotWidth_mux1h_782_nl) + (AccumDotWidth_mux1h_783_nl);
  assign z_out_242 = nl_z_out_242[21:0];
  assign AccumDotWidth_mux_86_nl = MUX_v_22_2_2(z_out_266, z_out_255, fsm_output[8]);
  assign AccumDotWidth_mux_87_nl = MUX_v_22_2_2(z_out_275, z_out_307, fsm_output[8]);
  assign nl_z_out_243 = (AccumDotWidth_mux_86_nl) + (AccumDotWidth_mux_87_nl);
  assign z_out_243 = nl_z_out_243[21:0];
  assign nl_AccumDotWidth_acc_2402_nl = conv_s2s_21_22(z_out_1176_29_7[22:2]) + conv_s2s_21_22(z_out_1073_29_7[22:2]);
  assign AccumDotWidth_acc_2402_nl = nl_AccumDotWidth_acc_2402_nl[21:0];
  assign AccumDotWidth_mux1h_784_nl = MUX1HOT_v_22_6_2(z_out_791, z_out_391, z_out_722,
      z_out_738, (AccumDotWidth_acc_2402_nl), (z_out_945_29_7[21:0]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2403_nl = conv_s2s_21_22(z_out_879_29_7[22:2]) + conv_s2s_21_22(z_out_1030_29_7[22:2]);
  assign AccumDotWidth_acc_2403_nl = nl_AccumDotWidth_acc_2403_nl[21:0];
  assign AccumDotWidth_mux1h_785_nl = MUX1HOT_v_22_6_2(AccumDotWidth_acc_1203_itm,
      z_out_393, z_out_713, z_out_735, (AccumDotWidth_acc_2403_nl), (z_out_944_29_7[21:0]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_244 = (AccumDotWidth_mux1h_784_nl) + (AccumDotWidth_mux1h_785_nl);
  assign z_out_244 = nl_z_out_244[21:0];
  assign AccumDotWidth_mux1h_786_nl = MUX1HOT_v_22_6_2(z_out_309, z_out_389, z_out_689,
      z_out_732, z_out_363, (z_out_579_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_787_nl = MUX1HOT_v_22_6_2(AccumDotWidth_acc_1186_itm,
      z_out_390, z_out_682, z_out_707, z_out_359, (z_out_582_29_7[21:0]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_245 = (AccumDotWidth_mux1h_786_nl) + (AccumDotWidth_mux1h_787_nl);
  assign z_out_245 = nl_z_out_245[21:0];
  assign nl_MultLoop_acc_1364_nl = (z_out_949_29_7[21:0]) + (z_out_905_29_7[21:0]);
  assign MultLoop_acc_1364_nl = nl_MultLoop_acc_1364_nl[21:0];
  assign AccumDotWidth_mux_88_nl = MUX_v_22_2_2(z_out_517, (MultLoop_acc_1364_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1365_nl = (z_out_903_29_7[21:0]) + (z_out_902_29_7[21:0]);
  assign MultLoop_acc_1365_nl = nl_MultLoop_acc_1365_nl[21:0];
  assign AccumDotWidth_mux_89_nl = MUX_v_22_2_2(z_out_263, (MultLoop_acc_1365_nl),
      fsm_output[8]);
  assign nl_z_out_246 = (AccumDotWidth_mux_88_nl) + (AccumDotWidth_mux_89_nl);
  assign z_out_246 = nl_z_out_246[21:0];
  assign AccumDotWidth_mux1h_788_nl = MUX1HOT_v_22_4_2(z_out_367, z_out_729, z_out_699,
      MultLoop_612_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_789_nl = MUX1HOT_v_22_4_2(z_out_370, z_out_728, z_out_697,
      (z_out_900_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_247 = (AccumDotWidth_mux1h_788_nl) + (AccumDotWidth_mux1h_789_nl);
  assign z_out_247 = nl_z_out_247[21:0];
  assign AccumDotWidth_mux_90_nl = MUX_v_22_2_2(z_out_487, (z_out_1079_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_91_nl = MUX_v_22_2_2(MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      MultLoop_577_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      fsm_output[8]);
  assign nl_z_out_248 = (AccumDotWidth_mux_90_nl) + (AccumDotWidth_mux_91_nl);
  assign z_out_248 = nl_z_out_248[21:0];
  assign nl_AccumDotWidth_acc_2404_nl = conv_s2s_21_22(z_out_1163_29_7[22:2]) + conv_s2s_21_22(z_out_996_29_7[22:2]);
  assign AccumDotWidth_acc_2404_nl = nl_AccumDotWidth_acc_2404_nl[21:0];
  assign AccumDotWidth_mux1h_790_nl = MUX1HOT_v_22_5_2(z_out_403, (AccumDotWidth_acc_2404_nl),
      z_out_727, z_out_360, ({MultLoop_acc_1283_psp , (AccumDotWidth_acc_1837_itm[10:0])}),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_791_nl = MUX1HOT_v_22_5_2(z_out_400, z_out_375, z_out_726,
      z_out_358, (z_out_910_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_249 = (AccumDotWidth_mux1h_790_nl) + (AccumDotWidth_mux1h_791_nl);
  assign z_out_249 = nl_z_out_249[21:0];
  assign AccumDotWidth_mux1h_792_nl = MUX1HOT_v_22_6_2(z_out_545, z_out_491, z_out_555,
      z_out_746, z_out_546, (z_out_1035_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_793_nl = MUX1HOT_v_22_6_2(z_out_340, z_out_341, z_out_331,
      z_out_744, z_out_339, MultLoop_705_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_250 = (AccumDotWidth_mux1h_792_nl) + (AccumDotWidth_mux1h_793_nl);
  assign z_out_250 = nl_z_out_250[21:0];
  assign AccumDotWidth_mux1h_794_nl = MUX1HOT_v_22_7_2(z_out_503, z_out_430, z_out_433,
      z_out_371, z_out_741, z_out_492, ({MultLoop_acc_1284_psp , (AccumDotWidth_acc_1845_itm[10:0])}),
      {MultLoop_or_81_cse , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_795_nl = MUX1HOT_v_22_8_2(z_out_341, z_out_405, z_out_424,
      z_out_367, z_out_407, z_out_749, z_out_342, (z_out_971_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_251 = (AccumDotWidth_mux1h_794_nl) + (AccumDotWidth_mux1h_795_nl);
  assign z_out_251 = nl_z_out_251[21:0];
  assign AccumDotWidth_mux1h_796_nl = MUX1HOT_v_22_6_2(z_out_726, z_out_488, z_out_310,
      z_out_693, z_out_494, MultLoop_484_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_797_nl = MUX1HOT_v_22_6_2(z_out_729, z_out_339, z_out_314,
      z_out_742, z_out_341, (z_out_1037_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_252 = (AccumDotWidth_mux1h_796_nl) + (AccumDotWidth_mux1h_797_nl);
  assign z_out_252 = nl_z_out_252[21:0];
  assign AccumDotWidth_mux1h_798_nl = MUX1HOT_v_22_4_2(z_out_378, AccumDotWidth_acc_1164_itm,
      z_out_695, ({MultLoop_acc_1282_psp , (AccumDotWidth_acc_1426_itm[10:0])}),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2405_nl = conv_s2s_21_22(z_out_884_29_7[22:2]) + conv_s2s_21_22(z_out_1098_29_7[22:2]);
  assign AccumDotWidth_acc_2405_nl = nl_AccumDotWidth_acc_2405_nl[21:0];
  assign AccumDotWidth_mux1h_799_nl = MUX1HOT_v_22_4_2((AccumDotWidth_acc_2405_nl),
      z_out_427, z_out_694, (z_out_946_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_253 = (AccumDotWidth_mux1h_798_nl) + (AccumDotWidth_mux1h_799_nl);
  assign z_out_253 = nl_z_out_253[21:0];
  assign AccumDotWidth_mux1h_800_nl = MUX1HOT_v_22_6_2(z_out_727, z_out_489, z_out_567,
      z_out_696, z_out_500, (z_out_966_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_801_nl = MUX1HOT_v_22_6_2(z_out_724, z_out_347, z_out_336,
      z_out_698, z_out_489, MultLoop_867_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_254 = (AccumDotWidth_mux1h_800_nl) + (AccumDotWidth_mux1h_801_nl);
  assign z_out_254 = nl_z_out_254[21:0];
  assign AccumDotWidth_or_149_cse = (fsm_output[1]) | (fsm_output[7]);
  assign AccumDotWidth_mux1h_802_nl = MUX1HOT_v_22_6_2(z_out_489, z_out_461, z_out_500,
      z_out_700, z_out_490, (z_out_1104_29_7[21:0]), {nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_803_nl = MUX1HOT_v_22_6_2(z_out_345, z_out_343, z_out_340,
      z_out_329, z_out_692, MultLoop_833_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {AccumDotWidth_or_149_cse , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_255 = (AccumDotWidth_mux1h_802_nl) + (AccumDotWidth_mux1h_803_nl);
  assign z_out_255 = nl_z_out_255[21:0];
  assign AccumDotWidth_mux1h_804_nl = MUX1HOT_v_22_8_2(z_out_500, z_out_407, z_out_432,
      z_out_503, z_out_554, z_out_351, z_out_483, ({MultLoop_acc_1281_psp , (AccumDotWidth_acc_1135_itm[10:0])}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_805_nl = MUX1HOT_v_22_8_2(z_out_343, z_out_402, z_out_434,
      z_out_349, z_out_553, z_out_353, z_out_331, (z_out_607_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_256 = (AccumDotWidth_mux1h_804_nl) + (AccumDotWidth_mux1h_805_nl);
  assign z_out_256 = nl_z_out_256[21:0];
  assign AccumDotWidth_mux1h_806_nl = MUX1HOT_v_22_6_2(z_out_728, z_out_366, z_out_494,
      z_out_747, z_out_484, MultLoop_996_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_807_nl = MUX1HOT_v_22_6_2(z_out_723, z_out_724, z_out_484,
      z_out_743, z_out_343, (z_out_1016_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_257 = (AccumDotWidth_mux1h_806_nl) + (AccumDotWidth_mux1h_807_nl);
  assign z_out_257 = nl_z_out_257[21:0];
  assign nl_AccumDotWidth_acc_2406_nl = conv_s2s_21_22(z_out_1013_29_7[22:2]) + conv_s2s_21_22(z_out_874_29_7[22:2]);
  assign AccumDotWidth_acc_2406_nl = nl_AccumDotWidth_acc_2406_nl[21:0];
  assign AccumDotWidth_mux1h_808_nl = MUX1HOT_v_22_5_2(z_out_401, (AccumDotWidth_acc_2406_nl),
      z_out_731, z_out_359, AccumDotWidth_acc_1326_itm, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2407_nl = conv_s2s_21_22(z_out_886_29_7[22:2]) + conv_s2s_21_22(z_out_1100_29_7[22:2]);
  assign AccumDotWidth_acc_2407_nl = nl_AccumDotWidth_acc_2407_nl[21:0];
  assign AccumDotWidth_mux1h_809_nl = MUX1HOT_v_22_5_2(z_out_404, (AccumDotWidth_acc_2407_nl),
      z_out_730, z_out_356, (z_out_874_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_258 = (AccumDotWidth_mux1h_808_nl) + (AccumDotWidth_mux1h_809_nl);
  assign z_out_258 = nl_z_out_258[21:0];
  assign AccumDotWidth_mux1h_810_nl = MUX1HOT_v_22_5_2(z_out_423, z_out_492, z_out_805,
      z_out_461, (z_out_891_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_811_nl = MUX1HOT_v_22_5_2(z_out_435, z_out_342, z_out_804,
      z_out_347, MultLoop_235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_259 = (AccumDotWidth_mux1h_810_nl) + (AccumDotWidth_mux1h_811_nl);
  assign z_out_259 = nl_z_out_259[21:0];
  assign AccumDotWidth_mux1h_812_nl = MUX1HOT_v_22_6_2(z_out_402, z_out_490, z_out_493,
      z_out_691, z_out_488, MultLoop_228_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_813_nl = MUX1HOT_v_22_6_2(z_out_401, z_out_345, z_out_490,
      z_out_690, z_out_344, (z_out_926_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_260 = (AccumDotWidth_mux1h_812_nl) + (AccumDotWidth_mux1h_813_nl);
  assign z_out_260 = nl_z_out_260[21:0];
  assign AccumDotWidth_or_150_cse = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[7]);
  assign AccumDotWidth_mux1h_814_nl = MUX1HOT_v_22_5_2(z_out_493, z_out_376, z_out_492,
      z_out_745, (z_out_925_29_7[21:0]), {AccumDotWidth_or_150_cse , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_815_nl = MUX1HOT_v_22_7_2(z_out_340, z_out_377, z_out_343,
      z_out_488, z_out_750, z_out_503, MultLoop_227_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_261 = (AccumDotWidth_mux1h_814_nl) + (AccumDotWidth_mux1h_815_nl);
  assign z_out_261 = nl_z_out_261[21:0];
  assign AccumDotWidth_or_151_nl = (fsm_output[1]) | (fsm_output[5]) | (fsm_output[7]);
  assign AccumDotWidth_mux1h_816_nl = MUX1HOT_v_22_4_2(z_out_491, z_out_549, z_out_494,
      z_out_555, {(AccumDotWidth_or_151_nl) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[8])});
  assign nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[655:648]));
  assign MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[663:656]));
  assign MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1366_nl = (readslicef_29_22_7((MultLoop_82_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_83_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1366_nl = nl_MultLoop_acc_1366_nl[21:0];
  assign AccumDotWidth_mux1h_817_nl = MUX1HOT_v_22_6_2(z_out_342, z_out_350, z_out_351,
      z_out_489, z_out_340, (MultLoop_acc_1366_nl), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_262 = (AccumDotWidth_mux1h_816_nl) + (AccumDotWidth_mux1h_817_nl);
  assign z_out_262 = nl_z_out_262[21:0];
  assign AccumDotWidth_or_152_cse = (fsm_output[6:5]!=2'b00);
  assign AccumDotWidth_mux1h_818_nl = MUX1HOT_v_22_8_2(z_out_726, z_out_347, z_out_336,
      z_out_334, z_out_354, z_out_258, z_out_355, z_out_329, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_819_nl = MUX1HOT_v_22_7_2(z_out_722, z_out_353, z_out_335,
      z_out_329, z_out_343, AccumDotWidth_acc_1937_itm, AccumDotWidth_acc_1300_itm,
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_152_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_263 = (AccumDotWidth_mux1h_818_nl) + (AccumDotWidth_mux1h_819_nl);
  assign z_out_263 = nl_z_out_263[21:0];
  assign nl_AccumDotWidth_acc_2408_nl = z_out_805 + z_out_684;
  assign AccumDotWidth_acc_2408_nl = nl_AccumDotWidth_acc_2408_nl[21:0];
  assign nl_MultLoop_acc_1368_nl = (z_out_901_29_7[21:0]) + MultLoop_611_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1368_nl = nl_MultLoop_acc_1368_nl[21:0];
  assign nl_MultLoop_acc_1367_nl = z_out_490 + (MultLoop_acc_1368_nl);
  assign MultLoop_acc_1367_nl = nl_MultLoop_acc_1367_nl[21:0];
  assign AccumDotWidth_mux1h_820_nl = MUX1HOT_v_22_8_2(z_out_723, z_out_339, (AccumDotWidth_acc_2408_nl),
      z_out_338, z_out_685, z_out_249, z_out_709, (MultLoop_acc_1367_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1369_nl = z_out_247 + z_out_488;
  assign MultLoop_acc_1369_nl = nl_MultLoop_acc_1369_nl[21:0];
  assign AccumDotWidth_mux1h_821_nl = MUX1HOT_v_22_8_2(z_out_724, z_out_351, z_out_257,
      z_out_337, z_out_687, z_out_347, z_out_708, (MultLoop_acc_1369_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_264 = (AccumDotWidth_mux1h_820_nl) + (AccumDotWidth_mux1h_821_nl);
  assign z_out_264 = nl_z_out_264[21:0];
  assign nl_AccumDotWidth_acc_2409_nl = z_out_553 + z_out_554;
  assign AccumDotWidth_acc_2409_nl = nl_AccumDotWidth_acc_2409_nl[21:0];
  assign AccumDotWidth_mux1h_822_nl = MUX1HOT_v_22_8_2(z_out_367, z_out_235, z_out_521,
      z_out_336, z_out_393, z_out_525, (AccumDotWidth_acc_2409_nl), z_out_510, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2410_nl = z_out_687 + z_out_728;
  assign AccumDotWidth_acc_2410_nl = nl_AccumDotWidth_acc_2410_nl[21:0];
  assign nl_AccumDotWidth_acc_2411_nl = z_out_686 + z_out_422;
  assign AccumDotWidth_acc_2411_nl = nl_AccumDotWidth_acc_2411_nl[21:0];
  assign AccumDotWidth_mux1h_823_nl = MUX1HOT_v_22_8_2(z_out_366, (AccumDotWidth_acc_2410_nl),
      (AccumDotWidth_acc_2411_nl), z_out_331, z_out_394, z_out_527, z_out_511, AccumDotWidth_acc_1198_itm,
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_265 = (AccumDotWidth_mux1h_822_nl) + (AccumDotWidth_mux1h_823_nl);
  assign z_out_265 = nl_z_out_265[21:0];
  assign nl_MultLoop_acc_1370_nl = z_out_484 + z_out_493;
  assign MultLoop_acc_1370_nl = nl_MultLoop_acc_1370_nl[21:0];
  assign AccumDotWidth_mux1h_824_nl = MUX1HOT_v_22_7_2(z_out_709, z_out_692, z_out_558,
      z_out_723, z_out_532, z_out_353, (MultLoop_acc_1370_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1371_nl = z_out_489 + z_out_491;
  assign MultLoop_acc_1371_nl = nl_MultLoop_acc_1371_nl[21:0];
  assign AccumDotWidth_mux1h_825_nl = MUX1HOT_v_22_7_2(z_out_705, z_out_693, z_out_339,
      z_out_703, z_out_531, z_out_351, (MultLoop_acc_1371_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_266 = (AccumDotWidth_mux1h_824_nl) + (AccumDotWidth_mux1h_825_nl);
  assign z_out_266 = nl_z_out_266[21:0];
  assign AccumDotWidth_or_153_cse = (fsm_output[1]) | (fsm_output[6]);
  assign nl_MultLoop_acc_1372_nl = z_out_462 + z_out_483;
  assign MultLoop_acc_1372_nl = nl_MultLoop_acc_1372_nl[21:0];
  assign AccumDotWidth_mux1h_826_nl = MUX1HOT_v_22_7_2(z_out_391, z_out_563, z_out_732,
      z_out_708, z_out_728, z_out_236, (MultLoop_acc_1372_nl), {(fsm_output[2]) ,
      AccumDotWidth_or_153_cse , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1373_nl = z_out_461 + z_out_494;
  assign MultLoop_acc_1373_nl = nl_MultLoop_acc_1373_nl[21:0];
  assign AccumDotWidth_mux1h_827_nl = MUX1HOT_v_22_8_2(z_out_395, z_out_526, z_out_740,
      z_out_709, z_out_727, z_out_348, z_out_327, (MultLoop_acc_1373_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_267 = (AccumDotWidth_mux1h_826_nl) + (AccumDotWidth_mux1h_827_nl);
  assign z_out_267 = nl_z_out_267[21:0];
  assign MultLoop_mux1h_372_nl = MUX1HOT_v_22_7_2(z_out_118_28_7, z_out_47_28_7,
      z_out_634_28_7, z_out_93_28_7, z_out_51_28_7, z_out_55_28_7, z_out_111_28_7,
      {(fsm_output[7]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[3])});
  assign MultLoop_mux1h_373_nl = MUX1HOT_v_22_7_2(z_out_113_28_7, z_out_40_28_7,
      z_out_639_28_7, z_out_92_28_7, z_out_50_28_7, z_out_46_28_7, z_out_112_28_7,
      {(fsm_output[7]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nl_z_out_268 = (MultLoop_mux1h_372_nl) + (MultLoop_mux1h_373_nl);
  assign z_out_268 = nl_z_out_268[21:0];
  assign AccumDotWidth_mux1h_828_nl = MUX1HOT_v_22_7_2(z_out_368, z_out_236, z_out_321,
      z_out_521, z_out_726, z_out_510, z_out_332, {(fsm_output[2]) , AccumDotWidth_or_153_cse
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_829_nl = MUX1HOT_v_22_8_2(z_out_370, z_out_329, z_out_261,
      z_out_520, z_out_717, z_out_235, z_out_521, AccumDotWidth_acc_1201_itm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_269 = (AccumDotWidth_mux1h_828_nl) + (AccumDotWidth_mux1h_829_nl);
  assign z_out_269 = nl_z_out_269[21:0];
  assign nl_AccumDotWidth_acc_2412_nl = z_out_560 + z_out_328;
  assign AccumDotWidth_acc_2412_nl = nl_AccumDotWidth_acc_2412_nl[21:0];
  assign AccumDotWidth_mux1h_830_nl = MUX1HOT_v_22_7_2(z_out_372, z_out_234, z_out_236,
      z_out_531, z_out_397, (AccumDotWidth_acc_2412_nl), z_out_511, {(fsm_output[2])
      , AccumDotWidth_or_153_cse , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_831_nl = MUX1HOT_v_22_8_2(z_out_369, z_out_320, z_out_260,
      z_out_523, z_out_723, z_out_322, z_out_524, AccumDotWidth_acc_1371_itm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_270 = (AccumDotWidth_mux1h_830_nl) + (AccumDotWidth_mux1h_831_nl);
  assign z_out_270 = nl_z_out_270[21:0];
  assign AccumDotWidth_or_156_cse = (fsm_output[3]) | (fsm_output[8]);
  assign nl_AccumDotWidth_acc_2413_nl = z_out_799 + z_out_797;
  assign AccumDotWidth_acc_2413_nl = nl_AccumDotWidth_acc_2413_nl[21:0];
  assign AccumDotWidth_mux1h_832_nl = MUX1HOT_v_22_8_2(z_out_389, z_out_564, z_out_531,
      z_out_710, z_out_686, z_out_256, (AccumDotWidth_acc_2413_nl), z_out_236, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_833_nl = MUX1HOT_v_22_7_2(z_out_393, z_out_531, AccumDotWidth_acc_1203_itm,
      z_out_711, z_out_688, z_out_341, z_out_528, {(fsm_output[2]) , (fsm_output[1])
      , AccumDotWidth_or_156_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_271 = (AccumDotWidth_mux1h_832_nl) + (AccumDotWidth_mux1h_833_nl);
  assign z_out_271 = nl_z_out_271[21:0];
  assign nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0))
      * $signed((w4_rsci_idat_mxwt[4063:4056]));
  assign MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign MultLoop_mux1h_374_nl = MUX1HOT_v_22_5_2(z_out_141_28_7, (readslicef_29_22_7((MultLoop_508_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      z_out_112_28_7, z_out_638_28_7, z_out_808, {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1374_nl = z_out_480 + MultLoop_acc_123_itm;
  assign MultLoop_acc_1374_nl = nl_MultLoop_acc_1374_nl[21:0];
  assign MultLoop_mux1h_375_nl = MUX1HOT_v_22_5_2(z_out_115_28_7, z_out_658_28_7,
      z_out_634_28_7, z_out_655_28_7, (MultLoop_acc_1374_nl), {(fsm_output[3]) ,
      (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_272 = (MultLoop_mux1h_374_nl) + (MultLoop_mux1h_375_nl);
  assign z_out_272 = nl_z_out_272[21:0];
  assign AccumDotWidth_or_157_cse = (fsm_output[3]) | (fsm_output[6]);
  assign AccumDotWidth_mux1h_834_nl = MUX1HOT_v_22_6_2(z_out_699, z_out_547, z_out_691,
      z_out_342, z_out_417, z_out_514, {(fsm_output[1]) , AccumDotWidth_or_157_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_835_nl = MUX1HOT_v_22_7_2(z_out_695, z_out_355, z_out_696,
      z_out_349, z_out_545, z_out_414, MultLoop_acc_587_itm, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_273 = (AccumDotWidth_mux1h_834_nl) + (AccumDotWidth_mux1h_835_nl);
  assign z_out_273 = nl_z_out_273[21:0];
  assign nl_MultLoop_acc_1376_nl = (z_out_615_29_7[21:0]) + MultLoop_739_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1376_nl = nl_MultLoop_acc_1376_nl[21:0];
  assign nl_MultLoop_acc_1375_nl = z_out_503 + (MultLoop_acc_1376_nl);
  assign MultLoop_acc_1375_nl = nl_MultLoop_acc_1375_nl[21:0];
  assign AccumDotWidth_mux1h_836_nl = MUX1HOT_v_22_8_2(z_out_691, AccumDotWidth_acc_1164_itm,
      z_out_556, z_out_719, z_out_340, z_out_805, z_out_703, (MultLoop_acc_1375_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1378_nl = MultLoop_740_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + (z_out_610_29_7[21:0]);
  assign MultLoop_acc_1378_nl = nl_MultLoop_acc_1378_nl[21:0];
  assign nl_MultLoop_acc_1377_nl = (MultLoop_acc_1378_nl) + z_out_500;
  assign MultLoop_acc_1377_nl = nl_MultLoop_acc_1377_nl[21:0];
  assign AccumDotWidth_mux1h_837_nl = MUX1HOT_v_22_8_2(z_out_694, z_out_429, z_out_353,
      z_out_720, z_out_341, z_out_336, z_out_706, (MultLoop_acc_1377_nl), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_274 = (AccumDotWidth_mux1h_836_nl) + (AccumDotWidth_mux1h_837_nl);
  assign z_out_274 = nl_z_out_274[21:0];
  assign nl_MultLoop_acc_1380_nl = (z_out_1127_29_7[21:0]) + MultLoop_321_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1380_nl = nl_MultLoop_acc_1380_nl[21:0];
  assign nl_MultLoop_acc_1379_nl = (MultLoop_acc_1380_nl) + z_out_316;
  assign MultLoop_acc_1379_nl = nl_MultLoop_acc_1379_nl[21:0];
  assign AccumDotWidth_mux1h_838_nl = MUX1HOT_v_22_7_2(z_out_352, z_out_696, z_out_235,
      z_out_704, z_out_528, z_out_705, (MultLoop_acc_1379_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_839_nl = MUX1HOT_v_22_6_2(z_out_365, z_out_698, AccumDotWidth_acc_1220_itm,
      z_out_705, z_out_529, AccumDotWidth_acc_1916_itm, {(fsm_output[2]) , (fsm_output[1])
      , AccumDotWidth_or_156_cse , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_275 = (AccumDotWidth_mux1h_838_nl) + (AccumDotWidth_mux1h_839_nl);
  assign z_out_275 = nl_z_out_275[21:0];
  assign MultLoop_mux1h_376_nl = MUX1HOT_v_22_7_2(z_out_52_28_7, z_out_646_28_7,
      z_out_190_28_7, z_out_92_28_7, z_out_59_28_7, z_out_91_28_7, z_out_44_28_7,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[7])});
  assign MultLoop_mux1h_377_nl = MUX1HOT_v_22_7_2(z_out_53_28_7, z_out_647_28_7,
      z_out_189_28_7, z_out_661_28_7, z_out_54_28_7, z_out_90_28_7, z_out_67_28_7,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[7])});
  assign nl_z_out_276 = (MultLoop_mux1h_376_nl) + (MultLoop_mux1h_377_nl);
  assign z_out_276 = nl_z_out_276[21:0];
  assign MultLoop_mux1h_378_nl = MUX1HOT_v_22_5_2(z_out_83_28_7, z_out_48_28_7, z_out_47_28_7,
      z_out_91_28_7, z_out_642_28_7, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_379_nl = MUX1HOT_v_22_5_2(z_out_169_28_7, z_out_116_28_7,
      z_out_45_28_7, z_out_96_28_7, z_out_641_28_7, {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_277 = (MultLoop_mux1h_378_nl) + (MultLoop_mux1h_379_nl);
  assign z_out_277 = nl_z_out_277[21:0];
  assign nl_MultLoop_acc_1381_nl = z_out_240 + z_out_229;
  assign MultLoop_acc_1381_nl = nl_MultLoop_acc_1381_nl[21:0];
  assign MultLoop_mux_84_nl = MUX_v_22_2_2(MultLoop_acc_1121_itm, (MultLoop_acc_1381_nl),
      fsm_output[8]);
  assign nl_z_out_278 = MultLoop_acc_628_itm + (MultLoop_mux_84_nl);
  assign z_out_278 = nl_z_out_278[21:0];
  assign MultLoop_mux1h_380_nl = MUX1HOT_v_22_6_2(z_out_123_28_7, z_out_50_28_7,
      z_out_108_28_7, z_out_38_28_7, z_out_94_28_7, z_out_49_28_7, {(fsm_output[5])
      , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2])});
  assign MultLoop_mux1h_381_nl = MUX1HOT_v_22_6_2(z_out_121_28_7, z_out_51_28_7,
      z_out_115_28_7, z_out_39_28_7, z_out_93_28_7, z_out_48_28_7, {(fsm_output[5])
      , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2])});
  assign nl_z_out_279 = (MultLoop_mux1h_380_nl) + (MultLoop_mux1h_381_nl);
  assign z_out_279 = nl_z_out_279[21:0];
  assign MultLoop_mux_85_nl = MUX_v_22_2_2(z_out_285, z_out_818, fsm_output[8]);
  assign nl_MultLoop_acc_1382_nl = MultLoop_acc_128_itm + z_out_509;
  assign MultLoop_acc_1382_nl = nl_MultLoop_acc_1382_nl[21:0];
  assign MultLoop_mux_86_nl = MUX_v_22_2_2(z_out_456, (MultLoop_acc_1382_nl), fsm_output[8]);
  assign nl_z_out_280 = (MultLoop_mux_85_nl) + (MultLoop_mux_86_nl);
  assign z_out_280 = nl_z_out_280[21:0];
  assign MultLoop_mux_87_nl = MUX_v_22_2_2(MultLoop_acc_1010_itm, z_out_837, fsm_output[8]);
  assign nl_z_out_281 = MultLoop_acc_243_itm + (MultLoop_mux_87_nl);
  assign z_out_281 = nl_z_out_281[21:0];
  assign MultLoop_mux1h_382_nl = MUX1HOT_v_22_4_2(z_out_113_28_7, z_out_637_28_7,
      z_out_96_28_7, z_out_49_28_7, {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5])});
  assign MultLoop_mux1h_383_nl = MUX1HOT_v_22_4_2(z_out_108_28_7, z_out_641_28_7,
      z_out_98_28_7, z_out_45_28_7, {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_z_out_282 = (MultLoop_mux1h_382_nl) + (MultLoop_mux1h_383_nl);
  assign z_out_282 = nl_z_out_282[21:0];
  assign MultLoop_mux1h_384_nl = MUX1HOT_v_22_6_2(MultLoop_acc_356_itm, z_out_690,
      z_out_551, z_out_412, z_out_546, z_out_416, {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_MultLoop_acc_1383_nl = z_out_799 + z_out_801;
  assign MultLoop_acc_1383_nl = nl_MultLoop_acc_1383_nl[21:0];
  assign MultLoop_mux1h_385_nl = MUX1HOT_v_22_7_2(MultLoop_acc_1018_itm, z_out_689,
      z_out_683, z_out_417, z_out_560, z_out_415, (MultLoop_acc_1383_nl), {(fsm_output[5])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_283 = (MultLoop_mux1h_384_nl) + (MultLoop_mux1h_385_nl);
  assign z_out_283 = nl_z_out_283[21:0];
  assign MultLoop_mux1h_386_nl = MUX1HOT_v_22_7_2(z_out_114_28_7, z_out_112_28_7,
      z_out_88_28_7, z_out_192_28_7, z_out_106_28_7, z_out_648_28_7, z_out_44_28_7,
      {(fsm_output[3]) , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[2])});
  assign MultLoop_mux1h_387_nl = MUX1HOT_v_22_7_2(z_out_49_28_7, z_out_111_28_7,
      z_out_184_28_7, z_out_191_28_7, z_out_44_28_7, z_out_99_28_7, z_out_43_28_7,
      {(fsm_output[3]) , (fsm_output[7]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[2])});
  assign nl_z_out_284 = (MultLoop_mux1h_386_nl) + (MultLoop_mux1h_387_nl);
  assign z_out_284 = nl_z_out_284[21:0];
  assign MultLoop_mux1h_388_nl = MUX1HOT_v_22_3_2(z_out_501, MultLoop_acc_689_itm,
      z_out_516, {(fsm_output[5]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse
      , (fsm_output[6])});
  assign MultLoop_mux1h_389_nl = MUX1HOT_v_22_4_2(z_out_502, z_out_845, z_out_524,
      z_out_843, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_285 = (MultLoop_mux1h_388_nl) + (MultLoop_mux1h_389_nl);
  assign z_out_285 = nl_z_out_285[21:0];
  assign nl_MultLoop_acc_1385_nl = (z_out_854_29_7[21:0]) + (z_out_853_29_7[21:0]);
  assign MultLoop_acc_1385_nl = nl_MultLoop_acc_1385_nl[21:0];
  assign nl_MultLoop_acc_1386_nl = (z_out_856_29_7[21:0]) + (z_out_860_29_7[21:0]);
  assign MultLoop_acc_1386_nl = nl_MultLoop_acc_1386_nl[21:0];
  assign nl_MultLoop_acc_1384_nl = (MultLoop_acc_1385_nl) + (MultLoop_acc_1386_nl);
  assign MultLoop_acc_1384_nl = nl_MultLoop_acc_1384_nl[21:0];
  assign MultLoop_mux_88_nl = MUX_v_22_2_2(MultLoop_acc_1089_itm, (MultLoop_acc_1384_nl),
      fsm_output[8]);
  assign nl_z_out_286 = MultLoop_acc_483_itm + (MultLoop_mux_88_nl);
  assign z_out_286 = nl_z_out_286[21:0];
  assign MultLoop_mux1h_390_nl = MUX1HOT_v_22_4_2(z_out_650_28_7, z_out_101_28_7,
      z_out_97_28_7, z_out_126_28_7, {(fsm_output[1]) , (fsm_output[4]) , AccumDotWidth_or_25_cse
      , (fsm_output[5])});
  assign MultLoop_mux1h_391_nl = MUX1HOT_v_22_5_2(z_out_651_28_7, z_out_110_28_7,
      z_out_96_28_7, z_out_98_28_7, z_out_130_28_7, {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_287 = (MultLoop_mux1h_390_nl) + (MultLoop_mux1h_391_nl);
  assign z_out_287 = nl_z_out_287[21:0];
  assign nl_MultLoop_acc_1387_nl = z_out_118_28_7 + z_out_119_28_7;
  assign MultLoop_acc_1387_nl = nl_MultLoop_acc_1387_nl[21:0];
  assign MultLoop_mux1h_392_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1387_nl), z_out_276,
      z_out_465, z_out_198, MultLoop_acc_243_itm, z_out_221, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1388_nl = z_out_120_28_7 + z_out_37_28_7;
  assign MultLoop_acc_1388_nl = nl_MultLoop_acc_1388_nl[21:0];
  assign MultLoop_mux1h_393_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1388_nl), z_out_282,
      z_out_279, z_out_194, MultLoop_acc_1121_itm, z_out_300, {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[8])});
  assign nl_z_out_288 = (MultLoop_mux1h_392_nl) + (MultLoop_mux1h_393_nl);
  assign z_out_288 = nl_z_out_288[21:0];
  assign MultLoop_or_87_cse = (fsm_output[5]) | (fsm_output[4]) | (fsm_output[2]);
  assign nl_MultLoop_acc_1389_nl = z_out_38_28_7 + z_out_39_28_7;
  assign MultLoop_acc_1389_nl = nl_MultLoop_acc_1389_nl[21:0];
  assign MultLoop_mux1h_394_nl = MUX1HOT_v_22_6_2((MultLoop_acc_1389_nl), MultLoop_acc_181_itm,
      z_out_840, z_out_300, z_out_276, z_out_436, {(fsm_output[1]) , MultLoop_or_87_cse
      , (fsm_output[6]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1390_nl = z_out_66_28_7 + MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1390_nl = nl_MultLoop_acc_1390_nl[21:0];
  assign MultLoop_mux1h_395_nl = MUX1HOT_v_22_7_2(z_out_436, z_out_284, z_out_829,
      MultLoop_acc_1018_itm, z_out_209, (MultLoop_acc_1390_nl), z_out_457, {MultLoop_or_81_cse
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_289 = (MultLoop_mux1h_394_nl) + (MultLoop_mux1h_395_nl);
  assign z_out_289 = nl_z_out_289[21:0];
  assign MultLoop_or_89_cse = (fsm_output[6]) | (fsm_output[2]);
  assign MultLoop_mux1h_396_nl = MUX1HOT_v_22_6_2(MultLoop_acc_128_itm, z_out_478,
      z_out_203, MultLoop_acc_435_itm, z_out_199, z_out_455, {MultLoop_or_89_cse
      , (fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1391_nl = MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_39_28_7;
  assign MultLoop_acc_1391_nl = nl_MultLoop_acc_1391_nl[21:0];
  assign nl_MultLoop_acc_1392_nl = z_out_55_28_7 + z_out_64_28_7;
  assign MultLoop_acc_1392_nl = nl_MultLoop_acc_1392_nl[21:0];
  assign MultLoop_mux1h_397_nl = MUX1HOT_v_22_8_2(MultLoop_acc_1121_itm, z_out_455,
      z_out_197, (MultLoop_acc_1391_nl), MultLoop_acc_1012_itm, z_out_452, (MultLoop_acc_1392_nl),
      z_out_195, {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_290 = (MultLoop_mux1h_396_nl) + (MultLoop_mux1h_397_nl);
  assign z_out_290 = nl_z_out_290[21:0];
  assign MultLoop_mux1h_398_nl = MUX1HOT_v_22_5_2(z_out_305, z_out_300, z_out_197,
      z_out_833, z_out_196, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3])});
  assign MultLoop_mux1h_399_nl = MUX1HOT_v_22_5_2(z_out_220, z_out_196, z_out_277,
      z_out_834, z_out_199, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3])});
  assign nl_z_out_291 = (MultLoop_mux1h_398_nl) + (MultLoop_mux1h_399_nl);
  assign z_out_291 = nl_z_out_291[21:0];
  assign nl_MultLoop_acc_1394_nl = MultLoop_acc_36_itm + z_out_838;
  assign MultLoop_acc_1394_nl = nl_MultLoop_acc_1394_nl[21:0];
  assign nl_MultLoop_acc_1393_nl = z_out_813 + (MultLoop_acc_1394_nl);
  assign MultLoop_acc_1393_nl = nl_MultLoop_acc_1393_nl[21:0];
  assign MultLoop_mux1h_400_nl = MUX1HOT_v_22_5_2(z_out_284, z_out_195, MultLoop_acc_308_itm,
      z_out_831, (MultLoop_acc_1393_nl), {MultLoop_or_22_cse , (fsm_output[1]) ,
      MultLoop_or_87_cse , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1395_nl = z_out_35_28_7 + z_out_68_28_7;
  assign MultLoop_acc_1395_nl = nl_MultLoop_acc_1395_nl[21:0];
  assign MultLoop_mux1h_401_nl = MUX1HOT_v_22_8_2(z_out_279, z_out_210, z_out_201,
      z_out_443, z_out_830, MultLoop_acc_113_itm, (MultLoop_acc_1395_nl), z_out_209,
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[7]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_292 = (MultLoop_mux1h_400_nl) + (MultLoop_mux1h_401_nl);
  assign z_out_292 = nl_z_out_292[21:0];
  assign MultLoop_or_93_cse = (fsm_output[2]) | (fsm_output[5]);
  assign MultLoop_mux1h_402_nl = MUX1HOT_v_22_4_2(z_out_199, z_out_276, z_out_846,
      z_out_201, {(fsm_output[1]) , (fsm_output[4]) , MultLoop_or_93_cse , (fsm_output[3])});
  assign MultLoop_mux1h_403_nl = MUX1HOT_v_22_4_2(z_out_196, z_out_198, z_out_828,
      z_out_197, {(fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[2]) , (fsm_output[5])});
  assign nl_z_out_293 = (MultLoop_mux1h_402_nl) + (MultLoop_mux1h_403_nl);
  assign z_out_293 = nl_z_out_293[21:0];
  assign nl_MultLoop_acc_1396_nl = z_out_45_28_7 + z_out_48_28_7;
  assign MultLoop_acc_1396_nl = nl_MultLoop_acc_1396_nl[21:0];
  assign MultLoop_mux1h_404_nl = MUX1HOT_v_22_4_2((MultLoop_acc_1396_nl), z_out_209,
      z_out_277, z_out_306, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[3])});
  assign MultLoop_mux1h_405_nl = MUX1HOT_v_22_4_2(z_out_443, z_out_284, z_out_287,
      z_out_301, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_z_out_294 = (MultLoop_mux1h_404_nl) + (MultLoop_mux1h_405_nl);
  assign z_out_294 = nl_z_out_294[21:0];
  assign MultLoop_mux1h_406_nl = MUX1HOT_v_22_4_2(z_out_284, z_out_220, z_out_282,
      z_out_305, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign MultLoop_mux1h_407_nl = MUX1HOT_v_22_4_2(z_out_300, z_out_282, z_out_306,
      z_out_268, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_z_out_295 = (MultLoop_mux1h_406_nl) + (MultLoop_mux1h_407_nl);
  assign z_out_295 = nl_z_out_295[21:0];
  assign MultLoop_mux1h_408_nl = MUX1HOT_v_22_3_2(z_out_272, z_out_485, z_out_208,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_mux1h_409_nl = MUX1HOT_v_22_3_2(z_out_202, z_out_479, z_out_205,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_296 = (MultLoop_mux1h_408_nl) + (MultLoop_mux1h_409_nl);
  assign z_out_296 = nl_z_out_296[21:0];
  assign MultLoop_mux1h_410_nl = MUX1HOT_v_22_3_2(z_out_209, z_out_831, z_out_202,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign MultLoop_mux1h_411_nl = MUX1HOT_v_22_3_2(z_out_221, z_out_300, z_out_205,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_z_out_297 = (MultLoop_mux1h_410_nl) + (MultLoop_mux1h_411_nl);
  assign z_out_297 = nl_z_out_297[21:0];
  assign nl_MultLoop_acc_1397_nl = z_out_105_28_7 + z_out_645_28_7;
  assign MultLoop_acc_1397_nl = nl_MultLoop_acc_1397_nl[21:0];
  assign nl_MultLoop_acc_1398_nl = z_out_822 + z_out_444;
  assign MultLoop_acc_1398_nl = nl_MultLoop_acc_1398_nl[21:0];
  assign MultLoop_mux1h_412_nl = MUX1HOT_v_22_6_2(z_out_824, z_out_272, z_out_831,
      MultLoop_acc_54_itm, (MultLoop_acc_1397_nl), (MultLoop_acc_1398_nl), {(fsm_output[6])
      , (fsm_output[3]) , (fsm_output[2]) , AccumDotWidth_or_38_cse , (fsm_output[1])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1399_nl = z_out_106_28_7 + z_out_103_28_7;
  assign MultLoop_acc_1399_nl = nl_MultLoop_acc_1399_nl[21:0];
  assign nl_MultLoop_acc_1400_nl = MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_100_28_7;
  assign MultLoop_acc_1400_nl = nl_MultLoop_acc_1400_nl[21:0];
  assign nl_MultLoop_acc_1401_nl = z_out_93_28_7 + z_out_83_28_7;
  assign MultLoop_acc_1401_nl = nl_MultLoop_acc_1401_nl[21:0];
  assign MultLoop_mux1h_413_nl = MUX1HOT_v_22_7_2(z_out_832, (MultLoop_acc_1399_nl),
      MultLoop_acc_1095_itm, (MultLoop_acc_1400_nl), z_out_276, (MultLoop_acc_1401_nl),
      z_out_204, {(fsm_output[6]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_298 = (MultLoop_mux1h_412_nl) + (MultLoop_mux1h_413_nl);
  assign z_out_298 = nl_z_out_298[21:0];
  assign MultLoop_mux1h_414_nl = MUX1HOT_v_22_3_2(z_out_301, z_out_207, z_out_203,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign MultLoop_mux1h_415_nl = MUX1HOT_v_22_3_2(z_out_233, z_out_202, z_out_207,
      {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])});
  assign nl_z_out_299 = (MultLoop_mux1h_414_nl) + (MultLoop_mux1h_415_nl);
  assign z_out_299 = nl_z_out_299[21:0];
  assign nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1932_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9919:9912]));
  assign MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1937_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9927:9920]));
  assign MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1413_nl = (readslicef_29_22_7((MultLoop_1240_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1241_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1413_nl = nl_MultLoop_acc_1413_nl[21:0];
  assign nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1945_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9935:9928]));
  assign MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0]))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9943:9936]));
  assign MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1414_nl = (readslicef_29_22_7((MultLoop_1242_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1243_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1414_nl = nl_MultLoop_acc_1414_nl[21:0];
  assign nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9855:9848]));
  assign MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1406_nl = (readslicef_29_22_7((MultLoop_1232_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (z_out_621_29_7[21:0]);
  assign MultLoop_acc_1406_nl = nl_MultLoop_acc_1406_nl[21:0];
  assign nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9871:9864]));
  assign MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9879:9872]));
  assign MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1407_nl = (readslicef_29_22_7((MultLoop_1234_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1235_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1407_nl = nl_MultLoop_acc_1407_nl[21:0];
  assign nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9887:9880]));
  assign MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1871_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9895:9888]));
  assign MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1409_nl = (readslicef_29_22_7((MultLoop_1236_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1237_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1409_nl = nl_MultLoop_acc_1409_nl[21:0];
  assign nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1877_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9903:9896]));
  assign MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1916_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[9911:9904]));
  assign MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1410_nl = (readslicef_29_22_7((MultLoop_1238_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1239_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1410_nl = nl_MultLoop_acc_1410_nl[21:0];
  assign nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0]))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9951:9944]));
  assign MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9959:9952]));
  assign MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1416_nl = (readslicef_29_22_7((MultLoop_1244_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1245_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1416_nl = nl_MultLoop_acc_1416_nl[21:0];
  assign nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9967:9960]));
  assign MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9975:9968]));
  assign MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1417_nl = (readslicef_29_22_7((MultLoop_1246_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1247_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1417_nl = nl_MultLoop_acc_1417_nl[21:0];
  assign nl_MultLoop_acc_1403_nl = (MultLoop_acc_1413_nl) + (MultLoop_acc_1414_nl)
      + (MultLoop_acc_1406_nl) + (MultLoop_acc_1407_nl) + (MultLoop_acc_1409_nl)
      + (MultLoop_acc_1410_nl) + (MultLoop_acc_1416_nl) + (MultLoop_acc_1417_nl);
  assign MultLoop_acc_1403_nl = nl_MultLoop_acc_1403_nl[21:0];
  assign nl_MultLoop_acc_1402_nl = z_out_541 + (MultLoop_acc_1403_nl);
  assign MultLoop_acc_1402_nl = nl_MultLoop_acc_1402_nl[21:0];
  assign MultLoop_mux1h_416_nl = MUX1HOT_v_22_5_2(z_out_154_28_7, z_out_67_28_7,
      z_out_139_28_7, z_out_41_28_7, (MultLoop_acc_1402_nl), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign MultLoop_mux1h_417_nl = MUX1HOT_v_22_5_2(z_out_95_28_7, z_out_91_28_7, z_out_654_28_7,
      z_out_99_28_7, z_out_763, {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_300 = (MultLoop_mux1h_416_nl) + (MultLoop_mux1h_417_nl);
  assign z_out_300 = nl_z_out_300[21:0];
  assign MultLoop_mux1h_418_nl = MUX1HOT_v_22_4_2(z_out_49_28_7, z_out_635_28_7,
      z_out_93_28_7, z_out_137_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5])});
  assign MultLoop_mux1h_419_nl = MUX1HOT_v_22_4_2(z_out_95_28_7, z_out_649_28_7,
      z_out_90_28_7, z_out_119_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5])});
  assign nl_z_out_301 = (MultLoop_mux1h_418_nl) + (MultLoop_mux1h_419_nl);
  assign z_out_301 = nl_z_out_301[21:0];
  assign MultLoop_mux1h_420_nl = MUX1HOT_v_22_3_2(z_out_306, z_out_208, z_out_203,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_mux1h_421_nl = MUX1HOT_v_22_3_2(z_out_208, z_out_198, z_out_210,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_302 = (MultLoop_mux1h_420_nl) + (MultLoop_mux1h_421_nl);
  assign z_out_302 = nl_z_out_302[21:0];
  assign MultLoop_mux1h_422_nl = MUX1HOT_v_22_6_2(MultLoop_acc_562_itm, z_out_833,
      z_out_824, z_out_287, z_out_277, z_out_280, {AccumDotWidth_or_38_cse , (fsm_output[6])
      , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1418_nl = MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_122_28_7;
  assign MultLoop_acc_1418_nl = nl_MultLoop_acc_1418_nl[21:0];
  assign nl_MultLoop_acc_1419_nl = z_out_636_28_7 + z_out_77_28_7;
  assign MultLoop_acc_1419_nl = nl_MultLoop_acc_1419_nl[21:0];
  assign MultLoop_mux1h_423_nl = MUX1HOT_v_22_7_2((MultLoop_acc_1418_nl), z_out_834,
      (MultLoop_acc_1419_nl), z_out_832, z_out_204, z_out_287, z_out_272, {(fsm_output[5])
      , (fsm_output[6]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[8])});
  assign nl_z_out_303 = (MultLoop_mux1h_422_nl) + (MultLoop_mux1h_423_nl);
  assign z_out_303 = nl_z_out_303[21:0];
  assign MultLoop_mux1h_424_nl = MUX1HOT_v_22_3_2(z_out_305, z_out_457, z_out_276,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_mux1h_425_nl = MUX1HOT_v_22_3_2(z_out_203, z_out_268, z_out_221,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_304 = (MultLoop_mux1h_424_nl) + (MultLoop_mux1h_425_nl);
  assign z_out_304 = nl_z_out_304[21:0];
  assign MultLoop_mux1h_426_nl = MUX1HOT_v_22_4_2(z_out_105_28_7, z_out_94_28_7,
      z_out_661_28_7, z_out_109_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[3])});
  assign MultLoop_mux1h_427_nl = MUX1HOT_v_22_4_2(z_out_660_28_7, z_out_93_28_7,
      z_out_656_28_7, z_out_110_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[1])
      , (fsm_output[3])});
  assign nl_z_out_305 = (MultLoop_mux1h_426_nl) + (MultLoop_mux1h_427_nl);
  assign z_out_305 = nl_z_out_305[21:0];
  assign MultLoop_mux1h_428_nl = MUX1HOT_v_22_3_2(z_out_106_28_7, z_out_40_28_7,
      z_out_177_28_7, {AccumDotWidth_or_132_cse_1 , (fsm_output[5]) , (fsm_output[3])});
  assign MultLoop_mux1h_429_nl = MUX1HOT_v_22_4_2(z_out_90_28_7, z_out_663_28_7,
      z_out_43_28_7, z_out_92_28_7, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[3])});
  assign nl_z_out_306 = (MultLoop_mux1h_428_nl) + (MultLoop_mux1h_429_nl);
  assign z_out_306 = nl_z_out_306[21:0];
  assign AccumDotWidth_mux1h_840_nl = MUX1HOT_v_22_7_2(z_out_742, z_out_720, z_out_721,
      z_out_683, z_out_802, z_out_707, (z_out_1100_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_841_nl = MUX1HOT_v_22_7_2(z_out_697, z_out_721, z_out_715,
      z_out_345, z_out_807, z_out_711, (z_out_1097_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_307 = (AccumDotWidth_mux1h_840_nl) + (AccumDotWidth_mux1h_841_nl);
  assign z_out_307 = nl_z_out_307[21:0];
  assign AccumDotWidth_mux1h_842_nl = MUX1HOT_v_22_6_2(z_out_363, z_out_697, z_out_692,
      z_out_377, z_out_701, (z_out_584_29_7[21:0]), {(fsm_output[1]) , MultLoop_or_46_cse
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_843_nl = MUX1HOT_v_22_6_2(z_out_357, z_out_698, z_out_697,
      z_out_387, z_out_700, (z_out_585_29_7[21:0]), {(fsm_output[1]) , MultLoop_or_46_cse
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_308 = (AccumDotWidth_mux1h_842_nl) + (AccumDotWidth_mux1h_843_nl);
  assign z_out_308 = nl_z_out_308[21:0];
  assign AccumDotWidth_mux1h_844_nl = MUX1HOT_v_22_4_2(AccumDotWidth_acc_1300_itm,
      AccumDotWidth_acc_1392_itm, z_out_429, (z_out_985_29_7[21:0]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2415_nl = (nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2415_nl = nl_AccumDotWidth_acc_2415_nl[9:0];
  assign nl_AccumDotWidth_acc_2414_nl = AccumDotWidth_acc_1378_itm + conv_s2s_21_22({(AccumDotWidth_acc_2415_nl)
      , (nnet_relu_layer2_t_layer3_t_relu_config3_for_11_if_exu_pmx_20_0_lpi_1_dfm[10:0])});
  assign AccumDotWidth_acc_2414_nl = nl_AccumDotWidth_acc_2414_nl[21:0];
  assign AccumDotWidth_mux1h_845_nl = MUX1HOT_v_22_4_2(z_out_427, (AccumDotWidth_acc_2414_nl),
      AccumDotWidth_acc_1203_itm, (z_out_984_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_309 = (AccumDotWidth_mux1h_844_nl) + (AccumDotWidth_mux1h_845_nl);
  assign z_out_309 = nl_z_out_309[21:0];
  assign nl_AccumDotWidth_acc_2416_nl = conv_s2s_21_22(z_out_1099_29_7[22:2]) + conv_s2s_21_22(z_out_1182_29_7[22:2]);
  assign AccumDotWidth_acc_2416_nl = nl_AccumDotWidth_acc_2416_nl[21:0];
  assign AccumDotWidth_mux1h_846_nl = MUX1HOT_v_22_6_2(z_out_720, z_out_694, (AccumDotWidth_acc_2416_nl),
      z_out_731, z_out_352, (z_out_588_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2417_nl = conv_s2s_21_22(z_out_1064_29_7[22:2]) + conv_s2s_21_22(z_out_1070_29_7[22:2]);
  assign AccumDotWidth_acc_2417_nl = nl_AccumDotWidth_acc_2417_nl[21:0];
  assign AccumDotWidth_mux1h_847_nl = MUX1HOT_v_22_6_2(z_out_721, z_out_691, (AccumDotWidth_acc_2417_nl),
      z_out_733, z_out_366, (z_out_589_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_310 = (AccumDotWidth_mux1h_846_nl) + (AccumDotWidth_mux1h_847_nl);
  assign z_out_310 = nl_z_out_310[21:0];
  assign nl_AccumDotWidth_acc_2418_nl = conv_s2s_21_22(z_out_859_29_7[22:2]) + conv_s2s_21_22(z_out_903_29_7[22:2]);
  assign AccumDotWidth_acc_2418_nl = nl_AccumDotWidth_acc_2418_nl[21:0];
  assign AccumDotWidth_mux1h_848_nl = MUX1HOT_v_22_4_2(z_out_692, z_out_695, (AccumDotWidth_acc_2418_nl),
      (z_out_954_29_7[21:0]), {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2419_nl = conv_s2s_21_22(z_out_1141_29_9) + conv_s2s_21_22(z_out_976_29_7[22:2]);
  assign AccumDotWidth_acc_2419_nl = nl_AccumDotWidth_acc_2419_nl[21:0];
  assign AccumDotWidth_mux1h_849_nl = MUX1HOT_v_22_4_2(z_out_693, z_out_696, (AccumDotWidth_acc_2419_nl),
      (z_out_955_29_7[21:0]), {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_311 = (AccumDotWidth_mux1h_848_nl) + (AccumDotWidth_mux1h_849_nl);
  assign z_out_311 = nl_z_out_311[21:0];
  assign AccumDotWidth_mux_92_nl = MUX_v_22_2_2(z_out_361, (z_out_881_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_93_nl = MUX_v_22_2_2(z_out_364, (z_out_580_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_312 = (AccumDotWidth_mux_92_nl) + (AccumDotWidth_mux_93_nl);
  assign z_out_312 = nl_z_out_312[21:0];
  assign AccumDotWidth_mux1h_850_nl = MUX1HOT_v_22_4_2(z_out_364, z_out_413, z_out_724,
      (z_out_604_29_7[21:0]), {(fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse
      , (fsm_output[5]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_851_nl = MUX1HOT_v_22_5_2(z_out_363, z_out_414, z_out_716,
      z_out_412, (z_out_606_29_7[21:0]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_313 = (AccumDotWidth_mux1h_850_nl) + (AccumDotWidth_mux1h_851_nl);
  assign z_out_313 = nl_z_out_313[21:0];
  assign nl_AccumDotWidth_acc_2420_nl = conv_s2s_21_22(z_out_914_29_7[22:2]) + conv_s2s_21_22(z_out_856_29_7[22:2]);
  assign AccumDotWidth_acc_2420_nl = nl_AccumDotWidth_acc_2420_nl[21:0];
  assign AccumDotWidth_mux1h_852_nl = MUX1HOT_v_22_5_2(z_out_358, z_out_695, (AccumDotWidth_acc_2420_nl),
      z_out_738, (z_out_1098_29_7[21:0]), {AccumDotWidth_or_149_cse , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2421_nl = conv_s2s_21_22(z_out_994_29_7[22:2]) + conv_s2s_21_22(z_out_906_29_7[22:2]);
  assign AccumDotWidth_acc_2421_nl = nl_AccumDotWidth_acc_2421_nl[21:0];
  assign AccumDotWidth_mux1h_853_nl = MUX1HOT_v_22_5_2(z_out_350, z_out_696, (AccumDotWidth_acc_2421_nl),
      z_out_684, (z_out_1106_29_7[21:0]), {AccumDotWidth_or_149_cse , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_314 = (AccumDotWidth_mux1h_852_nl) + (AccumDotWidth_mux1h_853_nl);
  assign z_out_314 = nl_z_out_314[21:0];
  assign nl_AccumDotWidth_acc_2422_nl = conv_s2s_21_22(z_out_1005_29_7[22:2]) + conv_s2s_21_22(z_out_1047_29_9);
  assign AccumDotWidth_acc_2422_nl = nl_AccumDotWidth_acc_2422_nl[21:0];
  assign AccumDotWidth_mux1h_854_nl = MUX1HOT_v_22_6_2(z_out_356, z_out_722, z_out_706,
      z_out_681, (AccumDotWidth_acc_2422_nl), (z_out_908_29_7[21:0]), {AccumDotWidth_or_149_cse
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2423_nl = conv_s2s_21_22(z_out_1120_29_7[22:2]) + conv_s2s_21_22(z_out_589_29_7[22:2]);
  assign AccumDotWidth_acc_2423_nl = nl_AccumDotWidth_acc_2423_nl[21:0];
  assign AccumDotWidth_mux1h_855_nl = MUX1HOT_v_22_6_2(z_out_360, z_out_359, z_out_707,
      z_out_680, (AccumDotWidth_acc_2423_nl), (z_out_956_29_7[21:0]), {AccumDotWidth_or_149_cse
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_315 = (AccumDotWidth_mux1h_854_nl) + (AccumDotWidth_mux1h_855_nl);
  assign z_out_315 = nl_z_out_315[21:0];
  assign AccumDotWidth_mux1h_856_nl = MUX1HOT_v_22_7_2(z_out_364, z_out_365, z_out_699,
      z_out_691, z_out_378, z_out_710, (z_out_1124_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_857_nl = MUX1HOT_v_22_6_2(z_out_361, z_out_690, z_out_692,
      z_out_383, z_out_704, (z_out_1120_29_7[21:0]), {(fsm_output[1]) , AccumDotWidth_or_139_cse
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_316 = (AccumDotWidth_mux1h_856_nl) + (AccumDotWidth_mux1h_857_nl);
  assign z_out_316 = nl_z_out_316[21:0];
  assign AccumDotWidth_mux1h_858_nl = MUX1HOT_v_22_7_2(z_out_416, z_out_262, z_out_252,
      z_out_332, z_out_683, z_out_256, z_out_260, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1420_nl = (z_out_927_29_7[21:0]) + (z_out_928_29_7[21:0]);
  assign MultLoop_acc_1420_nl = nl_MultLoop_acc_1420_nl[21:0];
  assign AccumDotWidth_mux1h_859_nl = MUX1HOT_v_22_7_2(z_out_417, z_out_316, z_out_552,
      z_out_333, z_out_688, z_out_793, (MultLoop_acc_1420_nl), {(fsm_output[2]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_317 = (AccumDotWidth_mux1h_858_nl) + (AccumDotWidth_mux1h_859_nl);
  assign z_out_317 = nl_z_out_317[21:0];
  assign AccumDotWidth_mux1h_860_nl = MUX1HOT_v_22_7_2(z_out_418, z_out_255, z_out_254,
      z_out_259, z_out_273, z_out_262, z_out_795, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_861_nl = MUX1HOT_v_22_7_2(z_out_419, z_out_552, z_out_316,
      z_out_252, z_out_283, z_out_273, z_out_261, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_318 = (AccumDotWidth_mux1h_860_nl) + (AccumDotWidth_mux1h_861_nl);
  assign z_out_318 = nl_z_out_318[21:0];
  assign AccumDotWidth_mux1h_862_nl = MUX1HOT_v_22_7_2(z_out_307, z_out_342, z_out_250,
      z_out_524, z_out_686, z_out_252, z_out_804, {(fsm_output[1]) , (fsm_output[2])
      , MultLoop_or_46_cse , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_863_nl = MUX1HOT_v_22_8_2(z_out_273, z_out_398, z_out_310,
      z_out_553, z_out_527, z_out_687, z_out_274, z_out_259, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_319 = (AccumDotWidth_mux1h_862_nl) + (AccumDotWidth_mux1h_863_nl);
  assign z_out_319 = nl_z_out_319[21:0];
  assign AccumDotWidth_mux1h_864_nl = MUX1HOT_v_22_8_2(z_out_414, z_out_349, z_out_394,
      z_out_802, z_out_549, z_out_684, z_out_567, z_out_313, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1421_nl = (z_out_601_29_7[21:0]) + (z_out_602_29_7[21:0]);
  assign MultLoop_acc_1421_nl = nl_MultLoop_acc_1421_nl[21:0];
  assign AccumDotWidth_mux1h_865_nl = MUX1HOT_v_22_8_2(z_out_415, z_out_726, z_out_392,
      z_out_807, z_out_551, z_out_689, z_out_346, (MultLoop_acc_1421_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_320 = (AccumDotWidth_mux1h_864_nl) + (AccumDotWidth_mux1h_865_nl);
  assign z_out_320 = nl_z_out_320[21:0];
  assign AccumDotWidth_mux1h_866_nl = MUX1HOT_v_22_6_2(z_out_794, z_out_686, z_out_546,
      z_out_371, z_out_684, z_out_805, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1422_nl = (z_out_1085_29_7[21:0]) + (z_out_1084_29_7[21:0]);
  assign MultLoop_acc_1422_nl = nl_MultLoop_acc_1422_nl[21:0];
  assign AccumDotWidth_mux1h_867_nl = MUX1HOT_v_22_6_2(z_out_688, z_out_355, z_out_338,
      z_out_372, z_out_387, (MultLoop_acc_1422_nl), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_321 = (AccumDotWidth_mux1h_866_nl) + (AccumDotWidth_mux1h_867_nl);
  assign z_out_321 = nl_z_out_321[21:0];
  assign nl_MultLoop_acc_1423_nl = (z_out_1088_29_7[21:0]) + (z_out_1087_29_7[21:0]);
  assign MultLoop_acc_1423_nl = nl_MultLoop_acc_1423_nl[21:0];
  assign AccumDotWidth_mux1h_868_nl = MUX1HOT_v_22_3_2(z_out_848, z_out_373, (MultLoop_acc_1423_nl),
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_869_nl = MUX1HOT_v_22_3_2(z_out_328, z_out_374, z_out_797,
      {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_322 = (AccumDotWidth_mux1h_868_nl) + (AccumDotWidth_mux1h_869_nl);
  assign z_out_322 = nl_z_out_322[21:0];
  assign AccumDotWidth_mux1h_870_nl = MUX1HOT_v_22_7_2(z_out_686, z_out_369, z_out_260,
      z_out_558, AccumDotWidth_acc_1426_itm, z_out_556, z_out_793, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_871_nl = MUX1HOT_v_22_7_2(z_out_727, z_out_372, z_out_313,
      z_out_547, z_out_307, z_out_336, z_out_778, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_323 = (AccumDotWidth_mux1h_870_nl) + (AccumDotWidth_mux1h_871_nl);
  assign z_out_323 = nl_z_out_323[21:0];
  assign AccumDotWidth_mux_94_nl = MUX_v_22_2_2(z_out_807, z_out_780, fsm_output[8]);
  assign AccumDotWidth_mux_95_nl = MUX_v_22_2_2(z_out_802, z_out_791, fsm_output[8]);
  assign nl_z_out_324 = (AccumDotWidth_mux_94_nl) + (AccumDotWidth_mux_95_nl);
  assign z_out_324 = nl_z_out_324[21:0];
  assign AccumDotWidth_mux1h_872_nl = MUX1HOT_v_22_6_2(z_out_256, z_out_274, z_out_266,
      z_out_259, z_out_255, z_out_248, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1424_nl = (z_out_598_29_7[21:0]) + (z_out_593_29_7[21:0]);
  assign MultLoop_acc_1424_nl = nl_MultLoop_acc_1424_nl[21:0];
  assign AccumDotWidth_mux1h_873_nl = MUX1HOT_v_22_6_2(z_out_826, AccumDotWidth_acc_1133_itm,
      z_out_307, z_out_283, z_out_313, (MultLoop_acc_1424_nl), {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_325 = (AccumDotWidth_mux1h_872_nl) + (AccumDotWidth_mux1h_873_nl);
  assign z_out_325 = nl_z_out_325[21:0];
  assign nl_MultLoop_acc_1425_nl = (z_out_1010_29_7[21:0]) + (z_out_1015_29_7[21:0]);
  assign MultLoop_acc_1425_nl = nl_MultLoop_acc_1425_nl[21:0];
  assign AccumDotWidth_mux1h_874_nl = MUX1HOT_v_22_4_2(z_out_274, z_out_799, z_out_680,
      (MultLoop_acc_1425_nl), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1426_nl = (z_out_605_29_7[21:0]) + (z_out_608_29_7[21:0]);
  assign MultLoop_acc_1426_nl = nl_MultLoop_acc_1426_nl[21:0];
  assign AccumDotWidth_mux1h_875_nl = MUX1HOT_v_22_4_2(z_out_799, z_out_794, z_out_682,
      (MultLoop_acc_1426_nl), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_326 = (AccumDotWidth_mux1h_874_nl) + (AccumDotWidth_mux1h_875_nl);
  assign z_out_326 = nl_z_out_326[21:0];
  assign nl_MultLoop_acc_1427_nl = (z_out_603_29_7[21:0]) + (z_out_1121_29_7[21:0]);
  assign MultLoop_acc_1427_nl = nl_MultLoop_acc_1427_nl[21:0];
  assign AccumDotWidth_mux1h_876_nl = MUX1HOT_v_22_4_2(z_out_532, z_out_430, z_out_686,
      (MultLoop_acc_1427_nl), {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1428_nl = (z_out_1122_29_7[21:0]) + (z_out_1126_29_7[21:0]);
  assign MultLoop_acc_1428_nl = nl_MultLoop_acc_1428_nl[21:0];
  assign AccumDotWidth_mux1h_877_nl = MUX1HOT_v_22_4_2(z_out_556, z_out_431, z_out_386,
      (MultLoop_acc_1428_nl), {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_327 = (AccumDotWidth_mux1h_876_nl) + (AccumDotWidth_mux1h_877_nl);
  assign z_out_327 = nl_z_out_327[21:0];
  assign nl_MultLoop_acc_1429_nl = (z_out_953_29_7[21:0]) + (z_out_1125_29_7[21:0]);
  assign MultLoop_acc_1429_nl = nl_MultLoop_acc_1429_nl[21:0];
  assign AccumDotWidth_mux1h_878_nl = MUX1HOT_v_22_5_2(AccumDotWidth_acc_1326_itm,
      z_out_725, z_out_748, z_out_690, (MultLoop_acc_1429_nl), {(fsm_output[3]) ,
      AccumDotWidth_or_38_cse , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2424_nl = (z_out_907_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2424_nl = nl_AccumDotWidth_acc_2424_nl[9:0];
  assign nl_AccumDotWidth_acc_2425_nl = (z_out_992_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2425_nl = nl_AccumDotWidth_acc_2425_nl[9:0];
  assign nl_AccumDotWidth_acc_2426_nl = (z_out_582_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2426_nl = nl_AccumDotWidth_acc_2426_nl[9:0];
  assign nl_AccumDotWidth_acc_2427_nl = (z_out_885_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2427_nl = nl_AccumDotWidth_acc_2427_nl[9:0];
  assign AccumDotWidth_mux1h_879_nl = MUX1HOT_v_11_6_2(({{1{z_out_31[9]}}, z_out_31}),
      (signext_11_10(AccumDotWidth_acc_2424_nl)), (signext_11_10(AccumDotWidth_acc_2425_nl)),
      (signext_11_10(AccumDotWidth_acc_2426_nl)), (signext_11_10(AccumDotWidth_acc_2427_nl)),
      (MultLoop_acc_162_sdt[21:11]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_880_nl = MUX1HOT_v_11_6_2((nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm[10:0]),
      (z_out_907_29_7[12:2]), (z_out_992_29_9[10:0]), (z_out_582_29_7[12:2]), (z_out_885_29_7[12:2]),
      (MultLoop_acc_162_sdt[10:0]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_328 = (AccumDotWidth_mux1h_878_nl) + ({(AccumDotWidth_mux1h_879_nl)
      , (AccumDotWidth_mux1h_880_nl)});
  assign z_out_328 = nl_z_out_328[21:0];
  assign nl_AccumDotWidth_acc_2428_nl = conv_s2s_21_22(z_out_880_29_7[22:2]) + conv_s2s_21_22(z_out_610_29_7[22:2]);
  assign AccumDotWidth_acc_2428_nl = nl_AccumDotWidth_acc_2428_nl[21:0];
  assign nl_MultLoop_acc_1430_nl = (z_out_919_29_7[21:0]) + MultLoop_961_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1430_nl = nl_MultLoop_acc_1430_nl[21:0];
  assign AccumDotWidth_mux1h_881_nl = MUX1HOT_v_22_6_2(z_out_354, (AccumDotWidth_acc_2428_nl),
      z_out_395, z_out_734, z_out_379, (MultLoop_acc_1430_nl), {AccumDotWidth_or_153_cse
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2429_nl = conv_s2s_21_22(z_out_1037_29_7[22:2]) + conv_s2s_21_22(z_out_1074_29_7[22:2]);
  assign AccumDotWidth_acc_2429_nl = nl_AccumDotWidth_acc_2429_nl[21:0];
  assign nl_AccumDotWidth_acc_2430_nl = (z_out_900_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2430_nl = nl_AccumDotWidth_acc_2430_nl[9:0];
  assign nl_MultLoop_acc_1431_nl = (z_out_1184_29_7[21:0]) + (z_out_1173_29_7[21:0]);
  assign MultLoop_acc_1431_nl = nl_MultLoop_acc_1431_nl[21:0];
  assign AccumDotWidth_mux1h_882_nl = MUX1HOT_v_22_7_2(z_out_729, (AccumDotWidth_acc_2429_nl),
      z_out_396, z_out_400, (signext_22_21({(AccumDotWidth_acc_2430_nl) , (z_out_900_29_7[12:2])})),
      z_out_397, (MultLoop_acc_1431_nl), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_329 = (AccumDotWidth_mux1h_881_nl) + (AccumDotWidth_mux1h_882_nl);
  assign z_out_329 = nl_z_out_329[21:0];
  assign AccumDotWidth_mux1h_883_nl = MUX1HOT_v_22_5_2(z_out_273, z_out_806, z_out_393,
      z_out_807, z_out_554, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_46_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[367:360]));
  assign MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_47_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[375:368]));
  assign MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1432_nl = (readslicef_29_22_7((MultLoop_46_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_47_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1432_nl = nl_MultLoop_acc_1432_nl[21:0];
  assign AccumDotWidth_mux1h_884_nl = MUX1HOT_v_22_5_2(z_out_826, z_out_795, z_out_394,
      z_out_802, (MultLoop_acc_1432_nl), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_330 = (AccumDotWidth_mux1h_883_nl) + (AccumDotWidth_mux1h_884_nl);
  assign z_out_330 = nl_z_out_330[21:0];
  assign nl_AccumDotWidth_acc_2431_nl = conv_s2s_21_22(z_out_935_29_7[22:2]) + conv_s2s_21_22(z_out_609_29_7[22:2]);
  assign AccumDotWidth_acc_2431_nl = nl_AccumDotWidth_acc_2431_nl[21:0];
  assign nl_MultLoop_acc_1433_nl = (z_out_921_29_7[21:0]) + (z_out_920_29_7[21:0]);
  assign MultLoop_acc_1433_nl = nl_MultLoop_acc_1433_nl[21:0];
  assign AccumDotWidth_mux1h_885_nl = MUX1HOT_v_22_6_2(AccumDotWidth_acc_1274_itm,
      z_out_394, z_out_400, z_out_363, (AccumDotWidth_acc_2431_nl), (MultLoop_acc_1433_nl),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2432_nl = (z_out_901_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2432_nl = nl_AccumDotWidth_acc_2432_nl[9:0];
  assign nl_AccumDotWidth_acc_2433_nl = (z_out_901_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2433_nl = nl_AccumDotWidth_acc_2433_nl[9:0];
  assign nl_AccumDotWidth_acc_2434_nl = (z_out_608_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2434_nl = nl_AccumDotWidth_acc_2434_nl[9:0];
  assign nl_AccumDotWidth_acc_2435_nl = (z_out_862_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2435_nl = nl_AccumDotWidth_acc_2435_nl[9:0];
  assign AccumDotWidth_mux1h_886_nl = MUX1HOT_v_11_6_2(({{1{z_out_25[9]}}, z_out_25}),
      (signext_11_10(AccumDotWidth_acc_2432_nl)), (signext_11_10(AccumDotWidth_acc_2433_nl)),
      (signext_11_10(AccumDotWidth_acc_2434_nl)), (signext_11_10(AccumDotWidth_acc_2435_nl)),
      (MultLoop_acc_27_sdt[21:11]), {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_887_nl = MUX1HOT_v_11_5_2((nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm[10:0]),
      (z_out_901_29_7[12:2]), (z_out_608_29_7[12:2]), (z_out_862_29_7[12:2]), (MultLoop_acc_27_sdt[10:0]),
      {(fsm_output[3]) , AccumDotWidth_or_38_cse , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_331 = (AccumDotWidth_mux1h_885_nl) + ({(AccumDotWidth_mux1h_886_nl)
      , (AccumDotWidth_mux1h_887_nl)});
  assign z_out_331 = nl_z_out_331[21:0];
  assign AccumDotWidth_mux1h_888_nl = MUX1HOT_v_22_4_2(z_out_557, z_out_714, AccumDotWidth_acc_1877_itm,
      z_out_256, {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1434_nl = (z_out_616_29_7[21:0]) + (z_out_609_29_7[21:0]);
  assign MultLoop_acc_1434_nl = nl_MultLoop_acc_1434_nl[21:0];
  assign AccumDotWidth_mux1h_889_nl = MUX1HOT_v_22_4_2(z_out_559, z_out_717, z_out_794,
      (MultLoop_acc_1434_nl), {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_332 = (AccumDotWidth_mux1h_888_nl) + (AccumDotWidth_mux1h_889_nl);
  assign z_out_332 = nl_z_out_332[21:0];
  assign AccumDotWidth_mux1h_890_nl = MUX1HOT_v_22_6_2(z_out_368, z_out_390, z_out_560,
      z_out_716, z_out_795, z_out_487, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_891_nl = MUX1HOT_v_22_6_2(z_out_366, z_out_389, z_out_562,
      z_out_715, z_out_806, z_out_486, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_333 = (AccumDotWidth_mux1h_890_nl) + (AccumDotWidth_mux1h_891_nl);
  assign z_out_333 = nl_z_out_333[21:0];
  assign nl_MultLoop_acc_1435_nl = z_out_183_28_7 + z_out_182_28_7;
  assign MultLoop_acc_1435_nl = nl_MultLoop_acc_1435_nl[21:0];
  assign AccumDotWidth_mux1h_892_nl = MUX1HOT_v_22_4_2(z_out_739, z_out_736, z_out_718,
      (MultLoop_acc_1435_nl), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[343:336]));
  assign MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1436_nl = z_out_181_28_7 + (readslicef_29_22_7((MultLoop_43_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1436_nl = nl_MultLoop_acc_1436_nl[21:0];
  assign AccumDotWidth_mux1h_893_nl = MUX1HOT_v_22_4_2(z_out_737, (signext_22_21({z_out_27
      , (z_out_590_29_7[12:2])})), (signext_22_21({z_out_32 , (z_out_1133_29_9[10:0])})),
      (MultLoop_acc_1436_nl), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_334 = (AccumDotWidth_mux1h_892_nl) + (AccumDotWidth_mux1h_893_nl);
  assign z_out_334 = nl_z_out_334[21:0];
  assign nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[479:472]));
  assign MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[487:480]));
  assign MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1437_nl = (readslicef_29_22_7((MultLoop_60_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_61_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1437_nl = nl_MultLoop_acc_1437_nl[21:0];
  assign AccumDotWidth_mux1h_894_nl = MUX1HOT_v_22_5_2(z_out_711, z_out_736, z_out_719,
      (signext_22_21(z_out_1007_29_7[22:2])), (MultLoop_acc_1437_nl), {(fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[495:488]));
  assign MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[503:496]));
  assign MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1438_nl = (readslicef_29_22_7((MultLoop_62_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_63_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1438_nl = nl_MultLoop_acc_1438_nl[21:0];
  assign AccumDotWidth_mux1h_895_nl = MUX1HOT_v_22_5_2(z_out_702, z_out_732, z_out_720,
      (signext_22_21(z_out_970_29_7[22:2])), (MultLoop_acc_1438_nl), {(fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_335 = (AccumDotWidth_mux1h_894_nl) + (AccumDotWidth_mux1h_895_nl);
  assign z_out_335 = nl_z_out_335[21:0];
  assign nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[447:440]));
  assign MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[455:448]));
  assign MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1439_nl = (readslicef_29_22_7((MultLoop_56_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_57_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1439_nl = nl_MultLoop_acc_1439_nl[21:0];
  assign AccumDotWidth_mux1h_896_nl = MUX1HOT_v_22_6_2(z_out_706, z_out_397, z_out_424,
      z_out_422, z_out_693, (MultLoop_acc_1439_nl), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_897_nl = MUX1HOT_v_11_5_2((z_out_710[21:11]), (z_out_395[21:11]),
      ({{1{z_out_30[9]}}, z_out_30}), ({{1{z_out_33[9]}}, z_out_33}), (MultLoop_acc_1188_sdt[21:11]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_898_nl = MUX1HOT_v_11_6_2((z_out_710[10:0]), (z_out_395[10:0]),
      (z_out_908_29_7[12:2]), (z_out_609_29_7[12:2]), (z_out_883_29_7[12:2]), (MultLoop_acc_1188_sdt[10:0]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_336 = (AccumDotWidth_mux1h_896_nl) + ({(AccumDotWidth_mux1h_897_nl)
      , (AccumDotWidth_mux1h_898_nl)});
  assign z_out_336 = nl_z_out_336[21:0];
  assign nl_MultLoop_acc_1440_nl = z_out_168_28_7 + z_out_157_28_7;
  assign MultLoop_acc_1440_nl = nl_MultLoop_acc_1440_nl[21:0];
  assign AccumDotWidth_mux1h_899_nl = MUX1HOT_v_22_4_2(z_out_398, z_out_694, z_out_712,
      (MultLoop_acc_1440_nl), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2436_nl = (z_out_591_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2436_nl = nl_AccumDotWidth_acc_2436_nl[9:0];
  assign nl_AccumDotWidth_acc_2437_nl = (z_out_1137_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2437_nl = nl_AccumDotWidth_acc_2437_nl[9:0];
  assign nl_MultLoop_acc_1441_nl = (z_out_620_29_7[21:0]) + z_out_665_28_7;
  assign MultLoop_acc_1441_nl = nl_MultLoop_acc_1441_nl[21:0];
  assign AccumDotWidth_mux1h_900_nl = MUX1HOT_v_22_4_2(z_out_396, (signext_22_21({(AccumDotWidth_acc_2436_nl)
      , (z_out_591_29_7[12:2])})), (signext_22_21({(AccumDotWidth_acc_2437_nl) ,
      (z_out_1137_29_9[10:0])})), (MultLoop_acc_1441_nl), {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_337 = (AccumDotWidth_mux1h_899_nl) + (AccumDotWidth_mux1h_900_nl);
  assign z_out_337 = nl_z_out_337[21:0];
  assign nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[415:408]));
  assign MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[423:416]));
  assign MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1442_nl = (readslicef_29_22_7((MultLoop_52_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_53_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1442_nl = nl_MultLoop_acc_1442_nl[21:0];
  assign AccumDotWidth_mux1h_901_nl = MUX1HOT_v_22_4_2(z_out_399, z_out_734, z_out_424,
      (MultLoop_acc_1442_nl), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[431:424]));
  assign MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[439:432]));
  assign MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1443_nl = (readslicef_29_22_7((MultLoop_54_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_55_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1443_nl = nl_MultLoop_acc_1443_nl[21:0];
  assign AccumDotWidth_mux1h_902_nl = MUX1HOT_v_22_4_2(z_out_393, (signext_22_21({z_out_33
      , (z_out_989_29_9[10:0])})), (signext_22_21({z_out_27 , (z_out_1108_29_7[12:2])})),
      (MultLoop_acc_1443_nl), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_338 = (AccumDotWidth_mux1h_901_nl) + (AccumDotWidth_mux1h_902_nl);
  assign z_out_338 = nl_z_out_338[21:0];
  assign AccumDotWidth_mux1h_903_nl = MUX1HOT_v_11_7_2((signext_11_10(z_out_970_29_7[22:13])),
      (signext_11_10(z_out_955_29_7[22:13])), (signext_11_10(z_out_906_29_7[22:13])),
      ({{1{z_out_30[9]}}, z_out_30}), ({{1{z_out_27[9]}}, z_out_27}), (signext_11_10(z_out_1076_29_7[22:13])),
      (MultLoop_acc_1185_sdt[21:11]), {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[1])
      , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_904_nl = MUX1HOT_v_11_8_2((z_out_970_29_7[12:2]), (z_out_955_29_7[12:2]),
      (z_out_906_29_7[12:2]), (z_out_1028_29_7[12:2]), (z_out_1040_29_7[12:2]), (z_out_1076_29_7[12:2]),
      (z_out_1018_29_9[10:0]), (MultLoop_acc_1185_sdt[10:0]), {(fsm_output[2]) ,
      (fsm_output[6]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[527:520]));
  assign MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[535:528]));
  assign MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1444_nl = (readslicef_29_22_7((MultLoop_66_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_67_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1444_nl = nl_MultLoop_acc_1444_nl[21:0];
  assign AccumDotWidth_mux1h_905_nl = MUX1HOT_v_22_8_2((signext_22_21(z_out_908_29_7[22:2])),
      (signext_22_21(z_out_984_29_7[22:2])), (signext_22_21(z_out_895_29_7[22:2])),
      (signext_22_21(z_out_1051_29_7[22:2])), (signext_22_21(z_out_573_29_7[22:2])),
      (signext_22_21(z_out_587_29_7[22:2])), (signext_22_21(z_out_1125_29_7[22:2])),
      (MultLoop_acc_1444_nl), {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_339 = ({(AccumDotWidth_mux1h_903_nl) , (AccumDotWidth_mux1h_904_nl)})
      + (AccumDotWidth_mux1h_905_nl);
  assign z_out_339 = nl_z_out_339[21:0];
  assign AccumDotWidth_or_172_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[6]);
  assign AccumDotWidth_mux1h_906_nl = MUX1HOT_v_11_6_2((signext_11_10(z_out_944_29_7[22:13])),
      ({{1{z_out_30[9]}}, z_out_30}), ({{1{z_out_27[9]}}, z_out_27}), (signext_11_10(z_out_959_29_7[22:13])),
      ({{1{z_out_32[9]}}, z_out_32}), (MultLoop_acc_1193_sdt[21:11]), {(fsm_output[2])
      , (AccumDotWidth_or_172_nl) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_907_nl = MUX1HOT_v_11_8_2((z_out_944_29_7[12:2]), (z_out_1156_29_7[12:2]),
      (z_out_1033_29_9[10:0]), (z_out_618_29_7[12:2]), (z_out_959_29_7[12:2]), (z_out_588_29_7[12:2]),
      (z_out_1133_29_9[10:0]), (MultLoop_acc_1193_sdt[10:0]), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[399:392]));
  assign MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[407:400]));
  assign MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1445_nl = (readslicef_29_22_7((MultLoop_50_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_51_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1445_nl = nl_MultLoop_acc_1445_nl[21:0];
  assign AccumDotWidth_mux1h_908_nl = MUX1HOT_v_22_8_2((signext_22_21(z_out_1126_29_7[22:2])),
      (signext_22_21(z_out_1052_29_7[22:2])), (signext_22_21(z_out_1055_29_7[22:2])),
      (signext_22_21(z_out_954_29_7[22:2])), (signext_22_21(z_out_600_29_7[22:2])),
      (signext_22_21(z_out_595_29_7[22:2])), (signext_22_21(z_out_949_29_7[22:2])),
      (MultLoop_acc_1445_nl), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_340 = ({(AccumDotWidth_mux1h_906_nl) , (AccumDotWidth_mux1h_907_nl)})
      + (AccumDotWidth_mux1h_908_nl);
  assign z_out_340 = nl_z_out_340[21:0];
  assign nl_AccumDotWidth_acc_2438_nl = (z_out_1169_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[23:16]);
  assign AccumDotWidth_acc_2438_nl = nl_AccumDotWidth_acc_2438_nl[9:0];
  assign nl_AccumDotWidth_acc_2439_nl = (z_out_1039_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2439_nl = nl_AccumDotWidth_acc_2439_nl[9:0];
  assign nl_AccumDotWidth_acc_2440_nl = (z_out_1039_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2440_nl = nl_AccumDotWidth_acc_2440_nl[9:0];
  assign nl_AccumDotWidth_acc_2441_nl = (z_out_583_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2441_nl = nl_AccumDotWidth_acc_2441_nl[9:0];
  assign nl_AccumDotWidth_acc_2442_nl = (z_out_1137_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2442_nl = nl_AccumDotWidth_acc_2442_nl[9:0];
  assign AccumDotWidth_mux1h_909_nl = MUX1HOT_v_11_8_2((signext_11_10(z_out_978_29_9[20:11])),
      (signext_11_10(AccumDotWidth_acc_2438_nl)), (signext_11_10(AccumDotWidth_acc_2439_nl)),
      (signext_11_10(AccumDotWidth_acc_2440_nl)), (signext_11_10(z_out_1061_29_9[20:11])),
      (signext_11_10(AccumDotWidth_acc_2441_nl)), (signext_11_10(AccumDotWidth_acc_2442_nl)),
      (MultLoop_acc_1201_sdt[21:11]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_910_nl = MUX1HOT_v_11_7_2((z_out_978_29_9[10:0]), (z_out_1169_29_7[12:2]),
      (z_out_1039_29_7[12:2]), (z_out_1061_29_9[10:0]), (z_out_583_29_7[12:2]), (z_out_1137_29_9[10:0]),
      (MultLoop_acc_1201_sdt[10:0]), {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1446_nl = z_out_187_28_7 + z_out_186_28_7;
  assign MultLoop_acc_1446_nl = nl_MultLoop_acc_1446_nl[21:0];
  assign AccumDotWidth_mux1h_911_nl = MUX1HOT_v_22_8_2((signext_22_21(z_out_1010_29_7[22:2])),
      (signext_22_21(z_out_1184_29_7[22:2])), (signext_22_21(z_out_571_29_7[22:2])),
      (signext_22_21(z_out_568_29_7[22:2])), (signext_22_21(z_out_1149_29_7[22:2])),
      (signext_22_21(z_out_603_29_7[22:2])), (signext_22_21(z_out_1101_29_7[22:2])),
      (MultLoop_acc_1446_nl), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_341 = ({(AccumDotWidth_mux1h_909_nl) , (AccumDotWidth_mux1h_910_nl)})
      + (AccumDotWidth_mux1h_911_nl);
  assign z_out_341 = nl_z_out_341[21:0];
  assign nl_AccumDotWidth_acc_2443_nl = (z_out_892_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2443_nl = nl_AccumDotWidth_acc_2443_nl[9:0];
  assign nl_AccumDotWidth_acc_2444_nl = (z_out_868_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2444_nl = nl_AccumDotWidth_acc_2444_nl[9:0];
  assign nl_AccumDotWidth_acc_2445_nl = (z_out_1040_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2445_nl = nl_AccumDotWidth_acc_2445_nl[9:0];
  assign nl_AccumDotWidth_acc_2446_nl = (z_out_1043_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2446_nl = nl_AccumDotWidth_acc_2446_nl[9:0];
  assign nl_AccumDotWidth_acc_2447_nl = (z_out_591_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2447_nl = nl_AccumDotWidth_acc_2447_nl[9:0];
  assign nl_AccumDotWidth_acc_2448_nl = (z_out_863_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2448_nl = nl_AccumDotWidth_acc_2448_nl[9:0];
  assign AccumDotWidth_mux1h_912_nl = MUX1HOT_v_10_7_2((AccumDotWidth_acc_2443_nl),
      (AccumDotWidth_acc_2444_nl), (AccumDotWidth_acc_2445_nl), (AccumDotWidth_acc_2446_nl),
      (z_out_980_29_7[22:13]), (AccumDotWidth_acc_2447_nl), (AccumDotWidth_acc_2448_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_913_nl = MUX1HOT_v_11_7_2((z_out_892_29_7[12:2]), (z_out_868_29_7[12:2]),
      (z_out_1040_29_7[12:2]), (z_out_1043_29_7[12:2]), (z_out_980_29_7[12:2]), (z_out_591_29_7[12:2]),
      (z_out_863_29_7[12:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_914_nl = MUX1HOT_v_21_7_2(z_out_962_29_9, z_out_1139_29_9,
      (z_out_570_29_7[22:2]), (z_out_576_29_7[22:2]), (z_out_603_29_7[22:2]), (z_out_601_29_7[22:2]),
      (z_out_944_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_342 = conv_s2u_21_22({(AccumDotWidth_mux1h_912_nl) , (AccumDotWidth_mux1h_913_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_914_nl);
  assign z_out_342 = nl_z_out_342[21:0];
  assign nl_AccumDotWidth_acc_2449_nl = (z_out_1174_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2449_nl = nl_AccumDotWidth_acc_2449_nl[9:0];
  assign nl_AccumDotWidth_acc_2450_nl = (z_out_870_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2450_nl = nl_AccumDotWidth_acc_2450_nl[9:0];
  assign nl_AccumDotWidth_acc_2451_nl = (z_out_1026_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2451_nl = nl_AccumDotWidth_acc_2451_nl[9:0];
  assign nl_AccumDotWidth_acc_2452_nl = (z_out_1044_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2452_nl = nl_AccumDotWidth_acc_2452_nl[9:0];
  assign nl_AccumDotWidth_acc_2453_nl = (z_out_590_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2453_nl = nl_AccumDotWidth_acc_2453_nl[9:0];
  assign nl_AccumDotWidth_acc_2454_nl = (z_out_864_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2454_nl = nl_AccumDotWidth_acc_2454_nl[9:0];
  assign AccumDotWidth_mux1h_915_nl = MUX1HOT_v_10_7_2((AccumDotWidth_acc_2449_nl),
      (AccumDotWidth_acc_2450_nl), (AccumDotWidth_acc_2451_nl), (AccumDotWidth_acc_2452_nl),
      (z_out_1062_29_9[20:11]), (AccumDotWidth_acc_2453_nl), (AccumDotWidth_acc_2454_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_916_nl = MUX1HOT_v_11_7_2((z_out_1174_29_7[12:2]), (z_out_870_29_7[12:2]),
      (z_out_1026_29_7[12:2]), (z_out_1044_29_7[12:2]), (z_out_1062_29_9[10:0]),
      (z_out_590_29_7[12:2]), (z_out_864_29_7[12:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_917_nl = MUX1HOT_v_21_7_2(z_out_1141_29_9, (z_out_1127_29_7[22:2]),
      (z_out_1052_29_7[22:2]), (z_out_578_29_7[22:2]), (z_out_1146_29_7[22:2]), (z_out_602_29_7[22:2]),
      (z_out_940_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_343 = conv_s2u_21_22({(AccumDotWidth_mux1h_915_nl) , (AccumDotWidth_mux1h_916_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_917_nl);
  assign z_out_343 = nl_z_out_343[21:0];
  assign nl_AccumDotWidth_acc_2455_nl = (z_out_863_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[55:48]);
  assign AccumDotWidth_acc_2455_nl = nl_AccumDotWidth_acc_2455_nl[9:0];
  assign nl_AccumDotWidth_acc_2456_nl = (z_out_926_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2456_nl = nl_AccumDotWidth_acc_2456_nl[9:0];
  assign nl_AccumDotWidth_acc_2457_nl = (z_out_584_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2457_nl = nl_AccumDotWidth_acc_2457_nl[9:0];
  assign nl_AccumDotWidth_acc_2458_nl = (z_out_1159_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2458_nl = nl_AccumDotWidth_acc_2458_nl[9:0];
  assign AccumDotWidth_mux1h_918_nl = MUX1HOT_v_10_4_2((AccumDotWidth_acc_2455_nl),
      (AccumDotWidth_acc_2456_nl), (AccumDotWidth_acc_2457_nl), (AccumDotWidth_acc_2458_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_919_nl = MUX1HOT_v_11_4_2((z_out_863_29_7[12:2]), (z_out_926_29_7[12:2]),
      (z_out_584_29_7[12:2]), (z_out_1159_29_7[12:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_920_nl = MUX1HOT_v_21_4_2((z_out_879_29_7[22:2]), (z_out_1111_29_7[22:2]),
      (z_out_604_29_7[22:2]), (z_out_947_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_344 = conv_s2u_21_22({(AccumDotWidth_mux1h_918_nl) , (AccumDotWidth_mux1h_919_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_920_nl);
  assign z_out_344 = nl_z_out_344[21:0];
  assign nl_AccumDotWidth_acc_2459_nl = (z_out_1159_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[39:32]);
  assign AccumDotWidth_acc_2459_nl = nl_AccumDotWidth_acc_2459_nl[9:0];
  assign nl_AccumDotWidth_acc_2460_nl = (z_out_889_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2460_nl = nl_AccumDotWidth_acc_2460_nl[9:0];
  assign nl_AccumDotWidth_acc_2461_nl = (z_out_1042_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2461_nl = nl_AccumDotWidth_acc_2461_nl[9:0];
  assign nl_AccumDotWidth_acc_2462_nl = (z_out_594_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2462_nl = nl_AccumDotWidth_acc_2462_nl[9:0];
  assign nl_AccumDotWidth_acc_2463_nl = (z_out_1169_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2463_nl = nl_AccumDotWidth_acc_2463_nl[9:0];
  assign AccumDotWidth_mux1h_921_nl = MUX1HOT_v_10_7_2((z_out_955_29_7[22:13]), (AccumDotWidth_acc_2459_nl),
      (AccumDotWidth_acc_2460_nl), (AccumDotWidth_acc_2461_nl), (z_out_1060_29_9[20:11]),
      (AccumDotWidth_acc_2462_nl), (AccumDotWidth_acc_2463_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_922_nl = MUX1HOT_v_11_7_2((z_out_955_29_7[12:2]), (z_out_1159_29_7[12:2]),
      (z_out_889_29_7[12:2]), (z_out_1042_29_7[12:2]), (z_out_1060_29_9[10:0]), (z_out_594_29_7[12:2]),
      (z_out_1169_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_923_nl = MUX1HOT_v_21_6_2((z_out_1077_29_7[22:2]), (z_out_573_29_7[22:2]),
      (z_out_571_29_7[22:2]), (z_out_1158_29_7[22:2]), (z_out_599_29_7[22:2]), (z_out_945_29_7[22:2]),
      {(fsm_output[2]) , nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_345 = conv_s2u_21_22({(AccumDotWidth_mux1h_921_nl) , (AccumDotWidth_mux1h_922_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_923_nl);
  assign z_out_345 = nl_z_out_345[21:0];
  assign nl_AccumDotWidth_acc_2464_nl = conv_s2s_21_22(z_out_932_29_7[22:2]) + conv_s2s_21_22(z_out_616_29_7[22:2]);
  assign AccumDotWidth_acc_2464_nl = nl_AccumDotWidth_acc_2464_nl[21:0];
  assign AccumDotWidth_mux1h_924_nl = MUX1HOT_v_22_3_2(z_out_729, (AccumDotWidth_acc_2464_nl),
      z_out_694, {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2465_nl = (z_out_935_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2465_nl = nl_AccumDotWidth_acc_2465_nl[9:0];
  assign nl_AccumDotWidth_acc_2466_nl = (z_out_1128_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2466_nl = nl_AccumDotWidth_acc_2466_nl[9:0];
  assign nl_AccumDotWidth_acc_2467_nl = (z_out_882_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2467_nl = nl_AccumDotWidth_acc_2467_nl[9:0];
  assign AccumDotWidth_mux1h_925_nl = MUX1HOT_v_10_3_2((AccumDotWidth_acc_2465_nl),
      (AccumDotWidth_acc_2466_nl), (AccumDotWidth_acc_2467_nl), {(fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_926_nl = MUX1HOT_v_11_3_2((z_out_935_29_7[12:2]), (z_out_1128_29_7[12:2]),
      (z_out_882_29_7[12:2]), {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_346 = (AccumDotWidth_mux1h_924_nl) + conv_s2u_21_22({(AccumDotWidth_mux1h_925_nl)
      , (AccumDotWidth_mux1h_926_nl)});
  assign z_out_346 = nl_z_out_346[21:0];
  assign nl_AccumDotWidth_acc_2468_nl = (z_out_882_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2468_nl = nl_AccumDotWidth_acc_2468_nl[9:0];
  assign nl_AccumDotWidth_acc_2469_nl = (z_out_1036_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2469_nl = nl_AccumDotWidth_acc_2469_nl[9:0];
  assign nl_AccumDotWidth_acc_2470_nl = (z_out_587_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2470_nl = nl_AccumDotWidth_acc_2470_nl[9:0];
  assign nl_AccumDotWidth_acc_2471_nl = (z_out_1010_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2471_nl = nl_AccumDotWidth_acc_2471_nl[9:0];
  assign AccumDotWidth_mux1h_927_nl = MUX1HOT_v_21_7_2((z_out_1042_29_7[22:2]), (z_out_894_29_7[22:2]),
      ({(AccumDotWidth_acc_2468_nl) , (z_out_882_29_7[12:2])}), ({(AccumDotWidth_acc_2469_nl)
      , (z_out_1036_29_7[12:2])}), (z_out_1165_29_7[22:2]), ({(AccumDotWidth_acc_2470_nl)
      , (z_out_587_29_7[12:2])}), ({(AccumDotWidth_acc_2471_nl) , (z_out_1010_29_7[12:2])}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_928_nl = MUX1HOT_v_21_7_2((z_out_876_29_7[22:2]), (z_out_900_29_7[22:2]),
      (z_out_574_29_7[22:2]), (z_out_569_29_7[22:2]), (z_out_1097_29_7[22:2]), (z_out_597_29_7[22:2]),
      z_out_1135_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_347 = conv_s2u_21_22(AccumDotWidth_mux1h_927_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_928_nl);
  assign z_out_347 = nl_z_out_347[21:0];
  assign nl_AccumDotWidth_acc_2472_nl = conv_s2s_21_22(z_out_1003_29_9) + conv_s2s_21_22(z_out_879_29_7[22:2]);
  assign AccumDotWidth_acc_2472_nl = nl_AccumDotWidth_acc_2472_nl[21:0];
  assign AccumDotWidth_mux_96_nl = MUX_v_22_2_2(z_out_730, (AccumDotWidth_acc_2472_nl),
      fsm_output[6]);
  assign nl_AccumDotWidth_acc_2473_nl = (z_out_585_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2473_nl = nl_AccumDotWidth_acc_2473_nl[9:0];
  assign nl_AccumDotWidth_acc_2474_nl = (z_out_610_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2474_nl = nl_AccumDotWidth_acc_2474_nl[9:0];
  assign AccumDotWidth_mux_97_nl = MUX_v_10_2_2((AccumDotWidth_acc_2473_nl), (AccumDotWidth_acc_2474_nl),
      fsm_output[6]);
  assign AccumDotWidth_mux_98_nl = MUX_v_11_2_2((z_out_585_29_7[12:2]), (z_out_610_29_7[12:2]),
      fsm_output[6]);
  assign nl_z_out_348 = (AccumDotWidth_mux_96_nl) + conv_s2u_21_22({(AccumDotWidth_mux_97_nl)
      , (AccumDotWidth_mux_98_nl)});
  assign z_out_348 = nl_z_out_348[21:0];
  assign nl_AccumDotWidth_acc_2475_nl = (z_out_869_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2475_nl = nl_AccumDotWidth_acc_2475_nl[9:0];
  assign nl_AccumDotWidth_acc_2476_nl = (z_out_625_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2476_nl = nl_AccumDotWidth_acc_2476_nl[9:0];
  assign nl_AccumDotWidth_acc_2477_nl = (z_out_1036_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2477_nl = nl_AccumDotWidth_acc_2477_nl[9:0];
  assign nl_AccumDotWidth_acc_2478_nl = (z_out_1046_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2478_nl = nl_AccumDotWidth_acc_2478_nl[9:0];
  assign nl_AccumDotWidth_acc_2479_nl = (z_out_592_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2479_nl = nl_AccumDotWidth_acc_2479_nl[9:0];
  assign nl_AccumDotWidth_acc_2480_nl = (z_out_881_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2480_nl = nl_AccumDotWidth_acc_2480_nl[9:0];
  assign AccumDotWidth_mux1h_929_nl = MUX1HOT_v_10_7_2((AccumDotWidth_acc_2475_nl),
      (AccumDotWidth_acc_2476_nl), (AccumDotWidth_acc_2477_nl), (AccumDotWidth_acc_2478_nl),
      (z_out_1063_29_9[20:11]), (AccumDotWidth_acc_2479_nl), (AccumDotWidth_acc_2480_nl),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_930_nl = MUX1HOT_v_11_7_2((z_out_869_29_7[12:2]), (z_out_625_29_7[12:2]),
      (z_out_1036_29_7[12:2]), (z_out_1046_29_9[10:0]), (z_out_1063_29_9[10:0]),
      (z_out_592_29_7[12:2]), (z_out_881_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_931_nl = MUX1HOT_v_21_7_2((z_out_1109_29_7[22:2]), (z_out_919_29_7[22:2]),
      (z_out_569_29_7[22:2]), (z_out_577_29_7[22:2]), (z_out_1157_29_7[22:2]), (z_out_596_29_7[22:2]),
      (z_out_1087_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_349 = conv_s2u_21_22({(AccumDotWidth_mux1h_929_nl) , (AccumDotWidth_mux1h_930_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_931_nl);
  assign z_out_349 = nl_z_out_349[21:0];
  assign nl_AccumDotWidth_acc_2481_nl = (z_out_1031_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2481_nl = nl_AccumDotWidth_acc_2481_nl[9:0];
  assign nl_AccumDotWidth_acc_2482_nl = (z_out_1047_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2482_nl = nl_AccumDotWidth_acc_2482_nl[9:0];
  assign AccumDotWidth_mux1h_932_nl = MUX1HOT_v_21_7_2(z_out_1033_29_9, (z_out_1086_29_7[22:2]),
      (z_out_1114_29_7[22:2]), ({(AccumDotWidth_acc_2481_nl) , (z_out_1031_29_9[10:0])}),
      ({(AccumDotWidth_acc_2482_nl) , (z_out_1047_29_9[10:0])}), (z_out_938_29_7[22:2]),
      (z_out_1077_29_7[22:2]), {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_933_nl = MUX1HOT_v_21_7_2((z_out_1016_29_7[22:2]), (z_out_572_29_7[22:2]),
      (z_out_1117_29_7[22:2]), (z_out_1058_29_7[22:2]), (z_out_570_29_7[22:2]), (z_out_1180_29_7[22:2]),
      z_out_979_29_9, {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_z_out_350 = conv_s2u_21_22(AccumDotWidth_mux1h_932_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_933_nl);
  assign z_out_350 = nl_z_out_350[21:0];
  assign nl_AccumDotWidth_acc_2483_nl = (z_out_885_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2483_nl = nl_AccumDotWidth_acc_2483_nl[9:0];
  assign nl_AccumDotWidth_acc_2484_nl = (z_out_992_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2484_nl = nl_AccumDotWidth_acc_2484_nl[9:0];
  assign AccumDotWidth_mux1h_934_nl = MUX1HOT_v_21_7_2(z_out_1046_29_9, (z_out_899_29_7[22:2]),
      ({(AccumDotWidth_acc_2483_nl) , (z_out_885_29_7[12:2])}), ({(AccumDotWidth_acc_2484_nl)
      , (z_out_992_29_9[10:0])}), (z_out_1005_29_7[22:2]), (z_out_868_29_7[22:2]),
      (z_out_878_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_935_nl = MUX1HOT_v_21_6_2((z_out_900_29_7[22:2]), (z_out_897_29_7[22:2]),
      (z_out_568_29_7[22:2]), z_out_993_29_9, z_out_1144_29_9, (z_out_1027_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , AccumDotWidth_or_140_cse});
  assign nl_z_out_351 = conv_s2u_21_22(AccumDotWidth_mux1h_934_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_935_nl);
  assign z_out_351 = nl_z_out_351[21:0];
  assign AccumDotWidth_mux1h_936_nl = MUX1HOT_v_21_7_2((z_out_1025_29_7[22:2]), z_out_1143_29_9,
      (z_out_613_29_7[22:2]), (z_out_931_29_7[22:2]), ({z_out_31 , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0])}),
      (z_out_967_29_7[22:2]), (z_out_911_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_937_nl = MUX1HOT_v_21_7_2((z_out_1030_29_7[22:2]), (z_out_1076_29_7[22:2]),
      (z_out_908_29_7[22:2]), (z_out_937_29_7[22:2]), ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      (z_out_1107_29_7[22:2]), (z_out_1085_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_352 = conv_s2u_21_22(AccumDotWidth_mux1h_936_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_937_nl);
  assign z_out_352 = nl_z_out_352[21:0];
  assign nl_AccumDotWidth_acc_2485_nl = (z_out_1029_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2485_nl = nl_AccumDotWidth_acc_2485_nl[9:0];
  assign AccumDotWidth_mux1h_938_nl = MUX1HOT_v_21_7_2((z_out_1022_29_7[22:2]), (z_out_908_29_7[22:2]),
      ({(AccumDotWidth_acc_2485_nl) , (z_out_1029_29_7[12:2])}), (z_out_876_29_7[22:2]),
      (z_out_892_29_7[22:2]), (z_out_1034_29_7[22:2]), (z_out_1182_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_939_nl = MUX1HOT_v_21_7_2((z_out_614_29_7[22:2]), (z_out_898_29_7[22:2]),
      (z_out_1054_29_7[22:2]), (z_out_1025_29_7[22:2]), (z_out_854_29_7[22:2]), (z_out_894_29_7[22:2]),
      (z_out_1074_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_353 = conv_s2u_21_22(AccumDotWidth_mux1h_938_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_939_nl);
  assign z_out_353 = nl_z_out_353[21:0];
  assign nl_AccumDotWidth_acc_2486_nl = (z_out_624_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[7:0]);
  assign AccumDotWidth_acc_2486_nl = nl_AccumDotWidth_acc_2486_nl[9:0];
  assign nl_AccumDotWidth_acc_2487_nl = (z_out_621_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2487_nl = nl_AccumDotWidth_acc_2487_nl[9:0];
  assign AccumDotWidth_mux1h_940_nl = MUX1HOT_v_21_7_2((z_out_595_29_7[22:2]), ({(AccumDotWidth_acc_2486_nl)
      , (z_out_624_29_7[12:2])}), (z_out_608_29_7[22:2]), ({(AccumDotWidth_acc_2487_nl)
      , (z_out_621_29_7[12:2])}), (z_out_960_29_7[22:2]), (z_out_1130_29_7[22:2]),
      (z_out_581_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_941_nl = MUX1HOT_v_21_7_2((z_out_1159_29_7[22:2]), (z_out_912_29_7[22:2]),
      (z_out_870_29_7[22:2]), (z_out_599_29_7[22:2]), (z_out_598_29_7[22:2]), (z_out_1041_29_7[22:2]),
      (z_out_981_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_354 = conv_s2u_21_22(AccumDotWidth_mux1h_940_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_941_nl);
  assign z_out_354 = nl_z_out_354[21:0];
  assign nl_AccumDotWidth_acc_2488_nl = (z_out_1030_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2488_nl = nl_AccumDotWidth_acc_2488_nl[9:0];
  assign AccumDotWidth_mux1h_942_nl = MUX1HOT_v_21_7_2((z_out_893_29_7[22:2]), z_out_965_29_9,
      ({(AccumDotWidth_acc_2488_nl) , (z_out_1030_29_7[12:2])}), z_out_1063_29_9,
      (z_out_1069_29_7[22:2]), (z_out_1042_29_7[22:2]), (z_out_909_29_7[22:2]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_943_nl = MUX1HOT_v_21_7_2((z_out_918_29_7[22:2]), z_out_1136_29_9,
      (z_out_578_29_7[22:2]), (z_out_953_29_7[22:2]), (z_out_593_29_7[22:2]), (z_out_901_29_7[22:2]),
      (z_out_1084_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_355 = conv_s2u_21_22(AccumDotWidth_mux1h_942_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_943_nl);
  assign z_out_355 = nl_z_out_355[21:0];
  assign AccumDotWidth_mux1h_944_nl = MUX1HOT_v_21_7_2((z_out_1166_29_7[22:2]), (z_out_595_29_7[22:2]),
      (z_out_899_29_7[22:2]), (z_out_1171_29_7[22:2]), (z_out_1024_29_7[22:2]), (z_out_624_29_7[22:2]),
      (z_out_1172_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_945_nl = MUX1HOT_v_21_7_2((z_out_953_29_7[22:2]), (z_out_603_29_7[22:2]),
      (z_out_1025_29_7[22:2]), (z_out_1159_29_7[22:2]), (z_out_622_29_7[22:2]), (z_out_907_29_7[22:2]),
      (z_out_1086_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_356 = conv_s2u_21_22(AccumDotWidth_mux1h_944_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_945_nl);
  assign z_out_356 = nl_z_out_356[21:0];
  assign AccumDotWidth_mux1h_946_nl = MUX1HOT_v_21_7_2((z_out_974_29_7[22:2]), (z_out_1111_29_7[22:2]),
      (z_out_898_29_7[22:2]), (z_out_933_29_7[22:2]), (z_out_582_29_7[22:2]), (z_out_606_29_7[22:2]),
      (z_out_1163_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_947_nl = MUX1HOT_v_21_7_2((z_out_873_29_7[22:2]), (z_out_1115_29_7[22:2]),
      (z_out_1023_29_7[22:2]), (z_out_893_29_7[22:2]), z_out_1018_29_9, (z_out_1078_29_7[22:2]),
      (z_out_1090_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_357 = conv_s2u_21_22(AccumDotWidth_mux1h_946_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_947_nl);
  assign z_out_357 = nl_z_out_357[21:0];
  assign AccumDotWidth_mux1h_948_nl = MUX1HOT_v_21_7_2((z_out_995_29_7[22:2]), (z_out_1113_29_7[22:2]),
      (z_out_1016_29_7[22:2]), (z_out_1107_29_7[22:2]), (z_out_869_29_7[22:2]), (z_out_622_29_7[22:2]),
      (z_out_860_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_949_nl = MUX1HOT_v_21_7_2((z_out_927_29_7[22:2]), (z_out_1110_29_7[22:2]),
      (z_out_878_29_7[22:2]), (z_out_609_29_7[22:2]), (z_out_890_29_7[22:2]), z_out_904_29_9,
      (z_out_917_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_358 = conv_s2u_21_22(AccumDotWidth_mux1h_948_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_949_nl);
  assign z_out_358 = nl_z_out_358[21:0];
  assign AccumDotWidth_mux1h_950_nl = MUX1HOT_v_21_7_2((z_out_920_29_7[22:2]), (z_out_940_29_7[22:2]),
      (z_out_1181_29_7[22:2]), (z_out_867_29_7[22:2]), (z_out_1028_29_7[22:2]), (z_out_869_29_7[22:2]),
      (z_out_1107_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_951_nl = MUX1HOT_v_21_7_2((z_out_950_29_7[22:2]), (z_out_1124_29_7[22:2]),
      (z_out_864_29_7[22:2]), z_out_1032_29_9, (z_out_629_29_7[22:2]), (z_out_1024_29_7[22:2]),
      (z_out_968_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_359 = conv_s2u_21_22(AccumDotWidth_mux1h_950_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_951_nl);
  assign z_out_359 = nl_z_out_359[21:0];
  assign AccumDotWidth_mux1h_952_nl = MUX1HOT_v_21_7_2((z_out_601_29_7[22:2]), (z_out_597_29_7[22:2]),
      (z_out_609_29_7[22:2]), (z_out_1130_29_7[22:2]), z_out_1046_29_9, (z_out_876_29_7[22:2]),
      (z_out_572_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_953_nl = MUX1HOT_v_21_7_2((z_out_1015_29_7[22:2]), (z_out_592_29_7[22:2]),
      (z_out_872_29_7[22:2]), z_out_1018_29_9, (z_out_855_29_7[22:2]), (z_out_1025_29_7[22:2]),
      (z_out_980_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_360 = conv_s2u_21_22(AccumDotWidth_mux1h_952_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_953_nl);
  assign z_out_360 = nl_z_out_360[21:0];
  assign AccumDotWidth_mux1h_954_nl = MUX1HOT_v_21_7_2((z_out_915_29_7[22:2]), (z_out_1112_29_7[22:2]),
      (z_out_900_29_7[22:2]), (z_out_929_29_7[22:2]), (z_out_1147_29_7[22:2]), z_out_1031_29_9,
      (z_out_1186_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_955_nl = MUX1HOT_v_21_7_2(z_out_1066_29_9, (z_out_1119_29_7[22:2]),
      (z_out_1024_29_7[22:2]), (z_out_966_29_7[22:2]), (z_out_941_29_7[22:2]), (z_out_1014_29_7[22:2]),
      (z_out_1076_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_361 = conv_s2u_21_22(AccumDotWidth_mux1h_954_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_955_nl);
  assign z_out_361 = nl_z_out_361[21:0];
  assign AccumDotWidth_mux1h_956_nl = MUX1HOT_v_21_7_2((z_out_902_29_7[22:2]), (z_out_1182_29_7[22:2]),
      (z_out_879_29_7[22:2]), (z_out_1162_29_7[22:2]), z_out_1140_29_9, (z_out_1082_29_7[22:2]),
      (z_out_951_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_957_nl = MUX1HOT_v_21_7_2((z_out_1104_29_7[22:2]), (z_out_1049_29_7[22:2]),
      z_out_1018_29_9, (z_out_1187_29_7[22:2]), (z_out_1064_29_7[22:2]), (z_out_573_29_7[22:2]),
      z_out_1143_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_362 = conv_s2u_21_22(AccumDotWidth_mux1h_956_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_957_nl);
  assign z_out_362 = nl_z_out_362[21:0];
  assign AccumDotWidth_mux1h_958_nl = MUX1HOT_v_21_7_2((z_out_1113_29_7[22:2]), (z_out_905_29_7[22:2]),
      (z_out_967_29_7[22:2]), z_out_1140_29_9, (z_out_1001_29_7[22:2]), (z_out_922_29_7[22:2]),
      z_out_1062_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_959_nl = MUX1HOT_v_21_7_2((z_out_1157_29_7[22:2]), (z_out_1118_29_7[22:2]),
      (z_out_1079_29_7[22:2]), z_out_1020_29_9, z_out_1065_29_9, (z_out_925_29_7[22:2]),
      (z_out_902_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_363 = conv_s2u_21_22(AccumDotWidth_mux1h_958_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_959_nl);
  assign z_out_363 = nl_z_out_363[21:0];
  assign AccumDotWidth_mux1h_960_nl = MUX1HOT_v_21_7_2((z_out_856_29_7[22:2]), (z_out_1121_29_7[22:2]),
      (z_out_630_29_7[22:2]), (z_out_1054_29_7[22:2]), (z_out_1125_29_7[22:2]), (z_out_614_29_7[22:2]),
      (z_out_1058_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_961_nl = MUX1HOT_v_21_7_2((z_out_956_29_7[22:2]), (z_out_1116_29_7[22:2]),
      (z_out_1041_29_7[22:2]), (z_out_1024_29_7[22:2]), (z_out_1173_29_7[22:2]),
      (z_out_886_29_7[22:2]), (z_out_1022_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_364 = conv_s2u_21_22(AccumDotWidth_mux1h_960_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_961_nl);
  assign z_out_364 = nl_z_out_364[21:0];
  assign AccumDotWidth_mux1h_962_nl = MUX1HOT_v_21_7_2((z_out_1024_29_7[22:2]), (z_out_891_29_7[22:2]),
      (z_out_959_29_7[22:2]), (z_out_1168_29_7[22:2]), (z_out_581_29_7[22:2]), (z_out_861_29_7[22:2]),
      z_out_1065_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_963_nl = MUX1HOT_v_21_7_2(z_out_1033_29_9, (z_out_883_29_7[22:2]),
      (z_out_600_29_7[22:2]), (z_out_1156_29_7[22:2]), (z_out_998_29_7[22:2]), (z_out_969_29_7[22:2]),
      (z_out_573_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_365 = conv_s2u_21_22(AccumDotWidth_mux1h_962_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_963_nl);
  assign z_out_365 = nl_z_out_365[21:0];
  assign AccumDotWidth_mux1h_964_nl = MUX1HOT_v_21_7_2((z_out_1101_29_7[22:2]), (z_out_937_29_7[22:2]),
      (z_out_1177_29_7[22:2]), (z_out_1087_29_7[22:2]), (z_out_972_29_7[22:2]), (z_out_1001_29_7[22:2]),
      (z_out_854_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_965_nl = MUX1HOT_v_21_7_2((z_out_1093_29_7[22:2]), z_out_1062_29_9,
      (z_out_952_29_7[22:2]), (z_out_861_29_7[22:2]), (z_out_920_29_7[22:2]), (z_out_1115_29_7[22:2]),
      (z_out_957_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_366 = conv_s2u_21_22(AccumDotWidth_mux1h_964_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_965_nl);
  assign z_out_366 = nl_z_out_366[21:0];
  assign AccumDotWidth_mux1h_966_nl = MUX1HOT_v_21_7_2((z_out_1100_29_7[22:2]), (z_out_1180_29_7[22:2]),
      (z_out_1037_29_7[22:2]), (z_out_1108_29_7[22:2]), (z_out_913_29_7[22:2]), z_out_965_29_9,
      (z_out_1070_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_967_nl = MUX1HOT_v_21_7_2((z_out_1098_29_7[22:2]), (z_out_912_29_7[22:2]),
      (z_out_903_29_7[22:2]), (z_out_916_29_7[22:2]), (z_out_1090_29_7[22:2]), (z_out_981_29_7[22:2]),
      (z_out_1118_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_367 = conv_s2u_21_22(AccumDotWidth_mux1h_966_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_967_nl);
  assign z_out_367 = nl_z_out_367[21:0];
  assign AccumDotWidth_mux1h_968_nl = MUX1HOT_v_21_7_2((z_out_1027_29_7[22:2]), (z_out_914_29_7[22:2]),
      (z_out_1147_29_7[22:2]), (z_out_1050_29_7[22:2]), (z_out_863_29_7[22:2]), (z_out_957_29_7[22:2]),
      (z_out_958_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_969_nl = MUX1HOT_v_21_7_2((z_out_1022_29_7[22:2]), (z_out_1086_29_7[22:2]),
      (z_out_931_29_7[22:2]), (z_out_944_29_7[22:2]), (z_out_934_29_7[22:2]), (z_out_982_29_7[22:2]),
      (z_out_983_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_368 = conv_s2u_21_22(AccumDotWidth_mux1h_968_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_969_nl);
  assign z_out_368 = nl_z_out_368[21:0];
  assign AccumDotWidth_mux1h_970_nl = MUX1HOT_v_21_7_2((z_out_1096_29_7[22:2]), z_out_1138_29_9,
      (z_out_970_29_7[22:2]), z_out_1062_29_9, (z_out_1030_29_7[22:2]), (z_out_1088_29_7[22:2]),
      (z_out_908_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_971_nl = MUX1HOT_v_21_7_2((z_out_917_29_7[22:2]), z_out_989_29_9,
      (z_out_1076_29_7[22:2]), (z_out_941_29_7[22:2]), (z_out_625_29_7[22:2]), (z_out_580_29_7[22:2]),
      (z_out_592_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_369 = conv_s2u_21_22(AccumDotWidth_mux1h_970_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_971_nl);
  assign z_out_369 = nl_z_out_369[21:0];
  assign AccumDotWidth_mux1h_972_nl = MUX1HOT_v_21_7_2((z_out_1026_29_7[22:2]), (z_out_860_29_7[22:2]),
      z_out_1143_29_9, (z_out_1053_29_7[22:2]), (z_out_949_29_7[22:2]), (z_out_1007_29_7[22:2]),
      (z_out_1111_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_973_nl = MUX1HOT_v_21_7_2(z_out_1032_29_9, (z_out_593_29_7[22:2]),
      (z_out_586_29_7[22:2]), (z_out_1102_29_7[22:2]), (z_out_1164_29_7[22:2]), (z_out_1150_29_7[22:2]),
      (z_out_971_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_370 = conv_s2u_21_22(AccumDotWidth_mux1h_972_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_973_nl);
  assign z_out_370 = nl_z_out_370[21:0];
  assign AccumDotWidth_mux1h_974_nl = MUX1HOT_v_21_7_2((z_out_1095_29_7[22:2]), (z_out_954_29_7[22:2]),
      z_out_965_29_9, (z_out_1147_29_7[22:2]), (z_out_1075_29_7[22:2]), (z_out_618_29_7[22:2]),
      (z_out_1042_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_975_nl = MUX1HOT_v_21_7_2((z_out_1079_29_7[22:2]), (z_out_956_29_7[22:2]),
      (z_out_1111_29_7[22:2]), (z_out_940_29_7[22:2]), (z_out_1177_29_7[22:2]), (z_out_1044_29_7[22:2]),
      (z_out_866_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_371 = conv_s2u_21_22(AccumDotWidth_mux1h_974_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_975_nl);
  assign z_out_371 = nl_z_out_371[21:0];
  assign AccumDotWidth_mux1h_976_nl = MUX1HOT_v_21_7_2((z_out_981_29_7[22:2]), (z_out_959_29_7[22:2]),
      (z_out_587_29_7[22:2]), (z_out_1057_29_7[22:2]), (z_out_948_29_7[22:2]), (z_out_1119_29_7[22:2]),
      (z_out_602_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_977_nl = MUX1HOT_v_21_7_2((z_out_623_29_7[22:2]), (z_out_958_29_7[22:2]),
      (z_out_612_29_7[22:2]), (z_out_948_29_7[22:2]), (z_out_1167_29_7[22:2]), z_out_1134_29_9,
      (z_out_1008_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_372 = conv_s2u_21_22(AccumDotWidth_mux1h_976_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_977_nl);
  assign z_out_372 = nl_z_out_372[21:0];
  assign AccumDotWidth_mux1h_978_nl = MUX1HOT_v_21_7_2((z_out_864_29_7[22:2]), (z_out_982_29_7[22:2]),
      (z_out_961_29_7[22:2]), (z_out_1056_29_7[22:2]), (z_out_870_29_7[22:2]), (z_out_1076_29_7[22:2]),
      (z_out_575_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_979_nl = MUX1HOT_v_21_7_2((z_out_882_29_7[22:2]), (z_out_981_29_7[22:2]),
      (z_out_1114_29_7[22:2]), (z_out_947_29_7[22:2]), (z_out_880_29_7[22:2]), (z_out_996_29_7[22:2]),
      (z_out_985_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_373 = conv_s2u_21_22(AccumDotWidth_mux1h_978_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_979_nl);
  assign z_out_373 = nl_z_out_373[21:0];
  assign AccumDotWidth_mux1h_980_nl = MUX1HOT_v_21_7_2((z_out_943_29_7[22:2]), z_out_963_29_9,
      z_out_989_29_9, z_out_1060_29_9, (z_out_1122_29_7[22:2]), (z_out_889_29_7[22:2]),
      (z_out_952_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_981_nl = MUX1HOT_v_21_7_2(z_out_1067_29_9, (z_out_957_29_7[22:2]),
      (z_out_1110_29_7[22:2]), (z_out_943_29_7[22:2]), (z_out_1015_29_7[22:2]), (z_out_1023_29_7[22:2]),
      z_out_1066_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_374 = conv_s2u_21_22(AccumDotWidth_mux1h_980_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_981_nl);
  assign z_out_374 = nl_z_out_374[21:0];
  assign AccumDotWidth_mux1h_982_nl = MUX1HOT_v_21_7_2((z_out_960_29_7[22:2]), (z_out_584_29_7[22:2]),
      (z_out_1156_29_7[22:2]), z_out_1061_29_9, (z_out_964_29_7[22:2]), z_out_1065_29_9,
      z_out_1003_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_983_nl = MUX1HOT_v_21_7_2((z_out_961_29_7[22:2]), (z_out_620_29_7[22:2]),
      (z_out_923_29_7[22:2]), (z_out_945_29_7[22:2]), (z_out_1110_29_7[22:2]), (z_out_575_29_7[22:2]),
      (z_out_925_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_375 = conv_s2u_21_22(AccumDotWidth_mux1h_982_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_983_nl);
  assign z_out_375 = nl_z_out_375[21:0];
  assign AccumDotWidth_mux1h_984_nl = MUX1HOT_v_21_7_2((z_out_987_29_7[22:2]), (z_out_1099_29_7[22:2]),
      (z_out_596_29_7[22:2]), z_out_1142_29_9, (z_out_626_29_7[22:2]), (z_out_917_29_7[22:2]),
      (z_out_1164_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_985_nl = MUX1HOT_v_21_7_2(z_out_988_29_9, (z_out_998_29_7[22:2]),
      (z_out_1057_29_7[22:2]), (z_out_1123_29_7[22:2]), (z_out_977_29_7[22:2]), z_out_1142_29_9,
      (z_out_1088_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_376 = conv_s2u_21_22(AccumDotWidth_mux1h_984_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_985_nl);
  assign z_out_376 = nl_z_out_376[21:0];
  assign AccumDotWidth_mux1h_986_nl = MUX1HOT_v_21_7_2((z_out_980_29_7[22:2]), (z_out_952_29_7[22:2]),
      (z_out_1152_29_7[22:2]), (z_out_877_29_7[22:2]), (z_out_898_29_7[22:2]), (z_out_1071_29_7[22:2]),
      (z_out_601_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_987_nl = MUX1HOT_v_21_7_2((z_out_985_29_7[22:2]), (z_out_1054_29_7[22:2]),
      (z_out_941_29_7[22:2]), (z_out_926_29_7[22:2]), z_out_1031_29_9, (z_out_857_29_7[22:2]),
      (z_out_1014_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_377 = conv_s2u_21_22(AccumDotWidth_mux1h_986_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_987_nl);
  assign z_out_377 = nl_z_out_377[21:0];
  assign AccumDotWidth_mux1h_988_nl = MUX1HOT_v_21_7_2(z_out_965_29_9, (z_out_913_29_7[22:2]),
      z_out_1017_29_9, z_out_1141_29_9, (z_out_1074_29_7[22:2]), (z_out_1019_29_7[22:2]),
      (z_out_1054_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_989_nl = MUX1HOT_v_21_7_2((z_out_955_29_7[22:2]), (z_out_865_29_7[22:2]),
      (z_out_867_29_7[22:2]), (z_out_1122_29_7[22:2]), (z_out_592_29_7[22:2]), (z_out_916_29_7[22:2]),
      (z_out_937_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_378 = conv_s2u_21_22(AccumDotWidth_mux1h_988_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_989_nl);
  assign z_out_378 = nl_z_out_378[21:0];
  assign AccumDotWidth_mux1h_990_nl = MUX1HOT_v_21_7_2((z_out_969_29_7[22:2]), z_out_1137_29_9,
      z_out_988_29_9, (z_out_1161_29_7[22:2]), (z_out_984_29_7[22:2]), (z_out_859_29_7[22:2]),
      (z_out_995_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_991_nl = MUX1HOT_v_21_7_2((z_out_575_29_7[22:2]), (z_out_584_29_7[22:2]),
      z_out_1137_29_9, (z_out_1178_29_7[22:2]), (z_out_1038_29_7[22:2]), (z_out_971_29_7[22:2]),
      (z_out_932_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_379 = conv_s2u_21_22(AccumDotWidth_mux1h_990_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_991_nl);
  assign z_out_379 = nl_z_out_379[21:0];
  assign AccumDotWidth_mux1h_992_nl = MUX1HOT_v_21_7_2((z_out_984_29_7[22:2]), z_out_1141_29_9,
      (z_out_893_29_7[22:2]), (z_out_970_29_7[22:2]), (z_out_609_29_7[22:2]), (z_out_1113_29_7[22:2]),
      (z_out_1041_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_993_nl = MUX1HOT_v_21_7_2(z_out_992_29_9, (z_out_877_29_7[22:2]),
      (z_out_1071_29_7[22:2]), (z_out_951_29_7[22:2]), (z_out_605_29_7[22:2]), (z_out_1149_29_7[22:2]),
      (z_out_1117_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_380 = conv_s2u_21_22(AccumDotWidth_mux1h_992_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_993_nl);
  assign z_out_380 = nl_z_out_380[21:0];
  assign AccumDotWidth_mux1h_994_nl = MUX1HOT_v_21_7_2((z_out_1165_29_7[22:2]), (z_out_1153_29_7[22:2]),
      (z_out_1096_29_7[22:2]), (z_out_969_29_7[22:2]), (z_out_1127_29_7[22:2]), (z_out_958_29_7[22:2]),
      (z_out_921_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_995_nl = MUX1HOT_v_21_7_2((z_out_949_29_7[22:2]), (z_out_1147_29_7[22:2]),
      (z_out_856_29_7[22:2]), (z_out_950_29_7[22:2]), (z_out_911_29_7[22:2]), (z_out_986_29_7[22:2]),
      (z_out_1099_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_381 = conv_s2u_21_22(AccumDotWidth_mux1h_994_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_995_nl);
  assign z_out_381 = nl_z_out_381[21:0];
  assign AccumDotWidth_mux1h_996_nl = MUX1HOT_v_21_7_2((z_out_916_29_7[22:2]), (z_out_922_29_7[22:2]),
      (z_out_1115_29_7[22:2]), z_out_1144_29_9, (z_out_1151_29_7[22:2]), (z_out_946_29_7[22:2]),
      (z_out_959_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_997_nl = MUX1HOT_v_21_7_2(z_out_1006_29_9, (z_out_932_29_7[22:2]),
      (z_out_1148_29_7[22:2]), (z_out_1129_29_7[22:2]), (z_out_945_29_7[22:2]), z_out_1135_29_9,
      z_out_1136_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_382 = conv_s2u_21_22(AccumDotWidth_mux1h_996_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_997_nl);
  assign z_out_382 = nl_z_out_382[21:0];
  assign AccumDotWidth_mux1h_998_nl = MUX1HOT_v_21_7_2(z_out_979_29_9, (z_out_1154_29_7[22:2]),
      z_out_1188_29_9, (z_out_1082_29_7[22:2]), (z_out_903_29_7[22:2]), (z_out_1177_29_7[22:2]),
      (z_out_914_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_999_nl = MUX1HOT_v_21_7_2((z_out_1011_29_7[22:2]), (z_out_1146_29_7[22:2]),
      (z_out_877_29_7[22:2]), (z_out_925_29_7[22:2]), (z_out_1179_29_7[22:2]), (z_out_1111_29_7[22:2]),
      (z_out_1094_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_383 = conv_s2u_21_22(AccumDotWidth_mux1h_998_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_999_nl);
  assign z_out_383 = nl_z_out_383[21:0];
  assign AccumDotWidth_mux_99_nl = MUX_v_21_2_2((z_out_1103_29_7[22:2]), (z_out_592_29_7[22:2]),
      fsm_output[4]);
  assign AccumDotWidth_mux_100_nl = MUX_v_21_2_2((z_out_865_29_7[22:2]), (z_out_607_29_7[22:2]),
      fsm_output[4]);
  assign nl_z_out_384 = conv_s2u_21_22(AccumDotWidth_mux_99_nl) + conv_s2u_21_22(AccumDotWidth_mux_100_nl);
  assign z_out_384 = nl_z_out_384[21:0];
  assign AccumDotWidth_mux1h_1000_nl = MUX1HOT_v_21_7_2((z_out_945_29_7[22:2]), (z_out_1043_29_7[22:2]),
      (z_out_983_29_7[22:2]), (z_out_974_29_7[22:2]), (z_out_1080_29_7[22:2]), (z_out_948_29_7[22:2]),
      (z_out_964_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1001_nl = MUX1HOT_v_21_7_2((z_out_946_29_7[22:2]), (z_out_866_29_7[22:2]),
      (z_out_1106_29_7[22:2]), (z_out_902_29_7[22:2]), (z_out_858_29_7[22:2]), (z_out_1125_29_7[22:2]),
      z_out_1059_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_385 = conv_s2u_21_22(AccumDotWidth_mux1h_1000_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1001_nl);
  assign z_out_385 = nl_z_out_385[21:0];
  assign AccumDotWidth_mux1h_1002_nl = MUX1HOT_v_21_7_2((z_out_991_29_7[22:2]), (z_out_1104_29_7[22:2]),
      (z_out_1184_29_7[22:2]), (z_out_595_29_7[22:2]), (z_out_875_29_7[22:2]), (z_out_1172_29_7[22:2]),
      (z_out_910_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1003_nl = MUX1HOT_v_21_7_2((z_out_937_29_7[22:2]), (z_out_950_29_7[22:2]),
      (z_out_862_29_7[22:2]), (z_out_1051_29_7[22:2]), (z_out_923_29_7[22:2]), (z_out_1087_29_7[22:2]),
      (z_out_1100_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_386 = conv_s2u_21_22(AccumDotWidth_mux1h_1002_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1003_nl);
  assign z_out_386 = nl_z_out_386[21:0];
  assign AccumDotWidth_mux1h_1004_nl = MUX1HOT_v_21_7_2((z_out_1158_29_7[22:2]),
      (z_out_1152_29_7[22:2]), (z_out_1116_29_7[22:2]), (z_out_1160_29_7[22:2]),
      (z_out_1002_29_7[22:2]), (z_out_888_29_7[22:2]), (z_out_587_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1005_nl = MUX1HOT_v_21_7_2((z_out_590_29_7[22:2]), (z_out_1151_29_7[22:2]),
      (z_out_1149_29_7[22:2]), (z_out_1177_29_7[22:2]), (z_out_1187_29_7[22:2]),
      (z_out_1030_29_7[22:2]), (z_out_880_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_387 = conv_s2u_21_22(AccumDotWidth_mux1h_1004_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1005_nl);
  assign z_out_387 = nl_z_out_387[21:0];
  assign AccumDotWidth_mux1h_1006_nl = MUX1HOT_v_21_6_2((z_out_964_29_7[22:2]), (z_out_919_29_7[22:2]),
      (z_out_1164_29_7[22:2]), (z_out_1155_29_7[22:2]), (z_out_1123_29_7[22:2]),
      (z_out_928_29_7[22:2]), {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1007_nl = MUX1HOT_v_21_6_2((z_out_939_29_7[22:2]), (z_out_1082_29_7[22:2]),
      (z_out_1104_29_7[22:2]), (z_out_1096_29_7[22:2]), (z_out_1009_29_7[22:2]),
      (z_out_1103_29_7[22:2]), {AccumDotWidth_or_153_cse , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_z_out_388 = conv_s2u_21_22(AccumDotWidth_mux1h_1006_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1007_nl);
  assign z_out_388 = nl_z_out_388[21:0];
  assign AccumDotWidth_mux1h_1008_nl = MUX1HOT_v_21_7_2(z_out_942_29_9, (z_out_990_29_7[22:2]),
      (z_out_1145_29_7[22:2]), (z_out_606_29_7[22:2]), (z_out_909_29_7[22:2]), (z_out_571_29_7[22:2]),
      (z_out_618_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1009_nl = MUX1HOT_v_21_7_2((z_out_949_29_7[22:2]), (z_out_1052_29_7[22:2]),
      (z_out_853_29_7[22:2]), (z_out_1119_29_7[22:2]), (z_out_1082_29_7[22:2]), (z_out_863_29_7[22:2]),
      (z_out_898_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_389 = conv_s2u_21_22(AccumDotWidth_mux1h_1008_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1009_nl);
  assign z_out_389 = nl_z_out_389[21:0];
  assign AccumDotWidth_mux1h_1010_nl = MUX1HOT_v_21_7_2((z_out_1092_29_7[22:2]),
      (z_out_1016_29_7[22:2]), z_out_1003_29_9, (z_out_574_29_7[22:2]), z_out_1143_29_9,
      (z_out_1186_29_7[22:2]), (z_out_584_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1011_nl = MUX1HOT_v_21_7_2((z_out_1179_29_7[22:2]),
      (z_out_1012_29_7[22:2]), (z_out_1064_29_7[22:2]), z_out_962_29_9, (z_out_952_29_7[22:2]),
      z_out_1020_29_9, (z_out_615_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_390 = conv_s2u_21_22(AccumDotWidth_mux1h_1010_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1011_nl);
  assign z_out_390 = nl_z_out_390[21:0];
  assign AccumDotWidth_mux1h_1012_nl = MUX1HOT_v_21_7_2((z_out_959_29_7[22:2]), (z_out_1013_29_7[22:2]),
      (z_out_977_29_7[22:2]), (z_out_598_29_7[22:2]), (z_out_971_29_7[22:2]), z_out_1143_29_9,
      (z_out_588_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1013_nl = MUX1HOT_v_21_7_2((z_out_627_29_7[22:2]), z_out_1018_29_9,
      (z_out_925_29_7[22:2]), (z_out_1111_29_7[22:2]), (z_out_902_29_7[22:2]), z_out_979_29_9,
      (z_out_608_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_391 = conv_s2u_21_22(AccumDotWidth_mux1h_1012_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1013_nl);
  assign z_out_391 = nl_z_out_391[21:0];
  assign AccumDotWidth_mux1h_1014_nl = MUX1HOT_v_21_7_2((z_out_1034_29_7[22:2]),
      z_out_1132_29_9, z_out_1134_29_9, (z_out_575_29_7[22:2]), (z_out_1102_29_7[22:2]),
      (z_out_933_29_7[22:2]), (z_out_938_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1015_nl = MUX1HOT_v_21_7_2((z_out_1064_29_7[22:2]),
      (z_out_957_29_7[22:2]), (z_out_614_29_7[22:2]), z_out_963_29_9, (z_out_1160_29_7[22:2]),
      (z_out_920_29_7[22:2]), (z_out_1106_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_392 = conv_s2u_21_22(AccumDotWidth_mux1h_1014_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1015_nl);
  assign z_out_392 = nl_z_out_392[21:0];
  assign AccumDotWidth_mux1h_1016_nl = MUX1HOT_v_21_7_2((z_out_1150_29_7[22:2]),
      (z_out_600_29_7[22:2]), (z_out_1126_29_7[22:2]), z_out_942_29_9, (z_out_1052_29_7[22:2]),
      (z_out_1057_29_7[22:2]), (z_out_913_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1017_nl = MUX1HOT_v_21_7_2((z_out_948_29_7[22:2]), (z_out_1089_29_7[22:2]),
      (z_out_617_29_7[22:2]), (z_out_1183_29_7[22:2]), z_out_993_29_9, (z_out_941_29_7[22:2]),
      (z_out_1092_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_393 = conv_s2u_21_22(AccumDotWidth_mux1h_1016_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1017_nl);
  assign z_out_393 = nl_z_out_393[21:0];
  assign AccumDotWidth_mux1h_1018_nl = MUX1HOT_v_21_7_2((z_out_1155_29_7[22:2]),
      z_out_989_29_9, (z_out_968_29_7[22:2]), (z_out_986_29_7[22:2]), (z_out_597_29_7[22:2]),
      (z_out_1163_29_7[22:2]), (z_out_888_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1019_nl = MUX1HOT_v_21_7_2((z_out_1145_29_7[22:2]),
      (z_out_619_29_7[22:2]), (z_out_873_29_7[22:2]), z_out_1048_29_9, (z_out_1117_29_7[22:2]),
      (z_out_1085_29_7[22:2]), (z_out_975_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_394 = conv_s2u_21_22(AccumDotWidth_mux1h_1018_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1019_nl);
  assign z_out_394 = nl_z_out_394[21:0];
  assign AccumDotWidth_mux1h_1020_nl = MUX1HOT_v_21_7_2((z_out_1097_29_7[22:2]),
      (z_out_1051_29_7[22:2]), (z_out_1151_29_7[22:2]), z_out_979_29_9, (z_out_579_29_7[22:2]),
      z_out_1060_29_9, (z_out_900_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1021_nl = MUX1HOT_v_21_7_2(z_out_1138_29_9, (z_out_1058_29_7[22:2]),
      (z_out_926_29_7[22:2]), (z_out_1022_29_7[22:2]), (z_out_995_29_7[22:2]), (z_out_1099_29_7[22:2]),
      (z_out_590_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_395 = conv_s2u_21_22(AccumDotWidth_mux1h_1020_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1021_nl);
  assign z_out_395 = nl_z_out_395[21:0];
  assign AccumDotWidth_mux1h_1022_nl = MUX1HOT_v_21_7_2((z_out_604_29_7[22:2]), (z_out_1091_29_7[22:2]),
      (z_out_1002_29_7[22:2]), (z_out_1069_29_7[22:2]), (z_out_1068_29_7[22:2]),
      (z_out_581_29_7[22:2]), z_out_1020_29_9, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1023_nl = MUX1HOT_v_21_7_2((z_out_1080_29_7[22:2]),
      (z_out_1090_29_7[22:2]), (z_out_1045_29_7[22:2]), (z_out_588_29_7[22:2]), (z_out_1175_29_7[22:2]),
      (z_out_862_29_7[22:2]), (z_out_972_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_396 = conv_s2u_21_22(AccumDotWidth_mux1h_1022_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1023_nl);
  assign z_out_396 = nl_z_out_396[21:0];
  assign AccumDotWidth_mux1h_1024_nl = MUX1HOT_v_21_7_2((z_out_986_29_7[22:2]), (z_out_1082_29_7[22:2]),
      (z_out_960_29_7[22:2]), z_out_1017_29_9, (z_out_578_29_7[22:2]), (z_out_1181_29_7[22:2]),
      (z_out_1034_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1025_nl = MUX1HOT_v_21_7_2((z_out_628_29_7[22:2]), (z_out_1081_29_7[22:2]),
      (z_out_1113_29_7[22:2]), (z_out_1088_29_7[22:2]), (z_out_961_29_7[22:2]), z_out_1017_29_9,
      (z_out_899_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_397 = conv_s2u_21_22(AccumDotWidth_mux1h_1024_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1025_nl);
  assign z_out_397 = nl_z_out_397[21:0];
  assign AccumDotWidth_mux1h_1026_nl = MUX1HOT_v_21_7_2(z_out_1066_29_9, (z_out_909_29_7[22:2]),
      (z_out_974_29_7[22:2]), (z_out_1045_29_7[22:2]), (z_out_1008_29_7[22:2]), (z_out_612_29_7[22:2]),
      z_out_965_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1027_nl = MUX1HOT_v_21_7_2((z_out_1056_29_7[22:2]),
      (z_out_861_29_7[22:2]), (z_out_1075_29_7[22:2]), z_out_978_29_9, (z_out_613_29_7[22:2]),
      (z_out_885_29_7[22:2]), (z_out_891_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_398 = conv_s2u_21_22(AccumDotWidth_mux1h_1026_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1027_nl);
  assign z_out_398 = nl_z_out_398[21:0];
  assign AccumDotWidth_mux1h_1028_nl = MUX1HOT_v_21_7_2((z_out_1054_29_7[22:2]),
      (z_out_910_29_7[22:2]), z_out_1139_29_9, (z_out_619_29_7[22:2]), (z_out_895_29_7[22:2]),
      z_out_992_29_9, (z_out_1174_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1029_nl = MUX1HOT_v_21_7_2((z_out_1055_29_7[22:2]),
      (z_out_858_29_7[22:2]), (z_out_615_29_7[22:2]), (z_out_977_29_7[22:2]), z_out_1033_29_9,
      (z_out_1069_29_7[22:2]), (z_out_580_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_399 = conv_s2u_21_22(AccumDotWidth_mux1h_1028_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1029_nl);
  assign z_out_399 = nl_z_out_399[21:0];
  assign AccumDotWidth_mux1h_1030_nl = MUX1HOT_v_21_6_2((z_out_1038_29_7[22:2]),
      (z_out_987_29_7[22:2]), (z_out_995_29_7[22:2]), (z_out_985_29_7[22:2]), z_out_1033_29_9,
      (z_out_591_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1031_nl = MUX1HOT_v_21_6_2((z_out_1075_29_7[22:2]),
      (z_out_1112_29_7[22:2]), (z_out_891_29_7[22:2]), (z_out_1043_29_7[22:2]), (z_out_1011_29_7[22:2]),
      (z_out_616_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_400 = conv_s2u_21_22(AccumDotWidth_mux1h_1030_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1031_nl);
  assign z_out_400 = nl_z_out_400[21:0];
  assign AccumDotWidth_mux1h_1032_nl = MUX1HOT_v_21_4_2((z_out_960_29_7[22:2]), (z_out_1146_29_7[22:2]),
      (z_out_899_29_7[22:2]), (z_out_1180_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1033_nl = MUX1HOT_v_21_4_2(z_out_1004_29_9, (z_out_948_29_7[22:2]),
      (z_out_614_29_7[22:2]), z_out_989_29_9, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign nl_z_out_401 = conv_s2u_21_22(AccumDotWidth_mux1h_1032_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1033_nl);
  assign z_out_401 = nl_z_out_401[21:0];
  assign AccumDotWidth_mux1h_1034_nl = MUX1HOT_v_22_5_2(({{1{z_out_1048_29_9[20]}},
      z_out_1048_29_9}), (signext_22_21(z_out_601_29_7[22:2])), (signext_22_21(z_out_587_29_7[22:2])),
      z_out_360, (signext_22_21(z_out_1112_29_7[22:2])), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign nl_AccumDotWidth_acc_2489_nl = (z_out_584_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2489_nl = nl_AccumDotWidth_acc_2489_nl[9:0];
  assign AccumDotWidth_mux1h_1035_nl = MUX1HOT_v_21_5_2((z_out_1073_29_7[22:2]),
      z_out_1060_29_9, (z_out_1089_29_7[22:2]), ({(AccumDotWidth_acc_2489_nl) , (z_out_584_29_7[12:2])}),
      (z_out_1148_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6])});
  assign nl_z_out_402 = (AccumDotWidth_mux1h_1034_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1035_nl);
  assign z_out_402 = nl_z_out_402[21:0];
  assign AccumDotWidth_mux1h_1036_nl = MUX1HOT_v_21_4_2((z_out_1131_29_7[22:2]),
      (z_out_1091_29_7[22:2]), (z_out_889_29_7[22:2]), (z_out_1070_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1037_nl = MUX1HOT_v_21_4_2(z_out_1017_29_9, (z_out_895_29_7[22:2]),
      (z_out_615_29_7[22:2]), z_out_1059_29_9, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign nl_z_out_403 = conv_s2u_21_22(AccumDotWidth_mux1h_1036_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1037_nl);
  assign z_out_403 = nl_z_out_403[21:0];
  assign AccumDotWidth_mux1h_1038_nl = MUX1HOT_v_21_4_2((z_out_1064_29_7[22:2]),
      (z_out_1086_29_7[22:2]), (z_out_589_29_7[22:2]), (z_out_853_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1039_nl = MUX1HOT_v_21_4_2((z_out_1051_29_7[22:2]),
      (z_out_1131_29_7[22:2]), (z_out_617_29_7[22:2]), (z_out_959_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign nl_z_out_404 = conv_s2u_21_22(AccumDotWidth_mux1h_1038_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1039_nl);
  assign z_out_404 = nl_z_out_404[21:0];
  assign AccumDotWidth_mux1h_1040_nl = MUX1HOT_v_21_4_2((z_out_1034_29_7[22:2]),
      (z_out_1108_29_7[22:2]), (z_out_884_29_7[22:2]), (z_out_975_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1041_nl = MUX1HOT_v_21_4_2(z_out_1063_29_9, (z_out_1012_29_7[22:2]),
      (z_out_616_29_7[22:2]), (z_out_918_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign nl_z_out_405 = conv_s2u_21_22(AccumDotWidth_mux1h_1040_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1041_nl);
  assign z_out_405 = nl_z_out_405[21:0];
  assign AccumDotWidth_mux_101_nl = MUX_v_21_2_2(z_out_1140_29_9, (z_out_582_29_7[22:2]),
      fsm_output[4]);
  assign AccumDotWidth_mux_102_nl = MUX_v_21_2_2((z_out_1009_29_7[22:2]), (z_out_611_29_7[22:2]),
      fsm_output[4]);
  assign nl_z_out_406 = conv_s2u_21_22(AccumDotWidth_mux_101_nl) + conv_s2u_21_22(AccumDotWidth_mux_102_nl);
  assign z_out_406 = nl_z_out_406[21:0];
  assign nl_AccumDotWidth_acc_2490_nl = conv_s2s_21_22(z_out_988_29_9) + conv_s2s_21_22(z_out_1048_29_9);
  assign AccumDotWidth_acc_2490_nl = nl_AccumDotWidth_acc_2490_nl[21:0];
  assign AccumDotWidth_mux1h_1042_nl = MUX1HOT_v_22_5_2((signext_22_21(z_out_1107_29_7[22:2])),
      ({{1{z_out_1133_29_9[20]}}, z_out_1133_29_9}), (signext_22_21(z_out_890_29_7[22:2])),
      (AccumDotWidth_acc_2490_nl), (signext_22_21(z_out_910_29_7[22:2])), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign nl_AccumDotWidth_acc_2491_nl = (z_out_899_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2491_nl = nl_AccumDotWidth_acc_2491_nl[9:0];
  assign AccumDotWidth_mux1h_1043_nl = MUX1HOT_v_21_5_2((z_out_1014_29_7[22:2]),
      z_out_1020_29_9, (z_out_610_29_7[22:2]), ({(AccumDotWidth_acc_2491_nl) , (z_out_899_29_7[12:2])}),
      (z_out_1174_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6])});
  assign nl_z_out_407 = (AccumDotWidth_mux1h_1042_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1043_nl);
  assign z_out_407 = nl_z_out_407[21:0];
  assign AccumDotWidth_mux1h_1044_nl = MUX1HOT_v_21_4_2((z_out_881_29_7[22:2]), (z_out_1090_29_7[22:2]),
      (z_out_888_29_7[22:2]), (z_out_983_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1045_nl = MUX1HOT_v_21_4_2(z_out_1137_29_9, (z_out_910_29_7[22:2]),
      (z_out_608_29_7[22:2]), (z_out_980_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign nl_z_out_408 = conv_s2u_21_22(AccumDotWidth_mux1h_1044_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1045_nl);
  assign z_out_408 = nl_z_out_408[21:0];
  assign AccumDotWidth_mux_103_nl = MUX_v_21_2_2((z_out_1088_29_7[22:2]), (z_out_594_29_7[22:2]),
      fsm_output[4]);
  assign AccumDotWidth_mux_104_nl = MUX_v_21_2_2((z_out_1107_29_7[22:2]), (z_out_613_29_7[22:2]),
      fsm_output[4]);
  assign nl_z_out_409 = conv_s2u_21_22(AccumDotWidth_mux_103_nl) + conv_s2u_21_22(AccumDotWidth_mux_104_nl);
  assign z_out_409 = nl_z_out_409[21:0];
  assign AccumDotWidth_mux_105_nl = MUX_v_21_2_2((z_out_1083_29_7[22:2]), (z_out_882_29_7[22:2]),
      fsm_output[4]);
  assign AccumDotWidth_mux_106_nl = MUX_v_21_2_2((z_out_913_29_7[22:2]), z_out_988_29_9,
      fsm_output[4]);
  assign nl_z_out_410 = conv_s2u_21_22(AccumDotWidth_mux_105_nl) + conv_s2u_21_22(AccumDotWidth_mux_106_nl);
  assign z_out_410 = nl_z_out_410[21:0];
  assign AccumDotWidth_mux_107_nl = MUX_v_21_2_2((z_out_1122_29_7[22:2]), (z_out_593_29_7[22:2]),
      fsm_output[4]);
  assign AccumDotWidth_mux_108_nl = MUX_v_21_2_2((z_out_1015_29_7[22:2]), (z_out_1081_29_7[22:2]),
      fsm_output[4]);
  assign nl_z_out_411 = conv_s2u_21_22(AccumDotWidth_mux_107_nl) + conv_s2u_21_22(AccumDotWidth_mux_108_nl);
  assign z_out_411 = nl_z_out_411[21:0];
  assign AccumDotWidth_mux1h_1046_nl = MUX1HOT_v_21_5_2((z_out_911_29_7[22:2]), (z_out_606_29_7[22:2]),
      (z_out_959_29_7[22:2]), (z_out_1178_29_7[22:2]), (z_out_568_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1047_nl = MUX1HOT_v_21_5_2((z_out_1084_29_7[22:2]),
      (z_out_1050_29_7[22:2]), (z_out_1116_29_7[22:2]), (z_out_1010_29_7[22:2]),
      (z_out_961_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_412 = conv_s2u_21_22(AccumDotWidth_mux1h_1046_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1047_nl);
  assign z_out_412 = nl_z_out_412[21:0];
  assign AccumDotWidth_mux1h_1048_nl = MUX1HOT_v_21_5_2((z_out_583_29_7[22:2]), (z_out_1166_29_7[22:2]),
      (z_out_958_29_7[22:2]), (z_out_1131_29_7[22:2]), (z_out_1168_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1049_nl = MUX1HOT_v_21_5_2((z_out_980_29_7[22:2]), (z_out_1178_29_7[22:2]),
      (z_out_1115_29_7[22:2]), (z_out_1038_29_7[22:2]), (z_out_1081_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_413 = conv_s2u_21_22(AccumDotWidth_mux1h_1048_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1049_nl);
  assign z_out_413 = nl_z_out_413[21:0];
  assign AccumDotWidth_mux1h_1050_nl = MUX1HOT_v_21_6_2((z_out_984_29_7[22:2]), (z_out_881_29_7[22:2]),
      (z_out_1153_29_7[22:2]), (z_out_569_29_7[22:2]), (z_out_1052_29_7[22:2]), z_out_1063_29_9,
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1051_nl = MUX1HOT_v_21_6_2((z_out_626_29_7[22:2]), (z_out_1102_29_7[22:2]),
      (z_out_1124_29_7[22:2]), z_out_1004_29_9, (z_out_1145_29_7[22:2]), z_out_988_29_9,
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_414 = conv_s2u_21_22(AccumDotWidth_mux1h_1050_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1051_nl);
  assign z_out_414 = nl_z_out_414[21:0];
  assign AccumDotWidth_mux1h_1052_nl = MUX1HOT_v_21_4_2((z_out_1093_29_7[22:2]),
      (z_out_1162_29_7[22:2]), (z_out_923_29_7[22:2]), (z_out_874_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1053_nl = MUX1HOT_v_21_3_2((z_out_951_29_7[22:2]), (z_out_1176_29_7[22:2]),
      (z_out_1025_29_7[22:2]), {MultLoop_or_89_cse , (fsm_output[3]) , (fsm_output[7])});
  assign nl_z_out_415 = conv_s2u_21_22(AccumDotWidth_mux1h_1052_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1053_nl);
  assign z_out_415 = nl_z_out_415[21:0];
  assign AccumDotWidth_mux1h_1054_nl = MUX1HOT_v_21_4_2((z_out_996_29_7[22:2]), z_out_1144_29_9,
      (z_out_865_29_7[22:2]), z_out_1188_29_9, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1055_nl = MUX1HOT_v_21_4_2((z_out_1045_29_7[22:2]),
      (z_out_588_29_7[22:2]), (z_out_864_29_7[22:2]), (z_out_1075_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_416 = conv_s2u_21_22(AccumDotWidth_mux1h_1054_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1055_nl);
  assign z_out_416 = nl_z_out_416[21:0];
  assign AccumDotWidth_mux1h_1056_nl = MUX1HOT_v_21_6_2(z_out_942_29_9, (z_out_604_29_7[22:2]),
      (z_out_1154_29_7[22:2]), (z_out_1159_29_7[22:2]), (z_out_954_29_7[22:2]), (z_out_1171_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1057_nl = MUX1HOT_v_21_6_2((z_out_570_29_7[22:2]), (z_out_1056_29_7[22:2]),
      (z_out_1127_29_7[22:2]), (z_out_924_29_7[22:2]), (z_out_600_29_7[22:2]), (z_out_1089_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_417 = conv_s2u_21_22(AccumDotWidth_mux1h_1056_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1057_nl);
  assign z_out_417 = nl_z_out_417[21:0];
  assign AccumDotWidth_mux1h_1058_nl = MUX1HOT_v_21_3_2((z_out_598_29_7[22:2]), (z_out_1082_29_7[22:2]),
      (z_out_1161_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1059_nl = MUX1HOT_v_21_3_2((z_out_1069_29_7[22:2]),
      (z_out_928_29_7[22:2]), (z_out_1090_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[6])});
  assign nl_z_out_418 = conv_s2u_21_22(AccumDotWidth_mux1h_1058_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1059_nl);
  assign z_out_418 = nl_z_out_418[21:0];
  assign AccumDotWidth_mux1h_1060_nl = MUX1HOT_v_21_3_2((z_out_862_29_7[22:2]), (z_out_1084_29_7[22:2]),
      (z_out_1051_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1061_nl = MUX1HOT_v_21_3_2((z_out_888_29_7[22:2]), (z_out_934_29_7[22:2]),
      (z_out_1101_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])});
  assign nl_z_out_419 = conv_s2u_21_22(AccumDotWidth_mux1h_1060_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1061_nl);
  assign z_out_419 = nl_z_out_419[21:0];
  assign AccumDotWidth_mux_109_nl = MUX_v_21_2_2((z_out_921_29_7[22:2]), (z_out_883_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_110_nl = MUX_v_21_2_2((z_out_1087_29_7[22:2]), (z_out_949_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_420 = conv_s2u_21_22(AccumDotWidth_mux_109_nl) + conv_s2u_21_22(AccumDotWidth_mux_110_nl);
  assign z_out_420 = nl_z_out_420[21:0];
  assign AccumDotWidth_mux_111_nl = MUX_v_21_2_2((z_out_1168_29_7[22:2]), (z_out_971_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_112_nl = MUX_v_21_2_2((z_out_948_29_7[22:2]), (z_out_918_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_421 = conv_s2u_21_22(AccumDotWidth_mux_111_nl) + conv_s2u_21_22(AccumDotWidth_mux_112_nl);
  assign z_out_421 = nl_z_out_421[21:0];
  assign AccumDotWidth_mux1h_1062_nl = MUX1HOT_v_21_4_2((z_out_1041_29_7[22:2]),
      (z_out_997_29_7[22:2]), z_out_963_29_9, (z_out_1002_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1063_nl = MUX1HOT_v_21_4_2((z_out_568_29_7[22:2]), (z_out_1002_29_7[22:2]),
      (z_out_905_29_7[22:2]), (z_out_878_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6])});
  assign nl_z_out_422 = conv_s2u_21_22(AccumDotWidth_mux1h_1062_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1063_nl);
  assign z_out_422 = nl_z_out_422[21:0];
  assign AccumDotWidth_mux1h_1064_nl = MUX1HOT_v_21_4_2((z_out_1053_29_7[22:2]),
      (z_out_1001_29_7[22:2]), (z_out_603_29_7[22:2]), (z_out_1040_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1065_nl = MUX1HOT_v_21_4_2((z_out_946_29_7[22:2]), z_out_1003_29_9,
      z_out_1061_29_9, (z_out_960_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6])});
  assign nl_z_out_423 = conv_s2u_21_22(AccumDotWidth_mux1h_1064_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1065_nl);
  assign z_out_423 = nl_z_out_423[21:0];
  assign AccumDotWidth_mux1h_1066_nl = MUX1HOT_v_21_7_2((z_out_1068_29_7[22:2]),
      (z_out_1176_29_7[22:2]), (z_out_875_29_7[22:2]), z_out_1143_29_9, (z_out_987_29_7[22:2]),
      (z_out_896_29_7[22:2]), (z_out_1131_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1067_nl = MUX1HOT_v_21_7_2((z_out_582_29_7[22:2]), (z_out_1175_29_7[22:2]),
      (z_out_930_29_7[22:2]), (z_out_1016_29_7[22:2]), (z_out_1037_29_7[22:2]), (z_out_615_29_7[22:2]),
      (z_out_1150_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_424 = conv_s2u_21_22(AccumDotWidth_mux1h_1066_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1067_nl);
  assign z_out_424 = nl_z_out_424[21:0];
  assign nl_AccumDotWidth_acc_2492_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2492_nl = nl_AccumDotWidth_acc_2492_nl[9:0];
  assign nl_AccumDotWidth_acc_2493_nl = (nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2493_nl = nl_AccumDotWidth_acc_2493_nl[9:0];
  assign AccumDotWidth_mux_113_nl = MUX_v_10_2_2((AccumDotWidth_acc_2492_nl), (AccumDotWidth_acc_2493_nl),
      fsm_output[3]);
  assign AccumDotWidth_mux_114_nl = MUX_v_11_2_2((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0]),
      (nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm[10:0]),
      fsm_output[3]);
  assign nl_z_out_425 = conv_s2u_21_22({(AccumDotWidth_mux_113_nl) , (AccumDotWidth_mux_114_nl)})
      + conv_s2u_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm);
  assign z_out_425 = nl_z_out_425[21:0];
  assign nl_AccumDotWidth_acc_2494_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2494_nl = nl_AccumDotWidth_acc_2494_nl[9:0];
  assign nl_AccumDotWidth_acc_2495_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2495_nl = nl_AccumDotWidth_acc_2495_nl[9:0];
  assign AccumDotWidth_mux_115_nl = MUX_v_10_2_2((AccumDotWidth_acc_2494_nl), (AccumDotWidth_acc_2495_nl),
      fsm_output[3]);
  assign AccumDotWidth_mux_116_nl = MUX_v_11_2_2((ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0]),
      (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0]),
      fsm_output[3]);
  assign nl_z_out_426 = conv_s2u_21_22({(AccumDotWidth_mux_115_nl) , (AccumDotWidth_mux_116_nl)})
      + conv_s2u_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm);
  assign z_out_426 = nl_z_out_426[21:0];
  assign nl_AccumDotWidth_acc_2496_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2496_nl = nl_AccumDotWidth_acc_2496_nl[9:0];
  assign nl_AccumDotWidth_acc_2497_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2497_nl = nl_AccumDotWidth_acc_2497_nl[9:0];
  assign AccumDotWidth_mux_117_nl = MUX_v_10_2_2((AccumDotWidth_acc_2496_nl), (AccumDotWidth_acc_2497_nl),
      fsm_output[4]);
  assign AccumDotWidth_mux_118_nl = MUX_v_21_2_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      fsm_output[4]);
  assign nl_z_out_427 = conv_s2u_21_22({(AccumDotWidth_mux_117_nl) , (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0])})
      + conv_s2u_21_22(AccumDotWidth_mux_118_nl);
  assign z_out_427 = nl_z_out_427[21:0];
  assign nl_AccumDotWidth_acc_2498_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2498_nl = nl_AccumDotWidth_acc_2498_nl[9:0];
  assign nl_AccumDotWidth_acc_2499_nl = (ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]);
  assign AccumDotWidth_acc_2499_nl = nl_AccumDotWidth_acc_2499_nl[9:0];
  assign nl_AccumDotWidth_acc_2500_nl = (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2500_nl = nl_AccumDotWidth_acc_2500_nl[9:0];
  assign AccumDotWidth_mux1h_1068_nl = MUX1HOT_v_10_3_2((AccumDotWidth_acc_2498_nl),
      (AccumDotWidth_acc_2499_nl), (AccumDotWidth_acc_2500_nl), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign AccumDotWidth_AccumDotWidth_mux_21_nl = MUX_v_11_2_2((ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm[10:0]),
      (ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm[10:0]),
      fsm_output[4]);
  assign nl_z_out_428 = conv_s2u_21_22({(AccumDotWidth_mux1h_1068_nl) , (AccumDotWidth_AccumDotWidth_mux_21_nl)})
      + conv_s2u_21_22(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_slc_29_9_itm);
  assign z_out_428 = nl_z_out_428[21:0];
  assign nl_AccumDotWidth_acc_2501_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2501_nl = nl_AccumDotWidth_acc_2501_nl[9:0];
  assign nl_AccumDotWidth_acc_2502_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2502_nl = nl_AccumDotWidth_acc_2502_nl[9:0];
  assign nl_AccumDotWidth_acc_2503_nl = (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2503_nl = nl_AccumDotWidth_acc_2503_nl[9:0];
  assign AccumDotWidth_mux1h_1069_nl = MUX1HOT_v_10_3_2((AccumDotWidth_acc_2501_nl),
      (AccumDotWidth_acc_2502_nl), (AccumDotWidth_acc_2503_nl), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_429 = conv_s2u_21_22({(AccumDotWidth_mux1h_1069_nl) , (ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm[10:0])})
      + conv_s2u_21_22(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm);
  assign z_out_429 = nl_z_out_429[21:0];
  assign AccumDotWidth_mux1h_1070_nl = MUX1HOT_v_21_3_2((z_out_961_29_7[22:2]), (z_out_1081_29_7[22:2]),
      (z_out_1021_29_7[22:2]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1071_nl = MUX1HOT_v_21_3_2(z_out_1188_29_9, (z_out_909_29_7[22:2]),
      z_out_1046_29_9, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])});
  assign nl_z_out_430 = conv_s2u_21_22(AccumDotWidth_mux1h_1070_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1071_nl);
  assign z_out_430 = nl_z_out_430[21:0];
  assign AccumDotWidth_mux1h_1072_nl = MUX1HOT_v_21_5_2((z_out_968_29_7[22:2]), (z_out_1186_29_7[22:2]),
      (z_out_1129_29_7[22:2]), (z_out_869_29_7[22:2]), (z_out_1121_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1073_nl = MUX1HOT_v_21_5_2((z_out_1008_29_7[22:2]),
      (z_out_1177_29_7[22:2]), (z_out_1011_29_7[22:2]), (z_out_1028_29_7[22:2]),
      z_out_1139_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6])});
  assign nl_z_out_431 = conv_s2u_21_22(AccumDotWidth_mux1h_1072_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1073_nl);
  assign z_out_431 = nl_z_out_431[21:0];
  assign AccumDotWidth_mux_119_nl = MUX_v_21_2_2((z_out_886_29_7[22:2]), (z_out_1099_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_120_nl = MUX_v_21_2_2((z_out_1169_29_7[22:2]), (z_out_902_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_432 = conv_s2u_21_22(AccumDotWidth_mux_119_nl) + conv_s2u_21_22(AccumDotWidth_mux_120_nl);
  assign z_out_432 = nl_z_out_432[21:0];
  assign AccumDotWidth_mux_121_nl = MUX_v_21_2_2((z_out_1162_29_7[22:2]), (z_out_1172_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_122_nl = MUX_v_21_2_2((z_out_1085_29_7[22:2]), (z_out_1180_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_433 = conv_s2u_21_22(AccumDotWidth_mux_121_nl) + conv_s2u_21_22(AccumDotWidth_mux_122_nl);
  assign z_out_433 = nl_z_out_433[21:0];
  assign AccumDotWidth_mux_123_nl = MUX_v_21_2_2((z_out_1146_29_7[22:2]), (z_out_1095_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_124_nl = MUX_v_21_2_2((z_out_586_29_7[22:2]), (z_out_585_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_434 = conv_s2u_21_22(AccumDotWidth_mux_123_nl) + conv_s2u_21_22(AccumDotWidth_mux_124_nl);
  assign z_out_434 = nl_z_out_434[21:0];
  assign AccumDotWidth_mux_125_nl = MUX_v_21_2_2((z_out_973_29_7[22:2]), (z_out_887_29_7[22:2]),
      fsm_output[3]);
  assign AccumDotWidth_mux_126_nl = MUX_v_21_2_2((z_out_1070_29_7[22:2]), (z_out_1101_29_7[22:2]),
      fsm_output[3]);
  assign nl_z_out_435 = conv_s2u_21_22(AccumDotWidth_mux_125_nl) + conv_s2u_21_22(AccumDotWidth_mux_126_nl);
  assign z_out_435 = nl_z_out_435[21:0];
  assign nl_MultLoop_acc_1449_nl = z_out_519 + MultLoop_acc_613_itm;
  assign MultLoop_acc_1449_nl = nl_MultLoop_acc_1449_nl[21:0];
  assign nl_MultLoop_acc_1448_nl = (MultLoop_acc_1449_nl) + MultLoop_acc_629_itm;
  assign MultLoop_acc_1448_nl = nl_MultLoop_acc_1448_nl[21:0];
  assign nl_MultLoop_acc_1447_nl = (MultLoop_acc_1448_nl) + MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1447_nl = nl_MultLoop_acc_1447_nl[21:0];
  assign MultLoop_mux1h_430_nl = MUX1HOT_v_22_4_2(z_out_40_28_7, MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_644_28_7, (MultLoop_acc_1447_nl), {(fsm_output[1]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1450_nl = MultLoop_acc_499_itm + z_out_756;
  assign MultLoop_acc_1450_nl = nl_MultLoop_acc_1450_nl[21:0];
  assign MultLoop_mux1h_431_nl = MUX1HOT_v_22_4_2(z_out_41_28_7, z_out_98_28_7, MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      (MultLoop_acc_1450_nl), {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[8])});
  assign nl_z_out_436 = (MultLoop_mux1h_430_nl) + (MultLoop_mux1h_431_nl);
  assign z_out_436 = nl_z_out_436[21:0];
  assign MultLoop_mux_89_nl = MUX_v_22_2_2(z_out_633_28_7, z_out_66_28_7, fsm_output[3]);
  assign MultLoop_mux_90_nl = MUX_v_22_2_2(MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_63_28_7, fsm_output[3]);
  assign nl_z_out_437 = (MultLoop_mux_89_nl) + (MultLoop_mux_90_nl);
  assign z_out_437 = nl_z_out_437[21:0];
  assign MultLoop_mux1h_432_nl = MUX1HOT_v_22_5_2(z_out_129_28_7, z_out_169_28_7,
      z_out_631_28_7, z_out_131_28_7, z_out_67_28_7, {(fsm_output[1]) , (fsm_output[7])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[5]) , (fsm_output[3])});
  assign MultLoop_mux1h_433_nl = MUX1HOT_v_22_6_2(z_out_130_28_7, z_out_176_28_7,
      z_out_633_28_7, z_out_113_28_7, z_out_132_28_7, z_out_74_28_7, {(fsm_output[1])
      , (fsm_output[7]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[3])});
  assign nl_z_out_438 = (MultLoop_mux1h_432_nl) + (MultLoop_mux1h_433_nl);
  assign z_out_438 = nl_z_out_438[21:0];
  assign MultLoop_mux1h_434_nl = MUX1HOT_v_22_3_2(z_out_641_28_7, z_out_642_28_7,
      z_out_79_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign MultLoop_mux1h_435_nl = MUX1HOT_v_22_3_2(MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_641_28_7, z_out_68_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[3])});
  assign nl_z_out_439 = (MultLoop_mux1h_434_nl) + (MultLoop_mux1h_435_nl);
  assign z_out_439 = nl_z_out_439[21:0];
  assign MultLoop_mux_91_nl = MUX_v_22_2_2(z_out_839, z_out_89_28_7, fsm_output[3]);
  assign MultLoop_mux_92_nl = MUX_v_22_2_2(z_out_832, z_out_78_28_7, fsm_output[3]);
  assign nl_z_out_440 = (MultLoop_mux_91_nl) + (MultLoop_mux_92_nl);
  assign z_out_440 = nl_z_out_440[21:0];
  assign MultLoop_mux1h_436_nl = MUX1HOT_v_22_4_2(z_out_135_28_7, z_out_632_28_7,
      z_out_47_28_7, z_out_650_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign MultLoop_mux1h_437_nl = MUX1HOT_v_22_4_2(z_out_122_28_7, z_out_145_28_7,
      z_out_120_28_7, z_out_189_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_441 = (MultLoop_mux1h_436_nl) + (MultLoop_mux1h_437_nl);
  assign z_out_441 = nl_z_out_441[21:0];
  assign MultLoop_mux1h_438_nl = MUX1HOT_v_22_5_2(z_out_131_28_7, z_out_77_28_7,
      z_out_648_28_7, z_out_132_28_7, z_out_67_28_7, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_439_nl = MUX1HOT_v_22_5_2(z_out_132_28_7, z_out_61_28_7,
      z_out_661_28_7, z_out_131_28_7, z_out_63_28_7, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_442 = (MultLoop_mux1h_438_nl) + (MultLoop_mux1h_439_nl);
  assign z_out_442 = nl_z_out_442[21:0];
  assign MultLoop_mux1h_440_nl = MUX1HOT_v_22_3_2(z_out_49_28_7, MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_632_28_7, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_441_nl = MUX1HOT_v_22_3_2(z_out_36_28_7, z_out_113_28_7,
      MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_443 = (MultLoop_mux1h_440_nl) + (MultLoop_mux1h_441_nl);
  assign z_out_443 = nl_z_out_443[21:0];
  assign AccumDotWidth_mux_127_nl = MUX_v_22_2_2(z_out_818, MultLoop_acc_308_itm,
      fsm_output[8]);
  assign AccumDotWidth_mux_128_nl = MUX_v_22_2_2(z_out_751, z_out_281, fsm_output[8]);
  assign nl_z_out_444 = (AccumDotWidth_mux_127_nl) + (AccumDotWidth_mux_128_nl);
  assign z_out_444 = nl_z_out_444[21:0];
  assign AccumDotWidth_mux_129_nl = MUX_v_22_2_2(z_out_808, z_out_759, fsm_output[8]);
  assign AccumDotWidth_mux_130_nl = MUX_v_22_2_2(z_out_519, z_out_533, fsm_output[8]);
  assign nl_z_out_445 = (AccumDotWidth_mux_129_nl) + (AccumDotWidth_mux_130_nl);
  assign z_out_445 = nl_z_out_445[21:0];
  assign MultLoop_mux1h_442_nl = MUX1HOT_v_22_3_2(z_out_136_28_7, z_out_814, z_out_638_28_7,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_443_nl = MUX1HOT_v_22_3_2(z_out_142_28_7, z_out_817, MultLoop_647_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_446 = (MultLoop_mux1h_442_nl) + (MultLoop_mux1h_443_nl);
  assign z_out_446 = nl_z_out_446[21:0];
  assign MultLoop_mux1h_444_nl = MUX1HOT_v_22_4_2(z_out_169_28_7, z_out_633_28_7,
      z_out_121_28_7, MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_mux1h_445_nl = MUX1HOT_v_22_4_2(MultLoop_1108_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_80_28_7, z_out_124_28_7, z_out_129_28_7, {(fsm_output[4]) , (fsm_output[3])
      , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_447 = (MultLoop_mux1h_444_nl) + (MultLoop_mux1h_445_nl);
  assign z_out_447 = nl_z_out_447[21:0];
  assign MultLoop_MultLoop_mux_14_nl = MUX_v_22_2_2(z_out_820, z_out_84_28_7, fsm_output[3]);
  assign MultLoop_mux1h_446_nl = MUX1HOT_v_22_3_2(z_out_826, z_out_82_28_7, z_out_823,
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_448 = (MultLoop_MultLoop_mux_14_nl) + (MultLoop_mux1h_446_nl);
  assign z_out_448 = nl_z_out_448[21:0];
  assign MultLoop_mux1h_447_nl = MUX1HOT_v_22_3_2(z_out_823, z_out_829, z_out_62_28_7,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign MultLoop_mux1h_448_nl = MUX1HOT_v_22_3_2(z_out_828, z_out_830, z_out_64_28_7,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_z_out_449 = (MultLoop_mux1h_447_nl) + (MultLoop_mux1h_448_nl);
  assign z_out_449 = nl_z_out_449[21:0];
  assign AccumDotWidth_mux1h_1074_nl = MUX1HOT_v_22_5_2(z_out_735, z_out_843, z_out_524,
      z_out_253, z_out_333, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1075_nl = MUX1HOT_v_22_5_2(z_out_731, z_out_841, z_out_516,
      z_out_344, MultLoop_acc_460_itm, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_450 = (AccumDotWidth_mux1h_1074_nl) + (AccumDotWidth_mux1h_1075_nl);
  assign z_out_450 = nl_z_out_450[21:0];
  assign MultLoop_mux1h_449_nl = MUX1HOT_v_22_3_2(z_out_73_28_7, z_out_88_28_7, z_out_137_28_7,
      {MultLoop_or_81_cse , (fsm_output[3]) , (fsm_output[4])});
  assign MultLoop_mux1h_450_nl = MUX1HOT_v_22_4_2(z_out_71_28_7, z_out_638_28_7,
      z_out_133_28_7, z_out_74_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5])});
  assign nl_z_out_451 = (MultLoop_mux1h_449_nl) + (MultLoop_mux1h_450_nl);
  assign z_out_451 = nl_z_out_451[21:0];
  assign MultLoop_mux1h_451_nl = MUX1HOT_v_22_5_2(z_out_70_28_7, z_out_52_28_7, z_out_35_28_7,
      z_out_83_28_7, z_out_79_28_7, {AccumDotWidth_or_132_cse_1 , (fsm_output[2])
      , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_452_nl = MUX1HOT_v_22_5_2(z_out_644_28_7, z_out_53_28_7,
      z_out_75_28_7, MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_639_28_7, {(fsm_output[1]) , (fsm_output[2]) , AccumDotWidth_or_38_cse
      , (fsm_output[7]) , (fsm_output[3])});
  assign nl_z_out_452 = (MultLoop_mux1h_451_nl) + (MultLoop_mux1h_452_nl);
  assign z_out_452 = nl_z_out_452[21:0];
  assign AccumDotWidth_mux1h_1076_nl = MUX1HOT_v_22_8_2(z_out_681, z_out_832, z_out_833,
      z_out_229, z_out_242, z_out_255, z_out_522, z_out_341, {(fsm_output[2]) , (fsm_output[5])
      , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1452_nl = z_out_185_28_7 + z_out_149_28_7;
  assign MultLoop_acc_1452_nl = nl_MultLoop_acc_1452_nl[21:0];
  assign nl_MultLoop_acc_1453_nl = z_out_165_28_7 + z_out_176_28_7;
  assign MultLoop_acc_1453_nl = nl_MultLoop_acc_1453_nl[21:0];
  assign nl_MultLoop_acc_1451_nl = (MultLoop_acc_1452_nl) + (MultLoop_acc_1453_nl);
  assign MultLoop_acc_1451_nl = nl_MultLoop_acc_1451_nl[21:0];
  assign AccumDotWidth_mux1h_1077_nl = MUX1HOT_v_22_7_2(z_out_680, z_out_821, z_out_323,
      z_out_259, z_out_340, z_out_517, (MultLoop_acc_1451_nl), {(fsm_output[2]) ,
      AccumDotWidth_or_38_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_453 = (AccumDotWidth_mux1h_1076_nl) + (AccumDotWidth_mux1h_1077_nl);
  assign z_out_453 = nl_z_out_453[21:0];
  assign nl_AccumDotWidth_acc_2504_nl = z_out_275 + z_out_266;
  assign AccumDotWidth_acc_2504_nl = nl_AccumDotWidth_acc_2504_nl[21:0];
  assign AccumDotWidth_mux1h_1078_nl = MUX1HOT_v_22_5_2(z_out_683, (AccumDotWidth_acc_2504_nl),
      z_out_247, z_out_333, z_out_262, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[671:664]));
  assign MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1871_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[679:672]));
  assign MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1455_nl = (readslicef_29_22_7((MultLoop_84_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_85_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1455_nl = nl_MultLoop_acc_1455_nl[21:0];
  assign nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1877_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[687:680]));
  assign MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(AccumDotWidth_acc_1916_itm[20:0])) * $signed((MultLoop_io_read_w4_rsc_cse_sva[695:688]));
  assign MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1456_nl = (readslicef_29_22_7((MultLoop_86_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_87_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1456_nl = nl_MultLoop_acc_1456_nl[21:0];
  assign nl_MultLoop_acc_1454_nl = (MultLoop_acc_1455_nl) + (MultLoop_acc_1456_nl);
  assign MultLoop_acc_1454_nl = nl_MultLoop_acc_1454_nl[21:0];
  assign AccumDotWidth_mux1h_1079_nl = MUX1HOT_v_22_5_2(z_out_682, z_out_528, z_out_345,
      AccumDotWidth_acc_1845_itm, (MultLoop_acc_1454_nl), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_454 = (AccumDotWidth_mux1h_1078_nl) + (AccumDotWidth_mux1h_1079_nl);
  assign z_out_454 = nl_z_out_454[21:0];
  assign MultLoop_mux1h_453_nl = MUX1HOT_v_22_4_2(z_out_58_28_7, z_out_810, z_out_846,
      z_out_817, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_454_nl = MUX1HOT_v_22_4_2(z_out_57_28_7, z_out_811, z_out_826,
      z_out_814, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_455 = (MultLoop_mux1h_453_nl) + (MultLoop_mux1h_454_nl);
  assign z_out_455 = nl_z_out_455[21:0];
  assign nl_AccumDotWidth_acc_2505_nl = z_out_283 + z_out_274;
  assign AccumDotWidth_acc_2505_nl = nl_AccumDotWidth_acc_2505_nl[21:0];
  assign nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[10047:10040]));
  assign MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[10055:10048]));
  assign MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1458_nl = (readslicef_29_22_7((MultLoop_1256_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1257_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1458_nl = nl_MultLoop_acc_1458_nl[21:0];
  assign nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[10063:10056]));
  assign MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1459_nl = (readslicef_29_22_7((MultLoop_1258_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + MultLoop_1259_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1459_nl = nl_MultLoop_acc_1459_nl[21:0];
  assign nl_MultLoop_acc_1457_nl = (MultLoop_acc_1458_nl) + (MultLoop_acc_1459_nl);
  assign MultLoop_acc_1457_nl = nl_MultLoop_acc_1457_nl[21:0];
  assign AccumDotWidth_mux1h_1080_nl = MUX1HOT_v_22_8_2(z_out_685, z_out_836, z_out_828,
      (AccumDotWidth_acc_2505_nl), z_out_526, z_out_254, z_out_332, (MultLoop_acc_1457_nl),
      {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1081_nl = MUX1HOT_v_22_8_2(z_out_686, z_out_842, z_out_836,
      z_out_516, z_out_529, z_out_349, z_out_526, MultLoop_acc_1095_itm, {(fsm_output[2])
      , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_456 = (AccumDotWidth_mux1h_1080_nl) + (AccumDotWidth_mux1h_1081_nl);
  assign z_out_456 = nl_z_out_456[21:0];
  assign nl_MultLoop_acc_1462_nl = z_out_518 + MultLoop_acc_597_itm;
  assign MultLoop_acc_1462_nl = nl_MultLoop_acc_1462_nl[21:0];
  assign nl_MultLoop_acc_1465_nl = (z_out_1064_29_7[21:0]) + (z_out_1045_29_7[21:0]);
  assign MultLoop_acc_1465_nl = nl_MultLoop_acc_1465_nl[21:0];
  assign nl_MultLoop_acc_1466_nl = (z_out_909_29_7[21:0]) + (z_out_916_29_7[21:0]);
  assign MultLoop_acc_1466_nl = nl_MultLoop_acc_1466_nl[21:0];
  assign nl_MultLoop_acc_1461_nl = (MultLoop_acc_1462_nl) + MultLoop_acc_596_itm
      + (MultLoop_acc_1465_nl) + (MultLoop_acc_1466_nl);
  assign MultLoop_acc_1461_nl = nl_MultLoop_acc_1461_nl[21:0];
  assign nl_MultLoop_acc_1460_nl = (MultLoop_acc_1461_nl) + z_out_752;
  assign MultLoop_acc_1460_nl = nl_MultLoop_acc_1460_nl[21:0];
  assign MultLoop_mux1h_455_nl = MUX1HOT_v_22_6_2(z_out_62_28_7, z_out_54_28_7, MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_640_28_7, z_out_100_28_7, (MultLoop_acc_1460_nl), {MultLoop_or_81_cse
      , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1467_nl = z_out_751 + MultLoop_acc_631_itm;
  assign MultLoop_acc_1467_nl = nl_MultLoop_acc_1467_nl[21:0];
  assign MultLoop_mux1h_456_nl = MUX1HOT_v_22_7_2(z_out_653_28_7, z_out_111_28_7,
      z_out_36_28_7, z_out_661_28_7, z_out_74_28_7, z_out_61_28_7, (MultLoop_acc_1467_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_457 = (MultLoop_mux1h_455_nl) + (MultLoop_mux1h_456_nl);
  assign z_out_457 = nl_z_out_457[21:0];
  assign nl_AccumDotWidth_acc_2506_nl = z_out_703 + z_out_707;
  assign AccumDotWidth_acc_2506_nl = nl_AccumDotWidth_acc_2506_nl[21:0];
  assign nl_MultLoop_acc_1468_nl = z_out_548 + z_out_550;
  assign MultLoop_acc_1468_nl = nl_MultLoop_acc_1468_nl[21:0];
  assign AccumDotWidth_mux1h_1082_nl = MUX1HOT_v_22_4_2(z_out_345, (AccumDotWidth_acc_2506_nl),
      z_out_260, (MultLoop_acc_1468_nl), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2507_nl = z_out_709 + z_out_705;
  assign AccumDotWidth_acc_2507_nl = nl_AccumDotWidth_acc_2507_nl[21:0];
  assign AccumDotWidth_mux1h_1083_nl = MUX1HOT_v_22_4_2(z_out_732, (AccumDotWidth_acc_2507_nl),
      z_out_342, z_out_527, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_458 = (AccumDotWidth_mux1h_1082_nl) + (AccumDotWidth_mux1h_1083_nl);
  assign z_out_458 = nl_z_out_458[21:0];
  assign MultLoop_mux1h_457_nl = MUX1HOT_v_22_3_2(z_out_833, z_out_319, z_out_334,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[8])});
  assign MultLoop_mux1h_458_nl = MUX1HOT_v_22_3_2(z_out_834, z_out_517, z_out_330,
      {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[8])});
  assign nl_z_out_459 = (MultLoop_mux1h_457_nl) + (MultLoop_mux1h_458_nl);
  assign z_out_459 = nl_z_out_459[21:0];
  assign nl_MultLoop_acc_1470_nl = z_out_148_28_7 + z_out_147_28_7;
  assign MultLoop_acc_1470_nl = nl_MultLoop_acc_1470_nl[21:0];
  assign nl_MultLoop_acc_1471_nl = z_out_146_28_7 + MultLoop_107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1471_nl = nl_MultLoop_acc_1471_nl[21:0];
  assign nl_MultLoop_acc_1469_nl = (MultLoop_acc_1470_nl) + (MultLoop_acc_1471_nl);
  assign MultLoop_acc_1469_nl = nl_MultLoop_acc_1469_nl[21:0];
  assign MultLoop_mux_93_nl = MUX_v_22_2_2(z_out_498, (MultLoop_acc_1469_nl), fsm_output[8]);
  assign MultLoop_mux_94_nl = MUX_v_22_2_2(z_out_499, MultLoop_acc_1222_itm, fsm_output[8]);
  assign nl_z_out_460 = (MultLoop_mux_93_nl) + (MultLoop_mux_94_nl);
  assign z_out_460 = nl_z_out_460[21:0];
  assign nl_AccumDotWidth_acc_2508_nl = conv_s2s_21_22(z_out_1010_29_7[22:2]) + conv_s2s_21_22(z_out_874_29_7[22:2]);
  assign AccumDotWidth_acc_2508_nl = nl_AccumDotWidth_acc_2508_nl[21:0];
  assign AccumDotWidth_mux1h_1084_nl = MUX1HOT_v_22_4_2(z_out_388, (AccumDotWidth_acc_2508_nl),
      z_out_380, (z_out_600_29_7[21:0]), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2509_nl = conv_s2s_21_22(z_out_880_29_7[22:2]) + conv_s2s_21_22(z_out_1100_29_7[22:2]);
  assign AccumDotWidth_acc_2509_nl = nl_AccumDotWidth_acc_2509_nl[21:0];
  assign AccumDotWidth_mux1h_1085_nl = MUX1HOT_v_22_4_2(z_out_392, (AccumDotWidth_acc_2509_nl),
      z_out_375, (z_out_1113_29_7[21:0]), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_461 = (AccumDotWidth_mux1h_1084_nl) + (AccumDotWidth_mux1h_1085_nl);
  assign z_out_461 = nl_z_out_461[21:0];
  assign AccumDotWidth_mux_131_nl = MUX_v_22_2_2(z_out_397, (z_out_595_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_132_nl = MUX_v_22_2_2(z_out_386, (z_out_596_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_462 = (AccumDotWidth_mux_131_nl) + (AccumDotWidth_mux_132_nl);
  assign z_out_462 = nl_z_out_462[21:0];
  assign nl_AccumDotWidth_acc_2510_nl = conv_s2s_21_22(z_out_987_29_7[22:2]) + conv_s2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm);
  assign AccumDotWidth_acc_2510_nl = nl_AccumDotWidth_acc_2510_nl[21:0];
  assign AccumDotWidth_mux1h_1086_nl = MUX1HOT_v_22_3_2((AccumDotWidth_acc_2510_nl),
      z_out_252, z_out_339, {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1472_nl = z_out_525 + z_out_544;
  assign MultLoop_acc_1472_nl = nl_MultLoop_acc_1472_nl[21:0];
  assign AccumDotWidth_mux1h_1087_nl = MUX1HOT_v_22_3_2(AccumDotWidth_acc_1916_itm,
      z_out_250, (MultLoop_acc_1472_nl), {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_463 = (AccumDotWidth_mux1h_1086_nl) + (AccumDotWidth_mux1h_1087_nl);
  assign z_out_463 = nl_z_out_463[21:0];
  assign nl_MultLoop_acc_1474_nl = z_out_674_28_7 + z_out_675_28_7;
  assign MultLoop_acc_1474_nl = nl_MultLoop_acc_1474_nl[21:0];
  assign nl_MultLoop_acc_1473_nl = z_out_492 + (MultLoop_acc_1474_nl);
  assign MultLoop_acc_1473_nl = nl_MultLoop_acc_1473_nl[21:0];
  assign AccumDotWidth_mux1h_1088_nl = MUX1HOT_v_22_4_2(z_out_394, z_out_333, z_out_257,
      (MultLoop_acc_1473_nl), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1476_nl = (z_out_623_29_7[21:0]) + z_out_160_28_7;
  assign MultLoop_acc_1476_nl = nl_MultLoop_acc_1476_nl[21:0];
  assign nl_MultLoop_acc_1477_nl = z_out_161_28_7 + z_out_162_28_7;
  assign MultLoop_acc_1477_nl = nl_MultLoop_acc_1477_nl[21:0];
  assign nl_MultLoop_acc_1475_nl = (MultLoop_acc_1476_nl) + (MultLoop_acc_1477_nl);
  assign MultLoop_acc_1475_nl = nl_MultLoop_acc_1475_nl[21:0];
  assign AccumDotWidth_mux1h_1089_nl = MUX1HOT_v_22_4_2(z_out_390, z_out_323, z_out_261,
      (MultLoop_acc_1475_nl), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_464 = (AccumDotWidth_mux1h_1088_nl) + (AccumDotWidth_mux1h_1089_nl);
  assign z_out_464 = nl_z_out_464[21:0];
  assign MultLoop_mux1h_459_nl = MUX1HOT_v_22_4_2(z_out_635_28_7, z_out_122_28_7,
      z_out_61_28_7, z_out_71_28_7, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5])});
  assign MultLoop_mux1h_460_nl = MUX1HOT_v_22_4_2(z_out_653_28_7, z_out_54_28_7,
      z_out_82_28_7, z_out_72_28_7, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[5])});
  assign nl_z_out_465 = (MultLoop_mux1h_459_nl) + (MultLoop_mux1h_460_nl);
  assign z_out_465 = nl_z_out_465[21:0];
  assign AccumDotWidth_mux1h_1090_nl = MUX1HOT_v_22_8_2(z_out_431, z_out_386, z_out_317,
      z_out_263, z_out_519, z_out_269, z_out_566, z_out_264, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1091_nl = MUX1HOT_v_22_7_2(z_out_422, z_out_388, z_out_523,
      z_out_264, z_out_508, z_out_270, z_out_450, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_466 = (AccumDotWidth_mux1h_1090_nl) + (AccumDotWidth_mux1h_1091_nl);
  assign z_out_466 = nl_z_out_466[21:0];
  assign nl_AccumDotWidth_acc_2511_nl = z_out_685 + z_out_681;
  assign AccumDotWidth_acc_2511_nl = nl_AccumDotWidth_acc_2511_nl[21:0];
  assign AccumDotWidth_mux1h_1092_nl = MUX1HOT_v_22_5_2(z_out_684, z_out_562, z_out_563,
      (AccumDotWidth_acc_2511_nl), z_out_845, {(fsm_output[1]) , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1093_nl = MUX1HOT_v_22_6_2(z_out_682, z_out_523, z_out_517,
      z_out_335, z_out_329, z_out_834, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_467 = (AccumDotWidth_mux1h_1092_nl) + (AccumDotWidth_mux1h_1093_nl);
  assign z_out_467 = nl_z_out_467[21:0];
  assign MultLoop_mux1h_461_nl = MUX1HOT_v_22_5_2(z_out_655_28_7, z_out_42_28_7,
      z_out_108_28_7, z_out_46_28_7, z_out_77_28_7, {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_462_nl = MUX1HOT_v_22_5_2(z_out_642_28_7, z_out_50_28_7,
      z_out_113_28_7, z_out_72_28_7, z_out_135_28_7, {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_468 = (MultLoop_mux1h_461_nl) + (MultLoop_mux1h_462_nl);
  assign z_out_468 = nl_z_out_468[21:0];
  assign nl_MultLoop_acc_1480_nl = (z_out_1176_29_7[21:0]) + (z_out_1175_29_7[21:0]);
  assign MultLoop_acc_1480_nl = nl_MultLoop_acc_1480_nl[21:0];
  assign nl_MultLoop_acc_1481_nl = (z_out_1178_29_7[21:0]) + (z_out_1179_29_7[21:0]);
  assign MultLoop_acc_1481_nl = nl_MultLoop_acc_1481_nl[21:0];
  assign nl_MultLoop_acc_1483_nl = (z_out_1180_29_7[21:0]) + (z_out_994_29_7[21:0]);
  assign MultLoop_acc_1483_nl = nl_MultLoop_acc_1483_nl[21:0];
  assign nl_MultLoop_acc_1484_nl = (z_out_997_29_7[21:0]) + (z_out_1000_29_7[21:0]);
  assign MultLoop_acc_1484_nl = nl_MultLoop_acc_1484_nl[21:0];
  assign nl_MultLoop_acc_1478_nl = (MultLoop_acc_1480_nl) + (MultLoop_acc_1481_nl)
      + (MultLoop_acc_1483_nl) + (MultLoop_acc_1484_nl);
  assign MultLoop_acc_1478_nl = nl_MultLoop_acc_1478_nl[21:0];
  assign AccumDotWidth_mux1h_1094_nl = MUX1HOT_v_22_6_2(z_out_355, z_out_693, z_out_562,
      z_out_566, z_out_556, (MultLoop_acc_1478_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1487_nl = (z_out_1002_29_7[21:0]) + (z_out_999_29_7[21:0]);
  assign MultLoop_acc_1487_nl = nl_MultLoop_acc_1487_nl[21:0];
  assign nl_MultLoop_acc_1486_nl = z_out_849 + (MultLoop_acc_1487_nl);
  assign MultLoop_acc_1486_nl = nl_MultLoop_acc_1486_nl[21:0];
  assign nl_MultLoop_acc_1485_nl = (MultLoop_acc_1486_nl) + z_out_331;
  assign MultLoop_acc_1485_nl = nl_MultLoop_acc_1485_nl[21:0];
  assign AccumDotWidth_mux1h_1095_nl = MUX1HOT_v_22_6_2(z_out_362, z_out_340, z_out_528,
      z_out_333, z_out_551, (MultLoop_acc_1485_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_469 = (AccumDotWidth_mux1h_1094_nl) + (AccumDotWidth_mux1h_1095_nl);
  assign z_out_469 = nl_z_out_469[21:0];
  assign AccumDotWidth_mux1h_1096_nl = MUX1HOT_v_22_3_2(z_out_387, z_out_539, z_out_267,
      {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1097_nl = MUX1HOT_v_22_3_2(z_out_381, z_out_513, z_out_266,
      {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_470 = (AccumDotWidth_mux1h_1096_nl) + (AccumDotWidth_mux1h_1097_nl);
  assign z_out_470 = nl_z_out_470[21:0];
  assign AccumDotWidth_mux1h_1098_nl = MUX1HOT_v_22_6_2(z_out_724, z_out_350, z_out_458,
      z_out_565, z_out_566, z_out_265, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1099_nl = MUX1HOT_v_22_5_2(z_out_359, z_out_339, z_out_543,
      z_out_564, MultLoop_acc_502_itm, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , AccumDotWidth_or_145_cse , (fsm_output[8])});
  assign nl_z_out_471 = (AccumDotWidth_mux1h_1098_nl) + (AccumDotWidth_mux1h_1099_nl);
  assign z_out_471 = nl_z_out_471[21:0];
  assign nl_MultLoop_acc_1490_nl = (z_out_1029_29_7[21:0]) + (z_out_932_29_7[21:0]);
  assign MultLoop_acc_1490_nl = nl_MultLoop_acc_1490_nl[21:0];
  assign nl_MultLoop_acc_1491_nl = (z_out_933_29_7[21:0]) + (z_out_1030_29_7[21:0]);
  assign MultLoop_acc_1491_nl = nl_MultLoop_acc_1491_nl[21:0];
  assign nl_MultLoop_acc_1493_nl = (z_out_1028_29_7[21:0]) + (z_out_1026_29_7[21:0]);
  assign MultLoop_acc_1493_nl = nl_MultLoop_acc_1493_nl[21:0];
  assign nl_MultLoop_acc_1494_nl = (z_out_1025_29_7[21:0]) + (z_out_1024_29_7[21:0]);
  assign MultLoop_acc_1494_nl = nl_MultLoop_acc_1494_nl[21:0];
  assign nl_MultLoop_acc_1488_nl = (MultLoop_acc_1490_nl) + (MultLoop_acc_1491_nl)
      + (MultLoop_acc_1493_nl) + (MultLoop_acc_1494_nl);
  assign MultLoop_acc_1488_nl = nl_MultLoop_acc_1488_nl[21:0];
  assign AccumDotWidth_mux1h_1100_nl = MUX1HOT_v_22_7_2(z_out_393, z_out_744, z_out_318,
      z_out_265, z_out_564, z_out_842, (MultLoop_acc_1488_nl), {(fsm_output[1]) ,
      (fsm_output[2]) , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1497_nl = (z_out_1023_29_7[21:0]) + (z_out_1022_29_7[21:0]);
  assign MultLoop_acc_1497_nl = nl_MultLoop_acc_1497_nl[21:0];
  assign nl_MultLoop_acc_1498_nl = (z_out_950_29_7[21:0]) + (z_out_938_29_7[21:0]);
  assign MultLoop_acc_1498_nl = nl_MultLoop_acc_1498_nl[21:0];
  assign nl_MultLoop_acc_1500_nl = (z_out_951_29_7[21:0]) + (z_out_964_29_7[21:0]);
  assign MultLoop_acc_1500_nl = nl_MultLoop_acc_1500_nl[21:0];
  assign nl_MultLoop_acc_1501_nl = (z_out_990_29_7[21:0]) + (z_out_1174_29_7[21:0]);
  assign MultLoop_acc_1501_nl = nl_MultLoop_acc_1501_nl[21:0];
  assign nl_MultLoop_acc_1495_nl = (MultLoop_acc_1497_nl) + (MultLoop_acc_1498_nl)
      + (MultLoop_acc_1500_nl) + (MultLoop_acc_1501_nl);
  assign MultLoop_acc_1495_nl = nl_MultLoop_acc_1495_nl[21:0];
  assign AccumDotWidth_mux1h_1101_nl = MUX1HOT_v_22_8_2(z_out_389, z_out_750, z_out_508,
      z_out_559, z_out_541, z_out_333, z_out_235, (MultLoop_acc_1495_nl), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_472 = (AccumDotWidth_mux1h_1100_nl) + (AccumDotWidth_mux1h_1101_nl);
  assign z_out_472 = nl_z_out_472[21:0];
  assign nl_MultLoop_acc_1502_nl = z_out_321 + z_out_322;
  assign MultLoop_acc_1502_nl = nl_MultLoop_acc_1502_nl[21:0];
  assign AccumDotWidth_mux1h_1102_nl = MUX1HOT_v_22_3_2(z_out_383, z_out_844, (MultLoop_acc_1502_nl),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1505_nl = (z_out_1094_29_7[21:0]) + (z_out_1008_29_7[21:0]);
  assign MultLoop_acc_1505_nl = nl_MultLoop_acc_1505_nl[21:0];
  assign nl_MultLoop_acc_1504_nl = (MultLoop_acc_1505_nl) + z_out_802;
  assign MultLoop_acc_1504_nl = nl_MultLoop_acc_1504_nl[21:0];
  assign nl_MultLoop_acc_1503_nl = z_out_323 + (MultLoop_acc_1504_nl);
  assign MultLoop_acc_1503_nl = nl_MultLoop_acc_1503_nl[21:0];
  assign AccumDotWidth_mux1h_1103_nl = MUX1HOT_v_22_3_2(z_out_385, z_out_332, (MultLoop_acc_1503_nl),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_473 = (AccumDotWidth_mux1h_1102_nl) + (AccumDotWidth_mux1h_1103_nl);
  assign z_out_473 = nl_z_out_473[21:0];
  assign nl_MultLoop_acc_1508_nl = (z_out_1042_29_7[21:0]) + (z_out_1038_29_7[21:0]);
  assign MultLoop_acc_1508_nl = nl_MultLoop_acc_1508_nl[21:0];
  assign nl_MultLoop_acc_1507_nl = (MultLoop_acc_1508_nl) + z_out_235;
  assign MultLoop_acc_1507_nl = nl_MultLoop_acc_1507_nl[21:0];
  assign nl_MultLoop_acc_1506_nl = (MultLoop_acc_1507_nl) + z_out_508;
  assign MultLoop_acc_1506_nl = nl_MultLoop_acc_1506_nl[21:0];
  assign AccumDotWidth_mux1h_1104_nl = MUX1HOT_v_22_6_2(z_out_385, z_out_341, z_out_350,
      z_out_319, z_out_229, (MultLoop_acc_1506_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[6]) , MultLoop_or_22_cse , (fsm_output[5]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1105_nl = MUX1HOT_v_22_7_2(z_out_681, z_out_347, z_out_339,
      z_out_522, z_out_563, z_out_229, z_out_842, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[6]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_474 = (AccumDotWidth_mux1h_1104_nl) + (AccumDotWidth_mux1h_1105_nl);
  assign z_out_474 = nl_z_out_474[21:0];
  assign AccumDotWidth_mux1h_1106_nl = MUX1HOT_v_22_6_2(z_out_434, z_out_464, z_out_565,
      z_out_816, z_out_325, z_out_270, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1107_nl = MUX1HOT_v_22_6_2(z_out_421, z_out_541, z_out_512,
      AccumDotWidth_acc_1135_itm, z_out_237, z_out_531, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_475 = (AccumDotWidth_mux1h_1106_nl) + (AccumDotWidth_mux1h_1107_nl);
  assign z_out_475 = nl_z_out_475[21:0];
  assign AccumDotWidth_mux1h_1108_nl = MUX1HOT_v_22_5_2(z_out_698, z_out_325, z_out_566,
      z_out_811, z_out_816, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1509_nl = z_out_326 + MultLoop_acc_841_itm;
  assign MultLoop_acc_1509_nl = nl_MultLoop_acc_1509_nl[21:0];
  assign AccumDotWidth_mux1h_1109_nl = MUX1HOT_v_22_5_2(z_out_692, z_out_238, z_out_515,
      z_out_467, (MultLoop_acc_1509_nl), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_476 = (AccumDotWidth_mux1h_1108_nl) + (AccumDotWidth_mux1h_1109_nl);
  assign z_out_476 = nl_z_out_476[21:0];
  assign MultLoop_mux1h_463_nl = MUX1HOT_v_22_4_2(z_out_89_28_7, z_out_647_28_7,
      z_out_118_28_7, z_out_86_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign MultLoop_mux1h_464_nl = MUX1HOT_v_22_4_2(z_out_79_28_7, z_out_648_28_7,
      z_out_142_28_7, z_out_88_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_477 = (MultLoop_mux1h_463_nl) + (MultLoop_mux1h_464_nl);
  assign z_out_477 = nl_z_out_477[21:0];
  assign MultLoop_mux1h_465_nl = MUX1HOT_v_22_4_2(z_out_55_28_7, z_out_637_28_7,
      z_out_125_28_7, z_out_97_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign MultLoop_mux1h_466_nl = MUX1HOT_v_22_4_2(z_out_59_28_7, z_out_636_28_7,
      z_out_124_28_7, z_out_85_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_478 = (MultLoop_mux1h_465_nl) + (MultLoop_mux1h_466_nl);
  assign z_out_478 = nl_z_out_478[21:0];
  assign MultLoop_mux1h_467_nl = MUX1HOT_v_22_4_2(z_out_115_28_7, z_out_35_28_7,
      z_out_657_28_7, z_out_138_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5])});
  assign MultLoop_mux1h_468_nl = MUX1HOT_v_22_4_2(z_out_81_28_7, z_out_34_28_7, z_out_663_28_7,
      z_out_139_28_7, {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_479 = (MultLoop_mux1h_467_nl) + (MultLoop_mux1h_468_nl);
  assign z_out_479 = nl_z_out_479[21:0];
  assign nl_MultLoop_acc_1510_nl = z_out_318 + z_out_317;
  assign MultLoop_acc_1510_nl = nl_MultLoop_acc_1510_nl[21:0];
  assign AccumDotWidth_mux_133_nl = MUX_v_22_2_2(z_out_815, (MultLoop_acc_1510_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1511_nl = z_out_319 + MultLoop_acc_79_itm;
  assign MultLoop_acc_1511_nl = nl_MultLoop_acc_1511_nl[21:0];
  assign AccumDotWidth_mux_134_nl = MUX_v_22_2_2(z_out_469, (MultLoop_acc_1511_nl),
      fsm_output[8]);
  assign nl_z_out_480 = (AccumDotWidth_mux_133_nl) + (AccumDotWidth_mux_134_nl);
  assign z_out_480 = nl_z_out_480[21:0];
  assign AccumDotWidth_mux1h_1110_nl = MUX1HOT_v_22_3_2(z_out_690, z_out_565, z_out_833,
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1514_nl = (z_out_586_29_7[21:0]) + (z_out_587_29_7[21:0]);
  assign MultLoop_acc_1514_nl = nl_MultLoop_acc_1514_nl[21:0];
  assign nl_MultLoop_acc_1513_nl = (MultLoop_acc_1514_nl) + z_out_310;
  assign MultLoop_acc_1513_nl = nl_MultLoop_acc_1513_nl[21:0];
  assign nl_MultLoop_acc_1515_nl = z_out_311 + z_out_315;
  assign MultLoop_acc_1515_nl = nl_MultLoop_acc_1515_nl[21:0];
  assign nl_MultLoop_acc_1512_nl = (MultLoop_acc_1513_nl) + (MultLoop_acc_1515_nl);
  assign MultLoop_acc_1512_nl = nl_MultLoop_acc_1512_nl[21:0];
  assign AccumDotWidth_mux1h_1111_nl = MUX1HOT_v_22_3_2(z_out_699, z_out_562, (MultLoop_acc_1512_nl),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_481 = (AccumDotWidth_mux1h_1110_nl) + (AccumDotWidth_mux1h_1111_nl);
  assign z_out_481 = nl_z_out_481[21:0];
  assign nl_MultLoop_acc_1516_nl = z_out_755 + z_out_823;
  assign MultLoop_acc_1516_nl = nl_MultLoop_acc_1516_nl[21:0];
  assign MultLoop_mux1h_469_nl = MUX1HOT_v_22_3_2(z_out_78_28_7, z_out_62_28_7, (MultLoop_acc_1516_nl),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1519_nl = z_out_340 + z_out_338;
  assign MultLoop_acc_1519_nl = nl_MultLoop_acc_1519_nl[21:0];
  assign nl_MultLoop_acc_1520_nl = z_out_336 + z_out_335;
  assign MultLoop_acc_1520_nl = nl_MultLoop_acc_1520_nl[21:0];
  assign nl_MultLoop_acc_1518_nl = (MultLoop_acc_1519_nl) + (MultLoop_acc_1520_nl);
  assign MultLoop_acc_1518_nl = nl_MultLoop_acc_1518_nl[21:0];
  assign nl_MultLoop_acc_1517_nl = z_out_542 + (MultLoop_acc_1518_nl);
  assign MultLoop_acc_1517_nl = nl_MultLoop_acc_1517_nl[21:0];
  assign MultLoop_mux1h_470_nl = MUX1HOT_v_22_3_2(z_out_64_28_7, z_out_89_28_7, (MultLoop_acc_1517_nl),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_482 = (MultLoop_mux1h_469_nl) + (MultLoop_mux1h_470_nl);
  assign z_out_482 = nl_z_out_482[21:0];
  assign nl_AccumDotWidth_acc_2512_nl = conv_s2s_21_22(z_out_1116_29_7[22:2]) + conv_s2s_21_22(z_out_1048_29_9);
  assign AccumDotWidth_acc_2512_nl = nl_AccumDotWidth_acc_2512_nl[21:0];
  assign AccumDotWidth_mux1h_1112_nl = MUX1HOT_v_22_3_2(z_out_689, (AccumDotWidth_acc_2512_nl),
      (z_out_597_29_7[21:0]), {(fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1113_nl = MUX1HOT_v_22_3_2(z_out_735, z_out_395, (z_out_599_29_7[21:0]),
      {(fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_483 = (AccumDotWidth_mux1h_1112_nl) + (AccumDotWidth_mux1h_1113_nl);
  assign z_out_483 = nl_z_out_483[21:0];
  assign nl_AccumDotWidth_acc_2513_nl = conv_s2s_21_22(z_out_1091_29_7[22:2]) + conv_s2s_21_22(z_out_861_29_7[22:2]);
  assign AccumDotWidth_acc_2513_nl = nl_AccumDotWidth_acc_2513_nl[21:0];
  assign AccumDotWidth_mux1h_1114_nl = MUX1HOT_v_22_5_2(z_out_682, z_out_696, (AccumDotWidth_acc_2513_nl),
      z_out_389, (z_out_1116_29_7[21:0]), {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2514_nl = conv_s2s_21_22(z_out_999_29_7[22:2]) + conv_s2s_21_22(z_out_862_29_7[22:2]);
  assign AccumDotWidth_acc_2514_nl = nl_AccumDotWidth_acc_2514_nl[21:0];
  assign AccumDotWidth_mux1h_1115_nl = MUX1HOT_v_22_5_2(z_out_680, z_out_695, (AccumDotWidth_acc_2514_nl),
      z_out_390, (z_out_1117_29_7[21:0]), {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_484 = (AccumDotWidth_mux1h_1114_nl) + (AccumDotWidth_mux1h_1115_nl);
  assign z_out_484 = nl_z_out_484[21:0];
  assign MultLoop_mux1h_471_nl = MUX1HOT_v_22_4_2(z_out_51_28_7, z_out_81_28_7, z_out_82_28_7,
      z_out_812, {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1521_nl = MultLoop_acc_626_itm + z_out_278;
  assign MultLoop_acc_1521_nl = nl_MultLoop_acc_1521_nl[21:0];
  assign MultLoop_mux1h_472_nl = MUX1HOT_v_22_4_2(z_out_56_28_7, z_out_83_28_7, z_out_61_28_7,
      (MultLoop_acc_1521_nl), {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[8])});
  assign nl_z_out_485 = (MultLoop_mux1h_471_nl) + (MultLoop_mux1h_472_nl);
  assign z_out_485 = nl_z_out_485[21:0];
  assign AccumDotWidth_mux_135_nl = MUX_v_22_2_2(MultLoop_acc_215_itm, (z_out_895_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_136_nl = MUX_v_22_2_2(z_out_331, (z_out_894_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_486 = (AccumDotWidth_mux_135_nl) + (AccumDotWidth_mux_136_nl);
  assign z_out_486 = nl_z_out_486[21:0];
  assign AccumDotWidth_mux_137_nl = MUX_v_22_2_2(MultLoop_acc_356_itm, (z_out_897_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_138_nl = MUX_v_22_2_2(z_out_328, (z_out_896_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_487 = (AccumDotWidth_mux_137_nl) + (AccumDotWidth_mux_138_nl);
  assign z_out_487 = nl_z_out_487[21:0];
  assign nl_AccumDotWidth_acc_2515_nl = conv_s2s_21_22(z_out_625_29_7[22:2]) + conv_s2s_21_22(z_out_895_29_7[22:2]);
  assign AccumDotWidth_acc_2515_nl = nl_AccumDotWidth_acc_2515_nl[21:0];
  assign MultLoop_mux1h_473_nl = MUX1HOT_v_22_6_2(z_out_150_28_7, z_out_670_28_7,
      z_out_404, z_out_385, (AccumDotWidth_acc_2515_nl), (z_out_899_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign MultLoop_mux1h_474_nl = MUX1HOT_v_22_6_2(z_out_158_28_7, z_out_671_28_7,
      z_out_403, z_out_387, z_out_391, (z_out_898_29_7[21:0]), {(fsm_output[6]) ,
      (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_488 = (MultLoop_mux1h_473_nl) + (MultLoop_mux1h_474_nl);
  assign z_out_488 = nl_z_out_488[21:0];
  assign nl_AccumDotWidth_acc_2516_nl = conv_s2s_21_22(z_out_611_29_7[22:2]) + conv_s2s_21_22(z_out_605_29_7[22:2]);
  assign AccumDotWidth_acc_2516_nl = nl_AccumDotWidth_acc_2516_nl[21:0];
  assign AccumDotWidth_mux1h_1116_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2516_nl),
      z_out_407, z_out_406, z_out_375, z_out_396, (z_out_1123_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2517_nl = conv_s2s_21_22(z_out_608_29_7[22:2]) + conv_s2s_21_22(z_out_610_29_7[22:2]);
  assign AccumDotWidth_acc_2517_nl = nl_AccumDotWidth_acc_2517_nl[21:0];
  assign nl_AccumDotWidth_acc_2518_nl = conv_s2s_21_22(z_out_950_29_7[22:2]) + conv_s2s_21_22(z_out_1144_29_9);
  assign AccumDotWidth_acc_2518_nl = nl_AccumDotWidth_acc_2518_nl[21:0];
  assign AccumDotWidth_mux1h_1117_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2517_nl),
      z_out_403, z_out_407, z_out_355, (AccumDotWidth_acc_2518_nl), (z_out_1112_29_7[21:0]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_489 = (AccumDotWidth_mux1h_1116_nl) + (AccumDotWidth_mux1h_1117_nl);
  assign z_out_489 = nl_z_out_489[21:0];
  assign nl_AccumDotWidth_acc_2519_nl = conv_s2s_21_22(z_out_991_29_7[22:2]) + conv_s2s_21_22(z_out_1118_29_7[22:2]);
  assign AccumDotWidth_acc_2519_nl = nl_AccumDotWidth_acc_2519_nl[21:0];
  assign nl_AccumDotWidth_acc_2520_nl = conv_s2s_21_22(z_out_623_29_7[22:2]) + conv_s2s_21_22(z_out_894_29_7[22:2]);
  assign AccumDotWidth_acc_2520_nl = nl_AccumDotWidth_acc_2520_nl[21:0];
  assign MultLoop_mux1h_475_nl = MUX1HOT_v_22_6_2(z_out_161_28_7, z_out_176_28_7,
      z_out_384, (AccumDotWidth_acc_2519_nl), (AccumDotWidth_acc_2520_nl), (z_out_878_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2521_nl = conv_s2s_21_22(z_out_583_29_7[22:2]) + conv_s2s_21_22(z_out_617_29_7[22:2]);
  assign AccumDotWidth_acc_2521_nl = nl_AccumDotWidth_acc_2521_nl[21:0];
  assign MultLoop_mux1h_476_nl = MUX1HOT_v_22_6_2(z_out_162_28_7, z_out_160_28_7,
      z_out_405, z_out_378, (AccumDotWidth_acc_2521_nl), (z_out_877_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_490 = (MultLoop_mux1h_475_nl) + (MultLoop_mux1h_476_nl);
  assign z_out_490 = nl_z_out_490[21:0];
  assign nl_AccumDotWidth_acc_2522_nl = conv_s2s_21_22(z_out_628_29_7[22:2]) + conv_s2s_21_22(z_out_1120_29_7[22:2]);
  assign AccumDotWidth_acc_2522_nl = nl_AccumDotWidth_acc_2522_nl[21:0];
  assign MultLoop_mux1h_477_nl = MUX1HOT_v_22_8_2(z_out_670_28_7, z_out_167_28_7,
      z_out_396, MultLoop_acc_102_itm, z_out_402, z_out_376, (AccumDotWidth_acc_2522_nl),
      (z_out_1111_29_7[21:0]), {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2523_nl = conv_s2s_21_22(z_out_1126_29_7[22:2]) + conv_s2s_21_22(z_out_1013_29_7[22:2]);
  assign AccumDotWidth_acc_2523_nl = nl_AccumDotWidth_acc_2523_nl[21:0];
  assign MultLoop_mux1h_478_nl = MUX1HOT_v_22_8_2(z_out_671_28_7, z_out_664_28_7,
      z_out_397, z_out_426, z_out_401, z_out_383, (AccumDotWidth_acc_2523_nl), (z_out_1110_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_491 = (MultLoop_mux1h_477_nl) + (MultLoop_mux1h_478_nl);
  assign z_out_491 = nl_z_out_491[21:0];
  assign AccumDotWidth_mux1h_1118_nl = MUX1HOT_v_22_4_2(z_out_409, z_out_382, z_out_397,
      z_out_672_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1119_nl = MUX1HOT_v_22_4_2(z_out_408, z_out_381, z_out_400,
      z_out_673_28_7, {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_492 = (AccumDotWidth_mux1h_1118_nl) + (AccumDotWidth_mux1h_1119_nl);
  assign z_out_492 = nl_z_out_492[21:0];
  assign nl_AccumDotWidth_acc_2524_nl = conv_s2s_21_22(z_out_613_29_7[22:2]) + conv_s2s_21_22(z_out_612_29_7[22:2]);
  assign AccumDotWidth_acc_2524_nl = nl_AccumDotWidth_acc_2524_nl[21:0];
  assign nl_AccumDotWidth_acc_2525_nl = conv_s2s_21_22(z_out_620_29_7[22:2]) + conv_s2s_21_22(z_out_974_29_7[22:2]);
  assign AccumDotWidth_acc_2525_nl = nl_AccumDotWidth_acc_2525_nl[21:0];
  assign nl_AccumDotWidth_acc_2526_nl = conv_s2s_21_22(z_out_1035_29_7[22:2]) + conv_s2s_21_22(z_out_1155_29_7[22:2]);
  assign AccumDotWidth_acc_2526_nl = nl_AccumDotWidth_acc_2526_nl[21:0];
  assign AccumDotWidth_mux1h_1120_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2524_nl),
      MultLoop_acc_181_itm, z_out_411, (AccumDotWidth_acc_2525_nl), (AccumDotWidth_acc_2526_nl),
      (z_out_1118_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2527_nl = conv_s2s_21_22(z_out_1015_29_7[22:2]) + conv_s2s_21_22(z_out_1010_29_7[22:2]);
  assign AccumDotWidth_acc_2527_nl = nl_AccumDotWidth_acc_2527_nl[21:0];
  assign nl_AccumDotWidth_acc_2529_nl = (nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2529_nl = nl_AccumDotWidth_acc_2529_nl[9:0];
  assign nl_AccumDotWidth_acc_2528_nl = conv_s2s_21_22({(AccumDotWidth_acc_2529_nl)
      , (nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm[10:0])})
      + conv_s2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm);
  assign AccumDotWidth_acc_2528_nl = nl_AccumDotWidth_acc_2528_nl[21:0];
  assign nl_AccumDotWidth_acc_2530_nl = conv_s2s_21_22(z_out_893_29_7[22:2]) + conv_s2s_21_22(z_out_1183_29_7[22:2]);
  assign AccumDotWidth_acc_2530_nl = nl_AccumDotWidth_acc_2530_nl[21:0];
  assign nl_AccumDotWidth_acc_2531_nl = conv_s2s_21_22(z_out_996_29_7[22:2]) + conv_s2s_21_22(z_out_598_29_7[22:2]);
  assign AccumDotWidth_acc_2531_nl = nl_AccumDotWidth_acc_2531_nl[21:0];
  assign AccumDotWidth_mux1h_1121_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2527_nl),
      (AccumDotWidth_acc_2528_nl), z_out_410, (AccumDotWidth_acc_2530_nl), (AccumDotWidth_acc_2531_nl),
      (z_out_1119_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_493 = (AccumDotWidth_mux1h_1120_nl) + (AccumDotWidth_mux1h_1121_nl);
  assign z_out_493 = nl_z_out_493[21:0];
  assign nl_AccumDotWidth_acc_2532_nl = conv_s2s_21_22(z_out_1008_29_7[22:2]) + conv_s2s_21_22(z_out_878_29_7[22:2]);
  assign AccumDotWidth_acc_2532_nl = nl_AccumDotWidth_acc_2532_nl[21:0];
  assign nl_AccumDotWidth_acc_2533_nl = conv_s2s_21_22(z_out_1153_29_7[22:2]) + conv_s2s_21_22(z_out_943_29_7[22:2]);
  assign AccumDotWidth_acc_2533_nl = nl_AccumDotWidth_acc_2533_nl[21:0];
  assign nl_AccumDotWidth_acc_2534_nl = conv_s2s_21_22(z_out_621_29_7[22:2]) + conv_s2s_21_22(z_out_1121_29_7[22:2]);
  assign AccumDotWidth_acc_2534_nl = nl_AccumDotWidth_acc_2534_nl[21:0];
  assign MultLoop_mux1h_479_nl = MUX1HOT_v_22_6_2(z_out_669_28_7, MultLoop_acc_372_itm,
      (AccumDotWidth_acc_2532_nl), (AccumDotWidth_acc_2533_nl), (AccumDotWidth_acc_2534_nl),
      (z_out_1114_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2536_nl = (nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2536_nl = nl_AccumDotWidth_acc_2536_nl[9:0];
  assign nl_AccumDotWidth_acc_2535_nl = AccumDotWidth_acc_1352_itm + conv_s2s_21_22({(AccumDotWidth_acc_2536_nl)
      , (nnet_relu_layer2_t_layer3_t_relu_config3_for_10_if_exu_pmx_20_0_lpi_1_dfm[10:0])});
  assign AccumDotWidth_acc_2535_nl = nl_AccumDotWidth_acc_2535_nl[21:0];
  assign nl_AccumDotWidth_acc_2537_nl = conv_s2s_21_22(z_out_886_29_7[22:2]) + conv_s2s_21_22(z_out_1031_29_9);
  assign AccumDotWidth_acc_2537_nl = nl_AccumDotWidth_acc_2537_nl[21:0];
  assign nl_AccumDotWidth_acc_2538_nl = conv_s2s_21_22(z_out_1124_29_7[22:2]) + conv_s2s_21_22(z_out_915_29_7[22:2]);
  assign AccumDotWidth_acc_2538_nl = nl_AccumDotWidth_acc_2538_nl[21:0];
  assign nl_AccumDotWidth_acc_2539_nl = conv_s2s_21_22(z_out_1134_29_9) + conv_s2s_21_22(z_out_1016_29_7[22:2]);
  assign AccumDotWidth_acc_2539_nl = nl_AccumDotWidth_acc_2539_nl[21:0];
  assign MultLoop_mux1h_480_nl = MUX1HOT_v_22_6_2(z_out_676_28_7, (AccumDotWidth_acc_2535_nl),
      (AccumDotWidth_acc_2537_nl), (AccumDotWidth_acc_2538_nl), (AccumDotWidth_acc_2539_nl),
      (z_out_1115_29_7[21:0]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_494 = (MultLoop_mux1h_479_nl) + (MultLoop_mux1h_480_nl);
  assign z_out_494 = nl_z_out_494[21:0];
  assign MultLoop_mux1h_481_nl = MUX1HOT_v_22_6_2(z_out_72_28_7, z_out_641_28_7,
      z_out_112_28_7, z_out_129_28_7, z_out_65_28_7, z_out_76_28_7, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_mux1h_482_nl = MUX1HOT_v_22_6_2(z_out_67_28_7, z_out_656_28_7,
      z_out_115_28_7, z_out_130_28_7, z_out_63_28_7, z_out_65_28_7, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_z_out_495 = (MultLoop_mux1h_481_nl) + (MultLoop_mux1h_482_nl);
  assign z_out_495 = nl_z_out_495[21:0];
  assign nl_MultLoop_acc_1522_nl = z_out_762 + MultLoop_acc_1018_itm;
  assign MultLoop_acc_1522_nl = nl_MultLoop_acc_1522_nl[21:0];
  assign MultLoop_mux_95_nl = MUX_v_22_2_2(z_out_84_28_7, (MultLoop_acc_1522_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1523_nl = MultLoop_acc_1007_itm + z_out_537;
  assign MultLoop_acc_1523_nl = nl_MultLoop_acc_1523_nl[21:0];
  assign MultLoop_mux_96_nl = MUX_v_22_2_2(z_out_87_28_7, (MultLoop_acc_1523_nl),
      fsm_output[8]);
  assign nl_z_out_496 = (MultLoop_mux_95_nl) + (MultLoop_mux_96_nl);
  assign z_out_496 = nl_z_out_496[21:0];
  assign MultLoop_mux1h_483_nl = MUX1HOT_v_22_4_2(z_out_137_28_7, z_out_81_28_7,
      z_out_66_28_7, z_out_71_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign MultLoop_mux1h_484_nl = MUX1HOT_v_22_4_2(z_out_68_28_7, z_out_631_28_7,
      z_out_64_28_7, z_out_73_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_497 = (MultLoop_mux1h_483_nl) + (MultLoop_mux1h_484_nl);
  assign z_out_497 = nl_z_out_497[21:0];
  assign MultLoop_mux1h_485_nl = MUX1HOT_v_22_4_2(z_out_672_28_7, z_out_153_28_7,
      MultLoop_acc_128_itm, (z_out_592_29_7[21:0]), {AccumDotWidth_or_152_cse , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[8])});
  assign MultLoop_mux1h_486_nl = MUX1HOT_v_22_4_2(z_out_673_28_7, z_out_148_28_7,
      z_out_425, (z_out_594_29_7[21:0]), {AccumDotWidth_or_152_cse , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_498 = (MultLoop_mux1h_485_nl) + (MultLoop_mux1h_486_nl);
  assign z_out_498 = nl_z_out_498[21:0];
  assign MultLoop_mux1h_487_nl = MUX1HOT_v_22_4_2(z_out_674_28_7, z_out_171_28_7,
      z_out_147_28_7, (z_out_590_29_7[21:0]), {AccumDotWidth_or_152_cse , (fsm_output[7])
      , (fsm_output[2]) , (fsm_output[8])});
  assign MultLoop_mux1h_488_nl = MUX1HOT_v_22_4_2(z_out_675_28_7, z_out_186_28_7,
      z_out_146_28_7, (z_out_591_29_7[21:0]), {AccumDotWidth_or_152_cse , (fsm_output[7])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nl_z_out_499 = (MultLoop_mux1h_487_nl) + (MultLoop_mux1h_488_nl);
  assign z_out_499 = nl_z_out_499[21:0];
  assign AccumDotWidth_mux1h_1122_nl = MUX1HOT_v_22_6_2(z_out_390, MultLoop_acc_243_itm,
      z_out_743, z_out_380, z_out_399, (z_out_611_29_7[21:0]), {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2541_nl = (nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm[20:11])
      + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2541_nl = nl_AccumDotWidth_acc_2541_nl[9:0];
  assign nl_AccumDotWidth_acc_2540_nl = AccumDotWidth_acc_1300_itm + conv_s2s_21_22({(AccumDotWidth_acc_2541_nl)
      , (nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm[10:0])});
  assign AccumDotWidth_acc_2540_nl = nl_AccumDotWidth_acc_2540_nl[21:0];
  assign AccumDotWidth_mux1h_1123_nl = MUX1HOT_v_22_6_2(z_out_391, (AccumDotWidth_acc_2540_nl),
      z_out_742, z_out_377, z_out_398, (z_out_612_29_7[21:0]), {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_500 = (AccumDotWidth_mux1h_1122_nl) + (AccumDotWidth_mux1h_1123_nl);
  assign z_out_500 = nl_z_out_500[21:0];
  assign MultLoop_mux1h_489_nl = MUX1HOT_v_22_4_2(z_out_151_28_7, z_out_667_28_7,
      (z_out_623_29_7[21:0]), (z_out_912_29_7[21:0]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign MultLoop_mux1h_490_nl = MUX1HOT_v_22_4_2(z_out_152_28_7, z_out_668_28_7,
      z_out_160_28_7, (z_out_913_29_7[21:0]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_501 = (MultLoop_mux1h_489_nl) + (MultLoop_mux1h_490_nl);
  assign z_out_501 = nl_z_out_501[21:0];
  assign MultLoop_mux1h_491_nl = MUX1HOT_v_22_4_2((z_out_620_29_7[21:0]), z_out_665_28_7,
      z_out_161_28_7, (z_out_613_29_7[21:0]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign MultLoop_mux1h_492_nl = MUX1HOT_v_22_4_2(z_out_149_28_7, z_out_666_28_7,
      z_out_162_28_7, (z_out_614_29_7[21:0]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_502 = (MultLoop_mux1h_491_nl) + (MultLoop_mux1h_492_nl);
  assign z_out_502 = nl_z_out_502[21:0];
  assign nl_AccumDotWidth_acc_2542_nl = conv_s2s_21_22(z_out_1014_29_7[22:2]) + conv_s2s_21_22(z_out_1017_29_9);
  assign AccumDotWidth_acc_2542_nl = nl_AccumDotWidth_acc_2542_nl[21:0];
  assign nl_AccumDotWidth_acc_2543_nl = conv_s2s_21_22(z_out_586_29_7[22:2]) + conv_s2s_21_22(z_out_1090_29_7[22:2]);
  assign AccumDotWidth_acc_2543_nl = nl_AccumDotWidth_acc_2543_nl[21:0];
  assign nl_AccumDotWidth_acc_2544_nl = conv_s2s_21_22(z_out_608_29_7[22:2]) + conv_s2s_21_22(z_out_615_29_7[22:2]);
  assign AccumDotWidth_acc_2544_nl = nl_AccumDotWidth_acc_2544_nl[21:0];
  assign nl_AccumDotWidth_acc_2545_nl = conv_s2s_21_22(z_out_1071_29_7[22:2]) + conv_s2s_21_22(z_out_1012_29_7[22:2]);
  assign AccumDotWidth_acc_2545_nl = nl_AccumDotWidth_acc_2545_nl[21:0];
  assign AccumDotWidth_mux1h_1124_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2542_nl),
      MultLoop_acc_1007_itm, (AccumDotWidth_acc_2543_nl), (AccumDotWidth_acc_2544_nl),
      (AccumDotWidth_acc_2545_nl), (z_out_619_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2546_nl = conv_s2s_21_22(z_out_1009_29_7[22:2]) + conv_s2s_21_22(z_out_1020_29_9);
  assign AccumDotWidth_acc_2546_nl = nl_AccumDotWidth_acc_2546_nl[21:0];
  assign nl_AccumDotWidth_acc_2547_nl = conv_s2s_21_22(z_out_885_29_7[22:2]) + conv_s2s_21_22(z_out_984_29_7[22:2]);
  assign AccumDotWidth_acc_2547_nl = nl_AccumDotWidth_acc_2547_nl[21:0];
  assign nl_AccumDotWidth_acc_2548_nl = conv_s2s_21_22(z_out_887_29_7[22:2]) + conv_s2s_21_22(z_out_1025_29_7[22:2]);
  assign AccumDotWidth_acc_2548_nl = nl_AccumDotWidth_acc_2548_nl[21:0];
  assign nl_AccumDotWidth_acc_2549_nl = conv_s2s_21_22(z_out_884_29_7[22:2]) + conv_s2s_21_22(z_out_1032_29_9);
  assign AccumDotWidth_acc_2549_nl = nl_AccumDotWidth_acc_2549_nl[21:0];
  assign AccumDotWidth_mux1h_1125_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2546_nl),
      z_out_428, (AccumDotWidth_acc_2547_nl), (AccumDotWidth_acc_2548_nl), (AccumDotWidth_acc_2549_nl),
      (z_out_570_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_503 = (AccumDotWidth_mux1h_1124_nl) + (AccumDotWidth_mux1h_1125_nl);
  assign z_out_503 = nl_z_out_503[21:0];
  assign nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9983:9976]));
  assign MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign MultLoop_mux1h_493_nl = MUX1HOT_v_22_3_2(z_out_159_28_7, z_out_674_28_7,
      (readslicef_29_22_7((MultLoop_1248_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[8])});
  assign nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9991:9984]));
  assign MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign MultLoop_mux1h_494_nl = MUX1HOT_v_22_3_2(z_out_160_28_7, z_out_166_28_7,
      (readslicef_29_22_7((MultLoop_1249_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[6]) , (fsm_output[2]) , (fsm_output[8])});
  assign nl_z_out_504 = (MultLoop_mux1h_493_nl) + (MultLoop_mux1h_494_nl);
  assign z_out_504 = nl_z_out_504[21:0];
  assign MultLoop_mux1h_495_nl = MUX1HOT_v_22_3_2(z_out_65_28_7, z_out_87_28_7, z_out_445,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_496_nl = MUX1HOT_v_22_3_2(z_out_102_28_7, z_out_84_28_7,
      z_out_809, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_505 = (MultLoop_mux1h_495_nl) + (MultLoop_mux1h_496_nl);
  assign z_out_505 = nl_z_out_505[21:0];
  assign MultLoop_mux1h_497_nl = MUX1HOT_v_22_4_2(z_out_66_28_7, z_out_660_28_7,
      z_out_87_28_7, z_out_79_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign MultLoop_mux1h_498_nl = MUX1HOT_v_22_4_2(z_out_633_28_7, z_out_658_28_7,
      z_out_82_28_7, z_out_78_28_7, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_506 = (MultLoop_mux1h_497_nl) + (MultLoop_mux1h_498_nl);
  assign z_out_506 = nl_z_out_506[21:0];
  assign MultLoop_or_107_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[5]);
  assign MultLoop_mux1h_499_nl = MUX1HOT_v_22_3_2(z_out_69_28_7, z_out_35_28_7, z_out_649_28_7,
      {(MultLoop_or_107_nl) , (fsm_output[2]) , (fsm_output[3])});
  assign MultLoop_mux1h_500_nl = MUX1HOT_v_22_5_2(z_out_75_28_7, z_out_34_28_7, z_out_80_28_7,
      z_out_650_28_7, z_out_70_28_7, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_507 = (MultLoop_mux1h_499_nl) + (MultLoop_mux1h_500_nl);
  assign z_out_507 = nl_z_out_507[21:0];
  assign AccumDotWidth_mux1h_1126_nl = MUX1HOT_v_22_6_2(z_out_547, z_out_555, z_out_308,
      z_out_321, z_out_417, z_out_252, {AccumDotWidth_or_149_cse , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1524_nl = (z_out_968_29_7[21:0]) + (z_out_974_29_7[21:0]);
  assign MultLoop_acc_1524_nl = nl_MultLoop_acc_1524_nl[21:0];
  assign AccumDotWidth_mux1h_1127_nl = MUX1HOT_v_22_7_2(z_out_551, z_out_532, z_out_273,
      z_out_264, z_out_414, z_out_549, (MultLoop_acc_1524_nl), {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_508 = (AccumDotWidth_mux1h_1126_nl) + (AccumDotWidth_mux1h_1127_nl);
  assign z_out_508 = nl_z_out_508[21:0];
  assign AccumDotWidth_mux1h_1128_nl = MUX1HOT_v_22_3_2(z_out_532, z_out_413, MultLoop_acc_181_itm,
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1527_nl = (z_out_574_29_7[21:0]) + (z_out_572_29_7[21:0]);
  assign MultLoop_acc_1527_nl = nl_MultLoop_acc_1527_nl[21:0];
  assign nl_MultLoop_acc_1528_nl = (z_out_571_29_7[21:0]) + (z_out_569_29_7[21:0]);
  assign MultLoop_acc_1528_nl = nl_MultLoop_acc_1528_nl[21:0];
  assign nl_MultLoop_acc_1530_nl = (z_out_568_29_7[21:0]) + (z_out_1169_29_7[21:0]);
  assign MultLoop_acc_1530_nl = nl_MultLoop_acc_1530_nl[21:0];
  assign nl_MultLoop_acc_1531_nl = (z_out_1182_29_7[21:0]) + (z_out_1177_29_7[21:0]);
  assign MultLoop_acc_1531_nl = nl_MultLoop_acc_1531_nl[21:0];
  assign nl_MultLoop_acc_1525_nl = (MultLoop_acc_1527_nl) + (MultLoop_acc_1528_nl)
      + (MultLoop_acc_1530_nl) + (MultLoop_acc_1531_nl);
  assign MultLoop_acc_1525_nl = nl_MultLoop_acc_1525_nl[21:0];
  assign AccumDotWidth_mux1h_1129_nl = MUX1HOT_v_22_3_2(z_out_560, z_out_412, (MultLoop_acc_1525_nl),
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_509 = (AccumDotWidth_mux1h_1128_nl) + (AccumDotWidth_mux1h_1129_nl);
  assign z_out_509 = nl_z_out_509[21:0];
  assign AccumDotWidth_mux1h_1130_nl = MUX1HOT_v_22_5_2(z_out_493, z_out_555, z_out_419,
      z_out_532, z_out_249, {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1532_nl = (z_out_1130_29_7[21:0]) + (z_out_1108_29_7[21:0]);
  assign MultLoop_acc_1532_nl = nl_MultLoop_acc_1532_nl[21:0];
  assign AccumDotWidth_mux1h_1131_nl = MUX1HOT_v_22_5_2(MultLoop_acc_105_itm, z_out_500,
      z_out_418, z_out_555, (MultLoop_acc_1532_nl), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_510 = (AccumDotWidth_mux1h_1130_nl) + (AccumDotWidth_mux1h_1131_nl);
  assign z_out_510 = nl_z_out_510[21:0];
  assign nl_MultLoop_acc_1533_nl = (z_out_880_29_7[21:0]) + MultLoop_449_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1533_nl = nl_MultLoop_acc_1533_nl[21:0];
  assign AccumDotWidth_mux1h_1132_nl = MUX1HOT_v_22_4_2(z_out_567, z_out_709, z_out_544,
      (MultLoop_acc_1533_nl), {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1534_nl = (z_out_884_29_7[21:0]) + (z_out_885_29_7[21:0]);
  assign MultLoop_acc_1534_nl = nl_MultLoop_acc_1534_nl[21:0];
  assign AccumDotWidth_mux1h_1133_nl = MUX1HOT_v_22_4_2(z_out_554, z_out_705, z_out_525,
      (MultLoop_acc_1534_nl), {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_511 = (AccumDotWidth_mux1h_1132_nl) + (AccumDotWidth_mux1h_1133_nl);
  assign z_out_511 = nl_z_out_511[21:0];
  assign nl_MultLoop_acc_1535_nl = (z_out_1107_29_7[21:0]) + (z_out_1109_29_7[21:0]);
  assign MultLoop_acc_1535_nl = nl_MultLoop_acc_1535_nl[21:0];
  assign AccumDotWidth_mux1h_1134_nl = MUX1HOT_v_22_3_2(z_out_486, z_out_255, (MultLoop_acc_1535_nl),
      {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1536_nl = (z_out_1091_29_7[21:0]) + (z_out_1078_29_7[21:0]);
  assign MultLoop_acc_1536_nl = nl_MultLoop_acc_1536_nl[21:0];
  assign AccumDotWidth_mux1h_1135_nl = MUX1HOT_v_22_3_2(MultLoop_acc_1121_itm, z_out_269,
      (MultLoop_acc_1536_nl), {(fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_512 = (AccumDotWidth_mux1h_1134_nl) + (AccumDotWidth_mux1h_1135_nl);
  assign z_out_512 = nl_z_out_512[21:0];
  assign AccumDotWidth_mux_139_nl = MUX_v_22_2_2(z_out_250, z_out_264, fsm_output[7]);
  assign AccumDotWidth_mux_140_nl = MUX_v_22_2_2(z_out_267, z_out_275, fsm_output[7]);
  assign nl_z_out_513 = (AccumDotWidth_mux_139_nl) + (AccumDotWidth_mux_140_nl);
  assign z_out_513 = nl_z_out_513[21:0];
  assign AccumDotWidth_mux1h_1136_nl = MUX1HOT_v_22_3_2(z_out_500, z_out_703, z_out_502,
      {(fsm_output[3]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1137_nl = MUX1HOT_v_22_3_2(MultLoop_acc_113_itm, z_out_701,
      z_out_501, {(fsm_output[3]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_514 = (AccumDotWidth_mux1h_1136_nl) + (AccumDotWidth_mux1h_1137_nl);
  assign z_out_514 = nl_z_out_514[21:0];
  assign nl_MultLoop_acc_1537_nl = (z_out_1168_29_7[21:0]) + (z_out_1155_29_7[21:0]);
  assign MultLoop_acc_1537_nl = nl_MultLoop_acc_1537_nl[21:0];
  assign AccumDotWidth_mux_141_nl = MUX_v_22_2_2(z_out_251, (MultLoop_acc_1537_nl),
      fsm_output[8]);
  assign nl_MultLoop_acc_1538_nl = (z_out_618_29_7[21:0]) + (z_out_617_29_7[21:0]);
  assign MultLoop_acc_1538_nl = nl_MultLoop_acc_1538_nl[21:0];
  assign AccumDotWidth_mux_142_nl = MUX_v_22_2_2(z_out_270, (MultLoop_acc_1538_nl),
      fsm_output[8]);
  assign nl_z_out_515 = (AccumDotWidth_mux_141_nl) + (AccumDotWidth_mux_142_nl);
  assign z_out_515 = nl_z_out_515[21:0];
  assign nl_MultLoop_acc_1539_nl = (z_out_1165_29_7[21:0]) + (z_out_1163_29_7[21:0]);
  assign MultLoop_acc_1539_nl = nl_MultLoop_acc_1539_nl[21:0];
  assign AccumDotWidth_mux1h_1138_nl = MUX1HOT_v_22_8_2(z_out_736, z_out_688, z_out_421,
      z_out_687, z_out_801, z_out_727, z_out_680, (MultLoop_acc_1539_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1540_nl = (z_out_1167_29_7[21:0]) + (z_out_1159_29_7[21:0]);
  assign MultLoop_acc_1540_nl = nl_MultLoop_acc_1540_nl[21:0];
  assign AccumDotWidth_mux1h_1139_nl = MUX1HOT_v_22_8_2(z_out_738, z_out_730, z_out_416,
      z_out_372, z_out_797, z_out_729, z_out_682, (MultLoop_acc_1540_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_516 = (AccumDotWidth_mux1h_1138_nl) + (AccumDotWidth_mux1h_1139_nl);
  assign z_out_516 = nl_z_out_516[21:0];
  assign nl_MultLoop_acc_1541_nl = (z_out_914_29_7[21:0]) + (z_out_915_29_7[21:0]);
  assign MultLoop_acc_1541_nl = nl_MultLoop_acc_1541_nl[21:0];
  assign AccumDotWidth_mux1h_1140_nl = MUX1HOT_v_22_6_2(z_out_725, z_out_683, z_out_412,
      z_out_308, z_out_730, (MultLoop_acc_1541_nl), {(fsm_output[2]) , AccumDotWidth_or_150_cse
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1542_nl = (z_out_1166_29_7[21:0]) + (z_out_1164_29_7[21:0]);
  assign MultLoop_acc_1542_nl = nl_MultLoop_acc_1542_nl[21:0];
  assign AccumDotWidth_mux1h_1141_nl = MUX1HOT_v_22_8_2(z_out_730, z_out_723, z_out_420,
      z_out_375, z_out_337, z_out_728, z_out_388, (MultLoop_acc_1542_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_517 = (AccumDotWidth_mux1h_1140_nl) + (AccumDotWidth_mux1h_1141_nl);
  assign z_out_517 = nl_z_out_517[21:0];
  assign nl_AccumDotWidth_acc_2550_nl = z_out_234 + z_out_235;
  assign AccumDotWidth_acc_2550_nl = nl_AccumDotWidth_acc_2550_nl[21:0];
  assign AccumDotWidth_mux1h_1142_nl = MUX1HOT_v_22_6_2(z_out_715, z_out_349, z_out_241,
      (AccumDotWidth_acc_2550_nl), z_out_516, z_out_250, {(fsm_output[2]) , (fsm_output[3])
      , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1543_nl = (z_out_1049_29_7[21:0]) + (z_out_1034_29_7[21:0]);
  assign MultLoop_acc_1543_nl = nl_MultLoop_acc_1543_nl[21:0];
  assign AccumDotWidth_mux1h_1143_nl = MUX1HOT_v_22_7_2(z_out_718, z_out_374, z_out_526,
      z_out_241, z_out_242, z_out_321, (MultLoop_acc_1543_nl), {(fsm_output[2]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_518 = (AccumDotWidth_mux1h_1142_nl) + (AccumDotWidth_mux1h_1143_nl);
  assign z_out_518 = nl_z_out_518[21:0];
  assign AccumDotWidth_mux1h_1144_nl = MUX1HOT_v_22_7_2(z_out_261, z_out_252, z_out_255,
      z_out_320, z_out_245, z_out_250, z_out_251, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1544_nl = (z_out_969_29_7[21:0]) + (z_out_970_29_7[21:0]);
  assign MultLoop_acc_1544_nl = nl_MultLoop_acc_1544_nl[21:0];
  assign AccumDotWidth_mux1h_1145_nl = MUX1HOT_v_22_7_2(z_out_794, z_out_254, z_out_558,
      z_out_323, z_out_521, z_out_263, (MultLoop_acc_1544_nl), {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_519 = (AccumDotWidth_mux1h_1144_nl) + (AccumDotWidth_mux1h_1145_nl);
  assign z_out_519 = nl_z_out_519[21:0];
  assign nl_AccumDotWidth_acc_2551_nl = conv_s2s_21_22(z_out_1141_29_9) + conv_s2s_21_22(z_out_1037_29_7[22:2]);
  assign AccumDotWidth_acc_2551_nl = nl_AccumDotWidth_acc_2551_nl[21:0];
  assign nl_MultLoop_acc_1545_nl = (z_out_887_29_7[21:0]) + (z_out_876_29_7[21:0]);
  assign MultLoop_acc_1545_nl = nl_MultLoop_acc_1545_nl[21:0];
  assign AccumDotWidth_mux1h_1146_nl = MUX1HOT_v_22_6_2(z_out_780, z_out_498, z_out_733,
      AccumDotWidth_acc_1181_itm, (AccumDotWidth_acc_2551_nl), (MultLoop_acc_1545_nl),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2552_nl = conv_s2s_21_22(z_out_1138_29_9) + conv_s2s_21_22(z_out_1008_29_7[22:2]);
  assign AccumDotWidth_acc_2552_nl = nl_AccumDotWidth_acc_2552_nl[21:0];
  assign nl_MultLoop_acc_1546_nl = (z_out_865_29_7[21:0]) + (z_out_1146_29_7[21:0]);
  assign MultLoop_acc_1546_nl = nl_MultLoop_acc_1546_nl[21:0];
  assign AccumDotWidth_mux1h_1147_nl = MUX1HOT_v_22_6_2(AccumDotWidth_acc_1167_itm,
      MultLoop_acc_1010_itm, z_out_741, z_out_352, (AccumDotWidth_acc_2552_nl), (MultLoop_acc_1546_nl),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_520 = (AccumDotWidth_mux1h_1146_nl) + (AccumDotWidth_mux1h_1147_nl);
  assign z_out_520 = nl_z_out_520[21:0];
  assign AccumDotWidth_mux1h_1148_nl = MUX1HOT_v_22_6_2(z_out_848, z_out_375, z_out_554,
      z_out_740, z_out_704, z_out_552, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1149_nl = MUX1HOT_v_22_6_2(z_out_849, z_out_376, z_out_553,
      z_out_738, z_out_706, z_out_551, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_521 = (AccumDotWidth_mux1h_1148_nl) + (AccumDotWidth_mux1h_1149_nl);
  assign z_out_521 = nl_z_out_521[21:0];
  assign AccumDotWidth_mux1h_1150_nl = MUX1HOT_v_22_5_2(z_out_806, z_out_314, z_out_551,
      z_out_322, z_out_805, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1151_nl = MUX1HOT_v_22_5_2(z_out_795, z_out_567, z_out_547,
      z_out_271, z_out_804, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7])});
  assign nl_z_out_522 = (AccumDotWidth_mux1h_1150_nl) + (AccumDotWidth_mux1h_1151_nl);
  assign z_out_522 = nl_z_out_522[21:0];
  assign AccumDotWidth_mux1h_1152_nl = MUX1HOT_v_22_6_2(z_out_549, z_out_408, z_out_311,
      z_out_545, z_out_416, z_out_557, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1153_nl = MUX1HOT_v_22_6_2(z_out_545, z_out_378, z_out_308,
      z_out_549, z_out_415, z_out_559, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_523 = (AccumDotWidth_mux1h_1152_nl) + (AccumDotWidth_mux1h_1153_nl);
  assign z_out_523 = nl_z_out_523[21:0];
  assign AccumDotWidth_mux1h_1154_nl = MUX1HOT_v_22_7_2(z_out_366, z_out_716, z_out_415,
      z_out_684, z_out_795, z_out_724, z_out_735, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1155_nl = MUX1HOT_v_22_7_2(z_out_367, z_out_720, z_out_418,
      z_out_368, z_out_851, z_out_722, z_out_732, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_524 = (AccumDotWidth_mux1h_1154_nl) + (AccumDotWidth_mux1h_1155_nl);
  assign z_out_524 = nl_z_out_524[21:0];
  assign nl_AccumDotWidth_acc_2553_nl = conv_s2s_21_22(z_out_962_29_9) + conv_s2s_21_22(z_out_1105_29_7[22:2]);
  assign AccumDotWidth_acc_2553_nl = nl_AccumDotWidth_acc_2553_nl[21:0];
  assign nl_AccumDotWidth_acc_2554_nl = conv_s2s_21_22(z_out_1096_29_7[22:2]) + conv_s2s_21_22(z_out_1097_29_7[22:2]);
  assign AccumDotWidth_acc_2554_nl = nl_AccumDotWidth_acc_2554_nl[21:0];
  assign nl_AccumDotWidth_acc_2555_nl = conv_s2s_21_22(z_out_1171_29_7[22:2]) + conv_s2s_21_22(z_out_1042_29_7[22:2]);
  assign AccumDotWidth_acc_2555_nl = nl_AccumDotWidth_acc_2555_nl[21:0];
  assign nl_AccumDotWidth_acc_2556_nl = conv_s2s_21_22(z_out_585_29_7[22:2]) + conv_s2s_21_22(z_out_1083_29_7[22:2]);
  assign AccumDotWidth_acc_2556_nl = nl_AccumDotWidth_acc_2556_nl[21:0];
  assign nl_AccumDotWidth_acc_2557_nl = conv_s2s_21_22(z_out_906_29_7[22:2]) + conv_s2s_21_22(z_out_1093_29_7[22:2]);
  assign AccumDotWidth_acc_2557_nl = nl_AccumDotWidth_acc_2557_nl[21:0];
  assign nl_AccumDotWidth_acc_2558_nl = conv_s2s_21_22(z_out_911_29_7[22:2]) + conv_s2s_21_22(z_out_1080_29_7[22:2]);
  assign AccumDotWidth_acc_2558_nl = nl_AccumDotWidth_acc_2558_nl[21:0];
  assign nl_AccumDotWidth_acc_2559_nl = conv_s2s_21_22(z_out_1068_29_7[22:2]) + conv_s2s_21_22(z_out_1114_29_7[22:2]);
  assign AccumDotWidth_acc_2559_nl = nl_AccumDotWidth_acc_2559_nl[21:0];
  assign AccumDotWidth_mux1h_1156_nl = MUX1HOT_v_22_8_2((AccumDotWidth_acc_2553_nl),
      (AccumDotWidth_acc_2554_nl), (AccumDotWidth_acc_2555_nl), (AccumDotWidth_acc_2556_nl),
      (AccumDotWidth_acc_2557_nl), (AccumDotWidth_acc_2558_nl), (AccumDotWidth_acc_2559_nl),
      z_out_180_28_7, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2560_nl = conv_s2s_21_22(z_out_1027_29_7[22:2]) + conv_s2s_21_22(z_out_1186_29_7[22:2]);
  assign AccumDotWidth_acc_2560_nl = nl_AccumDotWidth_acc_2560_nl[21:0];
  assign nl_AccumDotWidth_acc_2561_nl = conv_s2s_21_22(z_out_1023_29_7[22:2]) + conv_s2s_21_22(z_out_1029_29_7[22:2]);
  assign AccumDotWidth_acc_2561_nl = nl_AccumDotWidth_acc_2561_nl[21:0];
  assign nl_AccumDotWidth_acc_2562_nl = conv_s2s_21_22(z_out_939_29_7[22:2]) + conv_s2s_21_22(z_out_1070_29_7[22:2]);
  assign AccumDotWidth_acc_2562_nl = nl_AccumDotWidth_acc_2562_nl[21:0];
  assign nl_AccumDotWidth_acc_2563_nl = conv_s2s_21_22(z_out_887_29_7[22:2]) + conv_s2s_21_22(z_out_985_29_7[22:2]);
  assign AccumDotWidth_acc_2563_nl = nl_AccumDotWidth_acc_2563_nl[21:0];
  assign nl_AccumDotWidth_acc_2564_nl = conv_s2s_21_22(z_out_918_29_7[22:2]) + conv_s2s_21_22(z_out_1184_29_7[22:2]);
  assign AccumDotWidth_acc_2564_nl = nl_AccumDotWidth_acc_2564_nl[21:0];
  assign nl_AccumDotWidth_acc_2565_nl = conv_s2s_21_22(z_out_854_29_7[22:2]) + conv_s2s_21_22(z_out_963_29_9);
  assign AccumDotWidth_acc_2565_nl = nl_AccumDotWidth_acc_2565_nl[21:0];
  assign nl_AccumDotWidth_acc_2566_nl = conv_s2s_21_22(z_out_886_29_7[22:2]) + conv_s2s_21_22(z_out_1031_29_9);
  assign AccumDotWidth_acc_2566_nl = nl_AccumDotWidth_acc_2566_nl[21:0];
  assign AccumDotWidth_mux1h_1157_nl = MUX1HOT_v_22_8_2((AccumDotWidth_acc_2560_nl),
      (AccumDotWidth_acc_2561_nl), (AccumDotWidth_acc_2562_nl), (AccumDotWidth_acc_2563_nl),
      (AccumDotWidth_acc_2564_nl), (AccumDotWidth_acc_2565_nl), (AccumDotWidth_acc_2566_nl),
      z_out_178_28_7, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_525 = (AccumDotWidth_mux1h_1156_nl) + (AccumDotWidth_mux1h_1157_nl);
  assign z_out_525 = nl_z_out_525[21:0];
  assign AccumDotWidth_mux1h_1158_nl = MUX1HOT_v_22_6_2(z_out_713, z_out_560, z_out_413,
      z_out_688, z_out_799, z_out_361, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1159_nl = MUX1HOT_v_22_7_2(z_out_727, z_out_799, z_out_419,
      z_out_369, z_out_334, z_out_355, z_out_381, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_526 = (AccumDotWidth_mux1h_1158_nl) + (AccumDotWidth_mux1h_1159_nl);
  assign z_out_526 = nl_z_out_526[21:0];
  assign nl_AccumDotWidth_acc_2567_nl = conv_s2s_21_22(z_out_969_29_7[22:2]) + conv_s2s_21_22(z_out_939_29_7[22:2])
      + conv_s2s_21_22(z_out_1107_29_7[22:2]) + conv_s2s_21_22(z_out_1034_29_7[22:2]);
  assign AccumDotWidth_acc_2567_nl = nl_AccumDotWidth_acc_2567_nl[21:0];
  assign AccumDotWidth_mux1h_1160_nl = MUX1HOT_v_22_7_2(z_out_737, z_out_368, z_out_730,
      z_out_354, (AccumDotWidth_acc_2567_nl), z_out_711, z_out_552, {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2570_nl = conv_s2s_21_22(z_out_1071_29_7[22:2]) + conv_s2s_21_22(z_out_873_29_7[22:2])
      + conv_s2s_21_22(z_out_1126_29_7[22:2]) + conv_s2s_21_22(z_out_1017_29_9);
  assign AccumDotWidth_acc_2570_nl = nl_AccumDotWidth_acc_2570_nl[21:0];
  assign AccumDotWidth_mux1h_1161_nl = MUX1HOT_v_22_6_2(z_out_733, z_out_370, z_out_725,
      (AccumDotWidth_acc_2570_nl), z_out_702, z_out_553, {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , AccumDotWidth_or_132_cse_1 , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_527 = (AccumDotWidth_mux1h_1160_nl) + (AccumDotWidth_mux1h_1161_nl);
  assign z_out_527 = nl_z_out_527[21:0];
  assign AccumDotWidth_mux1h_1162_nl = MUX1HOT_v_22_5_2(z_out_729, z_out_685, z_out_417,
      z_out_793, z_out_708, {(fsm_output[2]) , AccumDotWidth_or_150_cse , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1163_nl = MUX1HOT_v_22_7_2(z_out_728, z_out_713, z_out_414,
      z_out_374, z_out_348, z_out_710, z_out_393, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_528 = (AccumDotWidth_mux1h_1162_nl) + (AccumDotWidth_mux1h_1163_nl);
  assign z_out_528 = nl_z_out_528[21:0];
  assign AccumDotWidth_mux1h_1164_nl = MUX1HOT_v_22_8_2(z_out_362, z_out_567, z_out_708,
      z_out_681, z_out_852, z_out_357, z_out_734, AccumDotWidth_acc_1392_itm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1547_nl = z_out_499 + z_out_498;
  assign MultLoop_acc_1547_nl = nl_MultLoop_acc_1547_nl[21:0];
  assign AccumDotWidth_mux1h_1165_nl = MUX1HOT_v_22_8_2(z_out_374, z_out_532, z_out_701,
      z_out_373, z_out_402, z_out_364, z_out_738, (MultLoop_acc_1547_nl), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_529 = (AccumDotWidth_mux1h_1164_nl) + (AccumDotWidth_mux1h_1165_nl);
  assign z_out_529 = nl_z_out_529[21:0];
  assign nl_AccumDotWidth_acc_2573_nl = z_out_536 + z_out_516;
  assign AccumDotWidth_acc_2573_nl = nl_AccumDotWidth_acc_2573_nl[21:0];
  assign AccumDotWidth_mux1h_1166_nl = MUX1HOT_v_22_8_2(z_out_705, z_out_684, z_out_737,
      z_out_511, (AccumDotWidth_acc_2573_nl), z_out_323, z_out_543, z_out_271, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1167_nl = MUX1HOT_v_22_7_2(z_out_708, z_out_354, z_out_736,
      z_out_321, z_out_240, z_out_234, AccumDotWidth_acc_1397_itm, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_152_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_530 = (AccumDotWidth_mux1h_1166_nl) + (AccumDotWidth_mux1h_1167_nl);
  assign z_out_530 = nl_z_out_530[21:0];
  assign nl_AccumDotWidth_acc_2574_nl = z_out_701 + z_out_706;
  assign AccumDotWidth_acc_2574_nl = nl_AccumDotWidth_acc_2574_nl[21:0];
  assign AccumDotWidth_mux1h_1168_nl = MUX1HOT_v_22_7_2(z_out_371, z_out_556, z_out_546,
      (AccumDotWidth_acc_2574_nl), z_out_726, z_out_687, AccumDotWidth_acc_1352_itm,
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2576_nl = (z_out_905_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2576_nl = nl_AccumDotWidth_acc_2576_nl[9:0];
  assign nl_AccumDotWidth_acc_2575_nl = z_out_704 + conv_s2s_21_22({(AccumDotWidth_acc_2576_nl)
      , (z_out_905_29_7[12:2])});
  assign AccumDotWidth_acc_2575_nl = nl_AccumDotWidth_acc_2575_nl[21:0];
  assign AccumDotWidth_mux1h_1169_nl = MUX1HOT_v_22_7_2(z_out_373, z_out_557, AccumDotWidth_acc_1201_itm,
      (AccumDotWidth_acc_2575_nl), z_out_723, z_out_383, z_out_520, {(fsm_output[2])
      , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_531 = (AccumDotWidth_mux1h_1168_nl) + (AccumDotWidth_mux1h_1169_nl);
  assign z_out_531 = nl_z_out_531[21:0];
  assign AccumDotWidth_mux1h_1170_nl = MUX1HOT_v_22_6_2(z_out_748, z_out_744, z_out_700,
      z_out_391, z_out_369, z_out_365, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1171_nl = MUX1HOT_v_22_5_2(z_out_744, z_out_745, z_out_693,
      z_out_390, z_out_368, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , AccumDotWidth_or_140_cse});
  assign nl_z_out_532 = (AccumDotWidth_mux1h_1170_nl) + (AccumDotWidth_mux1h_1171_nl);
  assign z_out_532 = nl_z_out_532[21:0];
  assign AccumDotWidth_mux1h_1172_nl = MUX1HOT_v_22_8_2(z_out_709, z_out_687, z_out_734,
      z_out_320, z_out_543, z_out_321, z_out_540, AccumDotWidth_acc_1164_itm, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1173_nl = MUX1HOT_v_22_8_2(z_out_722, z_out_688, z_out_738,
      z_out_527, z_out_236, z_out_337, z_out_242, z_out_835, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_533 = (AccumDotWidth_mux1h_1172_nl) + (AccumDotWidth_mux1h_1173_nl);
  assign z_out_533 = nl_z_out_533[21:0];
  assign AccumDotWidth_mux1h_1174_nl = MUX1HOT_v_22_8_2(z_out_423, z_out_700, z_out_330,
      z_out_234, z_out_318, z_out_557, z_out_564, z_out_269, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1175_nl = MUX1HOT_v_22_8_2(z_out_433, z_out_703, z_out_234,
      z_out_528, z_out_246, z_out_559, z_out_241, AccumDotWidth_acc_1235_itm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_534 = (AccumDotWidth_mux1h_1174_nl) + (AccumDotWidth_mux1h_1175_nl);
  assign z_out_534 = nl_z_out_534[21:0];
  assign nl_AccumDotWidth_acc_2577_nl = z_out_283 + z_out_842;
  assign AccumDotWidth_acc_2577_nl = nl_AccumDotWidth_acc_2577_nl[21:0];
  assign AccumDotWidth_mux1h_1176_nl = MUX1HOT_v_22_8_2(z_out_382, z_out_363, (AccumDotWidth_acc_2577_nl),
      z_out_229, z_out_317, z_out_318, z_out_539, z_out_831, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1177_nl = MUX1HOT_v_22_8_2(z_out_392, z_out_359, z_out_229,
      z_out_517, z_out_522, z_out_237, z_out_238, AccumDotWidth_acc_1167_itm, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_535 = (AccumDotWidth_mux1h_1176_nl) + (AccumDotWidth_mux1h_1177_nl);
  assign z_out_535 = nl_z_out_535[21:0];
  assign AccumDotWidth_mux1h_1178_nl = MUX1HOT_v_22_6_2(z_out_352, z_out_702, z_out_341,
      z_out_253, z_out_806, z_out_514, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1179_nl = MUX1HOT_v_22_6_2(z_out_365, z_out_714, z_out_400,
      AccumDotWidth_acc_1167_itm, z_out_794, z_out_520, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign nl_z_out_536 = (AccumDotWidth_mux1h_1178_nl) + (AccumDotWidth_mux1h_1179_nl);
  assign z_out_536 = nl_z_out_536[21:0];
  assign AccumDotWidth_mux1h_1180_nl = MUX1HOT_v_22_3_2(z_out_235, z_out_526, z_out_286,
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1550_nl = (z_out_855_29_7[21:0]) + (z_out_858_29_7[21:0]);
  assign MultLoop_acc_1550_nl = nl_MultLoop_acc_1550_nl[21:0];
  assign nl_MultLoop_acc_1551_nl = (z_out_859_29_7[21:0]) + (z_out_1073_29_7[21:0]);
  assign MultLoop_acc_1551_nl = nl_MultLoop_acc_1551_nl[21:0];
  assign nl_MultLoop_acc_1553_nl = (z_out_1074_29_7[21:0]) + (z_out_1075_29_7[21:0]);
  assign MultLoop_acc_1553_nl = nl_MultLoop_acc_1553_nl[21:0];
  assign nl_MultLoop_acc_1554_nl = (z_out_1081_29_7[21:0]) + (z_out_1077_29_7[21:0]);
  assign MultLoop_acc_1554_nl = nl_MultLoop_acc_1554_nl[21:0];
  assign nl_MultLoop_acc_1548_nl = (MultLoop_acc_1550_nl) + (MultLoop_acc_1551_nl)
      + (MultLoop_acc_1553_nl) + (MultLoop_acc_1554_nl);
  assign MultLoop_acc_1548_nl = nl_MultLoop_acc_1548_nl[21:0];
  assign AccumDotWidth_mux1h_1181_nl = MUX1HOT_v_22_3_2(z_out_516, z_out_331, (MultLoop_acc_1548_nl),
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_537 = (AccumDotWidth_mux1h_1180_nl) + (AccumDotWidth_mux1h_1181_nl);
  assign z_out_537 = nl_z_out_537[21:0];
  assign AccumDotWidth_mux1h_1182_nl = MUX1HOT_v_22_5_2(z_out_353, z_out_326, z_out_319,
      z_out_523, z_out_463, {(fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1183_nl = MUX1HOT_v_22_6_2(z_out_351, z_out_241, z_out_524,
      z_out_239, z_out_509, z_out_458, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_538 = (AccumDotWidth_mux1h_1182_nl) + (AccumDotWidth_mux1h_1183_nl);
  assign z_out_538 = nl_z_out_538[21:0];
  assign nl_MultLoop_acc_1557_nl = (z_out_1069_29_7[21:0]) + (z_out_1068_29_7[21:0]);
  assign MultLoop_acc_1557_nl = nl_MultLoop_acc_1557_nl[21:0];
  assign nl_MultLoop_acc_1558_nl = (z_out_1054_29_7[21:0]) + (z_out_1058_29_7[21:0]);
  assign MultLoop_acc_1558_nl = nl_MultLoop_acc_1558_nl[21:0];
  assign nl_MultLoop_acc_1556_nl = (MultLoop_acc_1557_nl) + (MultLoop_acc_1558_nl);
  assign MultLoop_acc_1556_nl = nl_MultLoop_acc_1556_nl[21:0];
  assign nl_MultLoop_acc_1555_nl = z_out_547 + (MultLoop_acc_1556_nl);
  assign MultLoop_acc_1555_nl = nl_MultLoop_acc_1555_nl[21:0];
  assign AccumDotWidth_mux1h_1184_nl = MUX1HOT_v_22_4_2(z_out_262, z_out_261, z_out_251,
      (MultLoop_acc_1555_nl), {AccumDotWidth_or_132_cse_1 , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1561_nl = (z_out_1055_29_7[21:0]) + (z_out_1052_29_7[21:0]);
  assign MultLoop_acc_1561_nl = nl_MultLoop_acc_1561_nl[21:0];
  assign nl_MultLoop_acc_1562_nl = (z_out_1050_29_7[21:0]) + (z_out_1057_29_7[21:0]);
  assign MultLoop_acc_1562_nl = nl_MultLoop_acc_1562_nl[21:0];
  assign nl_MultLoop_acc_1564_nl = (z_out_1051_29_7[21:0]) + (z_out_936_29_7[21:0]);
  assign MultLoop_acc_1564_nl = nl_MultLoop_acc_1564_nl[21:0];
  assign nl_MultLoop_acc_1565_nl = (z_out_937_29_7[21:0]) + (z_out_1053_29_7[21:0]);
  assign MultLoop_acc_1565_nl = nl_MultLoop_acc_1565_nl[21:0];
  assign nl_MultLoop_acc_1559_nl = (MultLoop_acc_1561_nl) + (MultLoop_acc_1562_nl)
      + (MultLoop_acc_1564_nl) + (MultLoop_acc_1565_nl);
  assign MultLoop_acc_1559_nl = nl_MultLoop_acc_1559_nl[21:0];
  assign AccumDotWidth_mux1h_1185_nl = MUX1HOT_v_22_5_2(z_out_565, z_out_797, z_out_262,
      z_out_842, (MultLoop_acc_1559_nl), {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_539 = (AccumDotWidth_mux1h_1184_nl) + (AccumDotWidth_mux1h_1185_nl);
  assign z_out_539 = nl_z_out_539[21:0];
  assign AccumDotWidth_mux1h_1186_nl = MUX1HOT_v_22_5_2(z_out_717, z_out_245, z_out_251,
      z_out_260, z_out_841, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1187_nl = MUX1HOT_v_22_5_2(z_out_719, z_out_244, z_out_328,
      z_out_315, AccumDotWidth_acc_1218_itm, {(fsm_output[2]) , (fsm_output[3]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_540 = (AccumDotWidth_mux1h_1186_nl) + (AccumDotWidth_mux1h_1187_nl);
  assign z_out_540 = nl_z_out_540[21:0];
  assign nl_MultLoop_acc_1568_nl = (z_out_627_29_7[21:0]) + (z_out_626_29_7[21:0]);
  assign MultLoop_acc_1568_nl = nl_MultLoop_acc_1568_nl[21:0];
  assign nl_MultLoop_acc_1569_nl = (z_out_625_29_7[21:0]) + (z_out_624_29_7[21:0]);
  assign MultLoop_acc_1569_nl = nl_MultLoop_acc_1569_nl[21:0];
  assign nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9759:9752]));
  assign MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9767:9760]));
  assign MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1571_nl = (readslicef_29_22_7((MultLoop_1220_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1221_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1571_nl = nl_MultLoop_acc_1571_nl[21:0];
  assign nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9775:9768]));
  assign MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9783:9776]));
  assign MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1572_nl = (readslicef_29_22_7((MultLoop_1222_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1223_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1572_nl = nl_MultLoop_acc_1572_nl[21:0];
  assign nl_MultLoop_acc_1566_nl = (MultLoop_acc_1568_nl) + (MultLoop_acc_1569_nl)
      + (MultLoop_acc_1571_nl) + (MultLoop_acc_1572_nl);
  assign MultLoop_acc_1566_nl = nl_MultLoop_acc_1566_nl[21:0];
  assign AccumDotWidth_mux1h_1188_nl = MUX1HOT_v_22_5_2(z_out_255, z_out_345, z_out_256,
      z_out_254, (MultLoop_acc_1566_nl), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse , (fsm_output[8])});
  assign nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9791:9784]));
  assign MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9799:9792]));
  assign MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1575_nl = (readslicef_29_22_7((MultLoop_1224_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1225_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1575_nl = nl_MultLoop_acc_1575_nl[21:0];
  assign nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9807:9800]));
  assign MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1576_nl = (readslicef_29_22_7((MultLoop_1226_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + z_out_193_28_7;
  assign MultLoop_acc_1576_nl = nl_MultLoop_acc_1576_nl[21:0];
  assign nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9831:9824]));
  assign MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1578_nl = (z_out_622_29_7[21:0]) + (readslicef_29_22_7((MultLoop_1229_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1578_nl = nl_MultLoop_acc_1578_nl[21:0];
  assign nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9839:9832]));
  assign MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9847:9840]));
  assign MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1579_nl = (readslicef_29_22_7((MultLoop_1230_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1231_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1579_nl = nl_MultLoop_acc_1579_nl[21:0];
  assign nl_MultLoop_acc_1573_nl = (MultLoop_acc_1575_nl) + (MultLoop_acc_1576_nl)
      + (MultLoop_acc_1578_nl) + (MultLoop_acc_1579_nl);
  assign MultLoop_acc_1573_nl = nl_MultLoop_acc_1573_nl[21:0];
  assign AccumDotWidth_mux1h_1189_nl = MUX1HOT_v_22_6_2(z_out_778, z_out_373, z_out_848,
      z_out_313, z_out_261, (MultLoop_acc_1573_nl), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_541 = (AccumDotWidth_mux1h_1188_nl) + (AccumDotWidth_mux1h_1189_nl);
  assign z_out_541 = nl_z_out_541[21:0];
  assign nl_AccumDotWidth_acc_2578_nl = z_out_850 + z_out_835 + z_out_778 + z_out_844;
  assign AccumDotWidth_acc_2578_nl = nl_AccumDotWidth_acc_2578_nl[21:0];
  assign AccumDotWidth_mux1h_1190_nl = MUX1HOT_v_22_5_2(z_out_355, z_out_342, z_out_242,
      (AccumDotWidth_acc_2578_nl), z_out_453, {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1191_nl = MUX1HOT_v_22_5_2(z_out_361, z_out_397, z_out_529,
      z_out_237, z_out_459, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_542 = (AccumDotWidth_mux1h_1190_nl) + (AccumDotWidth_mux1h_1191_nl);
  assign z_out_542 = nl_z_out_542[21:0];
  assign nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_48_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9599:9592]));
  assign MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_49_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9607:9600]));
  assign MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1582_nl = (readslicef_29_22_7((MultLoop_1200_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1201_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1582_nl = nl_MultLoop_acc_1582_nl[21:0];
  assign nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_50_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9615:9608]));
  assign MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_51_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9623:9616]));
  assign MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1583_nl = (readslicef_29_22_7((MultLoop_1202_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1203_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1583_nl = nl_MultLoop_acc_1583_nl[21:0];
  assign nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9631:9624]));
  assign MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9639:9632]));
  assign MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1585_nl = (readslicef_29_22_7((MultLoop_1204_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1205_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1585_nl = nl_MultLoop_acc_1585_nl[21:0];
  assign nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9647:9640]));
  assign MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9655:9648]));
  assign MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1586_nl = (readslicef_29_22_7((MultLoop_1206_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1207_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1586_nl = nl_MultLoop_acc_1586_nl[21:0];
  assign nl_MultLoop_acc_1580_nl = (MultLoop_acc_1582_nl) + (MultLoop_acc_1583_nl)
      + (MultLoop_acc_1585_nl) + (MultLoop_acc_1586_nl);
  assign MultLoop_acc_1580_nl = nl_MultLoop_acc_1580_nl[21:0];
  assign AccumDotWidth_mux1h_1192_nl = MUX1HOT_v_22_6_2(z_out_251, z_out_351, z_out_261,
      z_out_324, z_out_257, (MultLoop_acc_1580_nl), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9663:9656]));
  assign MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9671:9664]));
  assign MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1589_nl = (readslicef_29_22_7((MultLoop_1208_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1209_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1589_nl = nl_MultLoop_acc_1589_nl[21:0];
  assign nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9679:9672]));
  assign MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9687:9680]));
  assign MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1590_nl = (readslicef_29_22_7((MultLoop_1210_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1211_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1590_nl = nl_MultLoop_acc_1590_nl[21:0];
  assign nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9695:9688]));
  assign MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9703:9696]));
  assign MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1592_nl = (readslicef_29_22_7((MultLoop_1212_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_1213_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1592_nl = nl_MultLoop_acc_1592_nl[21:0];
  assign nl_MultLoop_acc_1593_nl = (z_out_629_29_7[21:0]) + (z_out_628_29_7[21:0]);
  assign MultLoop_acc_1593_nl = nl_MultLoop_acc_1593_nl[21:0];
  assign nl_MultLoop_acc_1587_nl = (MultLoop_acc_1589_nl) + (MultLoop_acc_1590_nl)
      + (MultLoop_acc_1592_nl) + (MultLoop_acc_1593_nl);
  assign MultLoop_acc_1587_nl = nl_MultLoop_acc_1587_nl[21:0];
  assign AccumDotWidth_mux1h_1193_nl = MUX1HOT_v_22_6_2(z_out_546, z_out_371, z_out_315,
      z_out_327, z_out_848, (MultLoop_acc_1587_nl), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_543 = (AccumDotWidth_mux1h_1192_nl) + (AccumDotWidth_mux1h_1193_nl);
  assign z_out_543 = nl_z_out_543[21:0];
  assign nl_AccumDotWidth_acc_2581_nl = conv_s2s_21_22(z_out_1045_29_7[22:2]) + conv_s2s_21_22(z_out_857_29_7[22:2]);
  assign AccumDotWidth_acc_2581_nl = nl_AccumDotWidth_acc_2581_nl[21:0];
  assign MultLoop_mux1h_501_nl = MUX1HOT_v_22_4_2(z_out_161_28_7, (AccumDotWidth_acc_2581_nl),
      z_out_335, z_out_174_28_7, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2582_nl = conv_s2s_21_22(z_out_1072_29_7[22:2]) + conv_s2s_21_22(z_out_586_29_7[22:2]);
  assign AccumDotWidth_acc_2582_nl = nl_AccumDotWidth_acc_2582_nl[21:0];
  assign nl_AccumDotWidth_acc_2583_nl = conv_s2s_21_22(z_out_994_29_7[22:2]) + conv_s2s_21_22(z_out_599_29_7[22:2]);
  assign AccumDotWidth_acc_2583_nl = nl_AccumDotWidth_acc_2583_nl[21:0];
  assign MultLoop_mux1h_502_nl = MUX1HOT_v_22_4_2(z_out_675_28_7, (AccumDotWidth_acc_2582_nl),
      (AccumDotWidth_acc_2583_nl), z_out_175_28_7, {(fsm_output[2]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_544 = (MultLoop_mux1h_501_nl) + (MultLoop_mux1h_502_nl);
  assign z_out_544 = nl_z_out_544[21:0];
  assign nl_AccumDotWidth_acc_2584_nl = conv_s2s_21_22(z_out_994_29_7[22:2]) + conv_s2s_21_22(z_out_998_29_7[22:2]);
  assign AccumDotWidth_acc_2584_nl = nl_AccumDotWidth_acc_2584_nl[21:0];
  assign AccumDotWidth_mux1h_1194_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2584_nl),
      z_out_411, AccumDotWidth_acc_1378_itm, z_out_712, z_out_408, z_out_376, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2585_nl = conv_s2s_21_22(z_out_1178_29_7[22:2]) + conv_s2s_21_22(z_out_1181_29_7[22:2]);
  assign AccumDotWidth_acc_2585_nl = nl_AccumDotWidth_acc_2585_nl[21:0];
  assign nl_AccumDotWidth_acc_2586_nl = conv_s2s_21_22(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm)
      + conv_s2s_21_22(z_out_924_29_7[22:2]);
  assign AccumDotWidth_acc_2586_nl = nl_AccumDotWidth_acc_2586_nl[21:0];
  assign AccumDotWidth_mux1h_1195_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2585_nl),
      z_out_409, (AccumDotWidth_acc_2586_nl), z_out_721, z_out_405, z_out_373, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_545 = (AccumDotWidth_mux1h_1194_nl) + (AccumDotWidth_mux1h_1195_nl);
  assign z_out_545 = nl_z_out_545[21:0];
  assign nl_AccumDotWidth_acc_2587_nl = conv_s2s_21_22(z_out_1179_29_7[22:2]) + conv_s2s_21_22(z_out_1183_29_7[22:2]);
  assign AccumDotWidth_acc_2587_nl = nl_AccumDotWidth_acc_2587_nl[21:0];
  assign AccumDotWidth_mux1h_1196_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2587_nl),
      AccumDotWidth_acc_1198_itm, z_out_719, z_out_401, AccumDotWidth_acc_1932_itm,
      {(fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) , (fsm_output[6]) ,
      (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2588_nl = conv_s2s_21_22(z_out_1182_29_7[22:2]) + conv_s2s_21_22(z_out_1188_29_9);
  assign AccumDotWidth_acc_2588_nl = nl_AccumDotWidth_acc_2588_nl[21:0];
  assign AccumDotWidth_mux1h_1197_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2588_nl),
      z_out_429, z_out_428, z_out_359, z_out_403, z_out_379, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_546 = (AccumDotWidth_mux1h_1196_nl) + (AccumDotWidth_mux1h_1197_nl);
  assign z_out_546 = nl_z_out_546[21:0];
  assign nl_MultLoop_acc_1594_nl = (z_out_1076_29_7[21:0]) + (z_out_1072_29_7[21:0]);
  assign MultLoop_acc_1594_nl = nl_MultLoop_acc_1594_nl[21:0];
  assign AccumDotWidth_mux1h_1198_nl = MUX1HOT_v_22_7_2(z_out_431, z_out_343, z_out_380,
      z_out_720, z_out_407, z_out_378, (MultLoop_acc_1594_nl), {nnet_relu_layer2_t_layer3_t_relu_config3_for_if_or_1_cse
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1595_nl = (z_out_1071_29_7[21:0]) + (z_out_1070_29_7[21:0]);
  assign MultLoop_acc_1595_nl = nl_MultLoop_acc_1595_nl[21:0];
  assign AccumDotWidth_mux1h_1199_nl = MUX1HOT_v_22_7_2(z_out_424, z_out_399, z_out_430,
      z_out_376, z_out_718, z_out_404, (MultLoop_acc_1595_nl), {AccumDotWidth_or_149_cse
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign nl_z_out_547 = (AccumDotWidth_mux1h_1198_nl) + (AccumDotWidth_mux1h_1199_nl);
  assign z_out_547 = nl_z_out_547[21:0];
  assign nl_AccumDotWidth_acc_2589_nl = conv_s2s_21_22(z_out_1089_29_7[22:2]) + conv_s2s_21_22(z_out_853_29_7[22:2]);
  assign AccumDotWidth_acc_2589_nl = nl_AccumDotWidth_acc_2589_nl[21:0];
  assign MultLoop_mux1h_503_nl = MUX1HOT_v_22_3_2(z_out_151_28_7, (AccumDotWidth_acc_2589_nl),
      z_out_171_28_7, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2590_nl = conv_s2s_21_22(z_out_1176_29_7[22:2]) + conv_s2s_21_22(z_out_864_29_7[22:2]);
  assign AccumDotWidth_acc_2590_nl = nl_AccumDotWidth_acc_2590_nl[21:0];
  assign MultLoop_mux1h_504_nl = MUX1HOT_v_22_3_2(z_out_152_28_7, (AccumDotWidth_acc_2590_nl),
      z_out_173_28_7, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_548 = (MultLoop_mux1h_503_nl) + (MultLoop_mux1h_504_nl);
  assign z_out_548 = nl_z_out_548[21:0];
  assign nl_AccumDotWidth_acc_2591_nl = conv_s2s_21_22(z_out_995_29_7[22:2]) + conv_s2s_21_22(z_out_1000_29_7[22:2]);
  assign AccumDotWidth_acc_2591_nl = nl_AccumDotWidth_acc_2591_nl[21:0];
  assign nl_AccumDotWidth_acc_2592_nl = conv_s2s_21_22(z_out_1181_29_7[22:2]) + conv_s2s_21_22(z_out_856_29_7[22:2]);
  assign AccumDotWidth_acc_2592_nl = nl_AccumDotWidth_acc_2592_nl[21:0];
  assign AccumDotWidth_mux1h_1200_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2591_nl),
      z_out_405, z_out_381, z_out_710, z_out_731, (AccumDotWidth_acc_2592_nl), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2593_nl = conv_s2s_21_22(z_out_1004_29_9) + conv_s2s_21_22(z_out_996_29_7[22:2]);
  assign AccumDotWidth_acc_2593_nl = nl_AccumDotWidth_acc_2593_nl[21:0];
  assign nl_AccumDotWidth_acc_2594_nl = conv_s2s_21_22(z_out_868_29_7[22:2]) + conv_s2s_21_22(z_out_1098_29_7[22:2]);
  assign AccumDotWidth_acc_2594_nl = nl_AccumDotWidth_acc_2594_nl[21:0];
  assign AccumDotWidth_mux1h_1201_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2593_nl),
      z_out_404, z_out_378, z_out_709, z_out_740, (AccumDotWidth_acc_2594_nl), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_549 = (AccumDotWidth_mux1h_1200_nl) + (AccumDotWidth_mux1h_1201_nl);
  assign z_out_549 = nl_z_out_549[21:0];
  assign nl_AccumDotWidth_acc_2595_nl = conv_s2s_21_22(z_out_1155_29_7[22:2]) + conv_s2s_21_22(z_out_940_29_7[22:2]);
  assign AccumDotWidth_acc_2595_nl = nl_AccumDotWidth_acc_2595_nl[21:0];
  assign MultLoop_mux1h_505_nl = MUX1HOT_v_22_3_2(z_out_150_28_7, (AccumDotWidth_acc_2595_nl),
      z_out_172_28_7, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2596_nl = conv_s2s_21_22(z_out_1109_29_7[22:2]) + conv_s2s_21_22(z_out_916_29_7[22:2]);
  assign AccumDotWidth_acc_2596_nl = nl_AccumDotWidth_acc_2596_nl[21:0];
  assign MultLoop_mux1h_506_nl = MUX1HOT_v_22_3_2(z_out_193_28_7, (AccumDotWidth_acc_2596_nl),
      z_out_170_28_7, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_z_out_550 = (MultLoop_mux1h_505_nl) + (MultLoop_mux1h_506_nl);
  assign z_out_550 = nl_z_out_550[21:0];
  assign nl_AccumDotWidth_acc_2597_nl = conv_s2s_21_22(z_out_1123_29_7[22:2]) + conv_s2s_21_22(z_out_1010_29_7[22:2]);
  assign AccumDotWidth_acc_2597_nl = nl_AccumDotWidth_acc_2597_nl[21:0];
  assign AccumDotWidth_mux1h_1202_nl = MUX1HOT_v_22_6_2(z_out_369, (AccumDotWidth_acc_2597_nl),
      z_out_387, z_out_711, z_out_391, z_out_367, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2598_nl = conv_s2s_21_22(z_out_1089_29_7[22:2]) + conv_s2s_21_22(z_out_922_29_7[22:2]);
  assign AccumDotWidth_acc_2598_nl = nl_AccumDotWidth_acc_2598_nl[21:0];
  assign AccumDotWidth_mux1h_1203_nl = MUX1HOT_v_22_6_2(z_out_377, (AccumDotWidth_acc_2598_nl),
      z_out_383, z_out_714, z_out_390, z_out_730, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_551 = (AccumDotWidth_mux1h_1202_nl) + (AccumDotWidth_mux1h_1203_nl);
  assign z_out_551 = nl_z_out_551[21:0];
  assign nl_AccumDotWidth_acc_2599_nl = conv_s2s_21_22(z_out_957_29_7[22:2]) + conv_s2s_21_22(z_out_597_29_7[22:2]);
  assign AccumDotWidth_acc_2599_nl = nl_AccumDotWidth_acc_2599_nl[21:0];
  assign nl_AccumDotWidth_acc_2600_nl = conv_s2s_21_22(z_out_957_29_7[22:2]) + conv_s2s_21_22(z_out_1113_29_7[22:2]);
  assign AccumDotWidth_acc_2600_nl = nl_AccumDotWidth_acc_2600_nl[21:0];
  assign nl_AccumDotWidth_acc_2601_nl = conv_s2s_21_22(z_out_1014_29_7[22:2]) + conv_s2s_21_22(z_out_617_29_7[22:2]);
  assign AccumDotWidth_acc_2601_nl = nl_AccumDotWidth_acc_2601_nl[21:0];
  assign nl_AccumDotWidth_acc_2602_nl = conv_s2s_21_22(z_out_990_29_7[22:2]) + conv_s2s_21_22(z_out_973_29_7[22:2]);
  assign AccumDotWidth_acc_2602_nl = nl_AccumDotWidth_acc_2602_nl[21:0];
  assign nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[607:600]));
  assign MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1204_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2599_nl),
      (AccumDotWidth_acc_2600_nl), (AccumDotWidth_acc_2601_nl), (AccumDotWidth_acc_2602_nl),
      (readslicef_29_22_7((MultLoop_76_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2603_nl = conv_s2s_21_22(z_out_1121_29_7[22:2]) + conv_s2s_21_22(z_out_921_29_7[22:2]);
  assign AccumDotWidth_acc_2603_nl = nl_AccumDotWidth_acc_2603_nl[21:0];
  assign nl_AccumDotWidth_acc_2604_nl = conv_s2s_21_22(z_out_1150_29_7[22:2]) + conv_s2s_21_22(z_out_1135_29_9);
  assign AccumDotWidth_acc_2604_nl = nl_AccumDotWidth_acc_2604_nl[21:0];
  assign nl_AccumDotWidth_acc_2605_nl = conv_s2s_21_22(z_out_885_29_7[22:2]) + conv_s2s_21_22(z_out_1026_29_7[22:2]);
  assign AccumDotWidth_acc_2605_nl = nl_AccumDotWidth_acc_2605_nl[21:0];
  assign nl_AccumDotWidth_acc_2606_nl = conv_s2s_21_22(z_out_997_29_7[22:2]) + conv_s2s_21_22(z_out_600_29_7[22:2]);
  assign AccumDotWidth_acc_2606_nl = nl_AccumDotWidth_acc_2606_nl[21:0];
  assign nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[615:608]));
  assign MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1205_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2603_nl),
      (AccumDotWidth_acc_2604_nl), (AccumDotWidth_acc_2605_nl), (AccumDotWidth_acc_2606_nl),
      (readslicef_29_22_7((MultLoop_77_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_552 = (AccumDotWidth_mux1h_1204_nl) + (AccumDotWidth_mux1h_1205_nl);
  assign z_out_552 = nl_z_out_552[21:0];
  assign nl_AccumDotWidth_acc_2607_nl = conv_s2s_21_22(z_out_1005_29_7[22:2]) + conv_s2s_21_22(z_out_1072_29_7[22:2]);
  assign AccumDotWidth_acc_2607_nl = nl_AccumDotWidth_acc_2607_nl[21:0];
  assign nl_AccumDotWidth_acc_2608_nl = conv_s2s_21_22(z_out_956_29_7[22:2]) + conv_s2s_21_22(z_out_1112_29_7[22:2]);
  assign AccumDotWidth_acc_2608_nl = nl_AccumDotWidth_acc_2608_nl[21:0];
  assign nl_AccumDotWidth_acc_2609_nl = conv_s2s_21_22(z_out_1019_29_7[22:2]) + conv_s2s_21_22(z_out_856_29_7[22:2]);
  assign AccumDotWidth_acc_2609_nl = nl_AccumDotWidth_acc_2609_nl[21:0];
  assign nl_AccumDotWidth_acc_2610_nl = conv_s2s_21_22(z_out_892_29_7[22:2]) + conv_s2s_21_22(z_out_579_29_7[22:2]);
  assign AccumDotWidth_acc_2610_nl = nl_AccumDotWidth_acc_2610_nl[21:0];
  assign nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[623:616]));
  assign MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1206_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2607_nl),
      (AccumDotWidth_acc_2608_nl), (AccumDotWidth_acc_2609_nl), (AccumDotWidth_acc_2610_nl),
      (readslicef_29_22_7((MultLoop_78_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2611_nl = conv_s2s_21_22(z_out_594_29_7[22:2]) + conv_s2s_21_22(z_out_1080_29_7[22:2]);
  assign AccumDotWidth_acc_2611_nl = nl_AccumDotWidth_acc_2611_nl[21:0];
  assign nl_AccumDotWidth_acc_2612_nl = conv_s2s_21_22(z_out_1149_29_7[22:2]) + conv_s2s_21_22(z_out_980_29_7[22:2]);
  assign AccumDotWidth_acc_2612_nl = nl_AccumDotWidth_acc_2612_nl[21:0];
  assign nl_AccumDotWidth_acc_2613_nl = conv_s2s_21_22(z_out_1079_29_7[22:2]) + conv_s2s_21_22(z_out_594_29_7[22:2]);
  assign AccumDotWidth_acc_2613_nl = nl_AccumDotWidth_acc_2613_nl[21:0];
  assign nl_AccumDotWidth_acc_2614_nl = conv_s2s_21_22(z_out_956_29_7[22:2]) + conv_s2s_21_22(z_out_984_29_7[22:2]);
  assign AccumDotWidth_acc_2614_nl = nl_AccumDotWidth_acc_2614_nl[21:0];
  assign nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[631:624]));
  assign MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1207_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2611_nl),
      (AccumDotWidth_acc_2612_nl), (AccumDotWidth_acc_2613_nl), (AccumDotWidth_acc_2614_nl),
      (readslicef_29_22_7((MultLoop_79_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_553 = (AccumDotWidth_mux1h_1206_nl) + (AccumDotWidth_mux1h_1207_nl);
  assign z_out_553 = nl_z_out_553[21:0];
  assign nl_AccumDotWidth_acc_2615_nl = conv_s2s_21_22(z_out_894_29_7[22:2]) + conv_s2s_21_22(z_out_1099_29_7[22:2]);
  assign AccumDotWidth_acc_2615_nl = nl_AccumDotWidth_acc_2615_nl[21:0];
  assign nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_3_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[351:344]));
  assign MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1208_nl = MUX1HOT_v_22_5_2(z_out_746, z_out_722, (AccumDotWidth_acc_2615_nl),
      z_out_394, (readslicef_29_22_7((MultLoop_44_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2616_nl = conv_s2s_21_22(z_out_937_29_7[22:2]) + conv_s2s_21_22(z_out_1185_29_7[22:2]);
  assign AccumDotWidth_acc_2616_nl = nl_AccumDotWidth_acc_2616_nl[21:0];
  assign nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_45_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[359:352]));
  assign MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1209_nl = MUX1HOT_v_22_5_2(z_out_743, z_out_713, (AccumDotWidth_acc_2616_nl),
      z_out_392, (readslicef_29_22_7((MultLoop_45_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_554 = (AccumDotWidth_mux1h_1208_nl) + (AccumDotWidth_mux1h_1209_nl);
  assign z_out_554 = nl_z_out_554[21:0];
  assign nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[639:632]));
  assign MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1210_nl = MUX1HOT_v_22_5_2(z_out_742, z_out_745, z_out_398,
      z_out_370, (readslicef_29_22_7((MultLoop_80_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[647:640]));
  assign MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign AccumDotWidth_mux1h_1211_nl = MUX1HOT_v_22_5_2(z_out_741, z_out_744, z_out_399,
      z_out_362, (readslicef_29_22_7((MultLoop_81_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_555 = (AccumDotWidth_mux1h_1210_nl) + (AccumDotWidth_mux1h_1211_nl);
  assign z_out_555 = nl_z_out_555[21:0];
  assign nl_AccumDotWidth_acc_2617_nl = conv_s2s_21_22(z_out_1128_29_7[22:2]) + conv_s2s_21_22(z_out_1014_29_7[22:2]);
  assign AccumDotWidth_acc_2617_nl = nl_AccumDotWidth_acc_2617_nl[21:0];
  assign AccumDotWidth_mux1h_1212_nl = MUX1HOT_v_22_5_2(z_out_373, (AccumDotWidth_acc_2617_nl),
      z_out_747, z_out_396, z_out_724, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , AccumDotWidth_or_152_cse , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1213_nl = MUX1HOT_v_22_5_2(z_out_374, z_out_408, z_out_746,
      z_out_388, z_out_726, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , AccumDotWidth_or_152_cse , (fsm_output[7])});
  assign nl_z_out_556 = (AccumDotWidth_mux1h_1212_nl) + (AccumDotWidth_mux1h_1213_nl);
  assign z_out_556 = nl_z_out_556[21:0];
  assign nl_AccumDotWidth_acc_2618_nl = conv_s2s_21_22(z_out_913_29_7[22:2]) + conv_s2s_21_22(z_out_865_29_7[22:2]);
  assign AccumDotWidth_acc_2618_nl = nl_AccumDotWidth_acc_2618_nl[21:0];
  assign AccumDotWidth_mux1h_1214_nl = MUX1HOT_v_22_6_2(z_out_378, z_out_398, (AccumDotWidth_acc_2618_nl),
      z_out_370, z_out_389, z_out_727, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2619_nl = conv_s2s_21_22(z_out_1000_29_7[22:2]) + conv_s2s_21_22(z_out_900_29_7[22:2]);
  assign AccumDotWidth_acc_2619_nl = nl_AccumDotWidth_acc_2619_nl[21:0];
  assign AccumDotWidth_mux1h_1215_nl = MUX1HOT_v_22_6_2(z_out_375, z_out_399, (AccumDotWidth_acc_2619_nl),
      z_out_367, z_out_392, z_out_722, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_557 = (AccumDotWidth_mux1h_1214_nl) + (AccumDotWidth_mux1h_1215_nl);
  assign z_out_557 = nl_z_out_557[21:0];
  assign AccumDotWidth_mux1h_1216_nl = MUX1HOT_v_22_6_2(z_out_380, z_out_406, z_out_386,
      z_out_702, z_out_395, z_out_731, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1217_nl = MUX1HOT_v_22_6_2(z_out_376, z_out_410, z_out_388,
      z_out_715, z_out_386, z_out_725, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_558 = (AccumDotWidth_mux1h_1216_nl) + (AccumDotWidth_mux1h_1217_nl);
  assign z_out_558 = nl_z_out_558[21:0];
  assign nl_MultLoop_acc_1596_nl = ({MultLoop_acc_1280_psp , (MultLoop_acc_88_itm[10:0])})
      + (z_out_577_29_7[21:0]);
  assign MultLoop_acc_1596_nl = nl_MultLoop_acc_1596_nl[21:0];
  assign AccumDotWidth_mux1h_1218_nl = MUX1HOT_v_22_7_2(z_out_749, z_out_309, z_out_392,
      z_out_365, z_out_733, z_out_729, (MultLoop_acc_1596_nl), {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1597_nl = (z_out_583_29_7[21:0]) + (z_out_575_29_7[21:0]);
  assign MultLoop_acc_1597_nl = nl_MultLoop_acc_1597_nl[21:0];
  assign AccumDotWidth_mux1h_1219_nl = MUX1HOT_v_22_7_2(z_out_745, AccumDotWidth_acc_1397_itm,
      z_out_391, z_out_368, z_out_725, z_out_728, (MultLoop_acc_1597_nl), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_559 = (AccumDotWidth_mux1h_1218_nl) + (AccumDotWidth_mux1h_1219_nl);
  assign z_out_559 = nl_z_out_559[21:0];
  assign AccumDotWidth_mux1h_1220_nl = MUX1HOT_v_22_6_2(z_out_741, z_out_494, z_out_694,
      z_out_366, z_out_399, z_out_713, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1221_nl = MUX1HOT_v_22_6_2(z_out_740, AccumDotWidth_acc_1371_itm,
      z_out_695, z_out_362, z_out_398, z_out_723, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_560 = (AccumDotWidth_mux1h_1220_nl) + (AccumDotWidth_mux1h_1221_nl);
  assign z_out_560 = nl_z_out_560[21:0];
  assign nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[767:760]));
  assign MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign MultLoop_mux_97_nl = MUX_v_22_2_2(z_out_162_28_7, (readslicef_29_22_7((MultLoop_96_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl))),
      fsm_output[8]);
  assign MultLoop_mux_98_nl = MUX_v_22_2_2(z_out_149_28_7, z_out_152_28_7, fsm_output[8]);
  assign nl_z_out_561 = (MultLoop_mux_97_nl) + (MultLoop_mux_98_nl);
  assign z_out_561 = nl_z_out_561[21:0];
  assign nl_MultLoop_acc_1599_nl = (z_out_1162_29_7[21:11]) + conv_s2s_8_11(InitAccum_io_read_b4_rsc_cse_sva[71:64]);
  assign MultLoop_acc_1599_nl = nl_MultLoop_acc_1599_nl[10:0];
  assign nl_MultLoop_acc_1598_nl = ({(MultLoop_acc_1599_nl) , (z_out_1162_29_7[10:0])})
      + (z_out_862_29_7[21:0]);
  assign MultLoop_acc_1598_nl = nl_MultLoop_acc_1598_nl[21:0];
  assign AccumDotWidth_mux1h_1222_nl = MUX1HOT_v_22_6_2(z_out_329, z_out_253, z_out_525,
      z_out_371, z_out_316, (MultLoop_acc_1598_nl), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1600_nl = (z_out_861_29_7[21:0]) + (z_out_857_29_7[21:0]);
  assign MultLoop_acc_1600_nl = nl_MultLoop_acc_1600_nl[21:0];
  assign AccumDotWidth_mux1h_1223_nl = MUX1HOT_v_22_6_2(z_out_344, z_out_685, z_out_350,
      z_out_374, z_out_308, (MultLoop_acc_1600_nl), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_562 = (AccumDotWidth_mux1h_1222_nl) + (AccumDotWidth_mux1h_1223_nl);
  assign z_out_562 = nl_z_out_562[21:0];
  assign nl_AccumDotWidth_acc_2625_nl = (z_out_891_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[63:56]);
  assign AccumDotWidth_acc_2625_nl = nl_AccumDotWidth_acc_2625_nl[9:0];
  assign nl_AccumDotWidth_acc_2620_nl = conv_s2s_21_22({(AccumDotWidth_acc_2625_nl)
      , (z_out_891_29_7[12:2])}) + conv_s2s_21_22(z_out_583_29_7[22:2]) + conv_s2s_21_22(z_out_1088_29_7[22:2])
      + conv_s2s_21_22(z_out_1089_29_7[22:2]) + conv_s2s_21_22(z_out_1080_29_7[22:2])
      + conv_s2s_21_22(z_out_585_29_7[22:2]);
  assign AccumDotWidth_acc_2620_nl = nl_AccumDotWidth_acc_2620_nl[21:0];
  assign nl_AccumDotWidth_acc_2629_nl = (z_out_907_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2629_nl = nl_AccumDotWidth_acc_2629_nl[9:0];
  assign nl_AccumDotWidth_acc_2627_nl = conv_s2s_21_22({(AccumDotWidth_acc_2629_nl)
      , (z_out_907_29_7[12:2])}) + conv_s2s_21_22(z_out_986_29_7[22:2]) + conv_s2s_21_22(z_out_1039_29_7[22:2]);
  assign AccumDotWidth_acc_2627_nl = nl_AccumDotWidth_acc_2627_nl[21:0];
  assign nl_AccumDotWidth_acc_2626_nl = z_out_552 + (AccumDotWidth_acc_2627_nl);
  assign AccumDotWidth_acc_2626_nl = nl_AccumDotWidth_acc_2626_nl[21:0];
  assign nl_MultLoop_acc_1602_nl = (z_out_1161_29_7[21:11]) + conv_s2s_8_11(InitAccum_io_read_b4_rsc_cse_sva[63:56]);
  assign MultLoop_acc_1602_nl = nl_MultLoop_acc_1602_nl[10:0];
  assign nl_MultLoop_acc_1601_nl = ({(MultLoop_acc_1602_nl) , (z_out_1161_29_7[10:0])})
      + (z_out_923_29_7[21:0]);
  assign MultLoop_acc_1601_nl = nl_MultLoop_acc_1601_nl[21:0];
  assign AccumDotWidth_mux1h_1224_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2620_nl),
      z_out_520, z_out_258, AccumDotWidth_acc_1274_itm, (AccumDotWidth_acc_2626_nl),
      z_out_400, (MultLoop_acc_1601_nl), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1225_nl = MUX1HOT_v_22_8_2(z_out_559, AccumDotWidth_acc_1169_itm,
      z_out_681, z_out_309, z_out_244, z_out_423, z_out_558, z_out_807, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_563 = (AccumDotWidth_mux1h_1224_nl) + (AccumDotWidth_mux1h_1225_nl);
  assign z_out_563 = nl_z_out_563[21:0];
  assign nl_AccumDotWidth_acc_2635_nl = (z_out_877_29_7[22:13]) + conv_s2s_8_10(b2_rsci_idat_mxwt[15:8]);
  assign AccumDotWidth_acc_2635_nl = nl_AccumDotWidth_acc_2635_nl[9:0];
  assign nl_AccumDotWidth_acc_2630_nl = conv_s2s_21_22({(AccumDotWidth_acc_2635_nl)
      , (z_out_877_29_7[12:2])}) + conv_s2s_21_22(z_out_983_29_7[22:2]) + conv_s2s_21_22(z_out_1008_29_7[22:2])
      + conv_s2s_21_22(z_out_1083_29_7[22:2]) + conv_s2s_21_22(z_out_1086_29_7[22:2])
      + conv_s2s_21_22(z_out_1084_29_7[22:2]);
  assign AccumDotWidth_acc_2630_nl = nl_AccumDotWidth_acc_2630_nl[21:0];
  assign nl_AccumDotWidth_acc_2636_nl = z_out_550 + z_out_548;
  assign AccumDotWidth_acc_2636_nl = nl_AccumDotWidth_acc_2636_nl[21:0];
  assign nl_AccumDotWidth_acc_2637_nl = conv_s2s_21_22(z_out_964_29_7[22:2]) + conv_s2s_21_22(z_out_912_29_7[22:2])
      + conv_s2s_21_22(z_out_999_29_7[22:2]) + conv_s2s_21_22(z_out_1116_29_7[22:2]);
  assign AccumDotWidth_acc_2637_nl = nl_AccumDotWidth_acc_2637_nl[21:0];
  assign nl_AccumDotWidth_acc_2645_nl = (z_out_877_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2645_nl = nl_AccumDotWidth_acc_2645_nl[9:0];
  assign nl_AccumDotWidth_acc_2640_nl = conv_s2s_21_22({(AccumDotWidth_acc_2645_nl)
      , (z_out_877_29_7[12:2])}) + conv_s2s_21_22(z_out_948_29_7[22:2]) + conv_s2s_21_22(z_out_627_29_7[22:2])
      + conv_s2s_21_22(z_out_905_29_7[22:2]) + conv_s2s_21_22(z_out_594_29_7[22:2])
      + conv_s2s_21_22(z_out_613_29_7[22:2]);
  assign AccumDotWidth_acc_2640_nl = nl_AccumDotWidth_acc_2640_nl[21:0];
  assign nl_MultLoop_acc_1604_nl = (z_out_1160_29_7[21:11]) + conv_s2s_8_11(InitAccum_io_read_b4_rsc_cse_sva[55:48]);
  assign MultLoop_acc_1604_nl = nl_MultLoop_acc_1604_nl[10:0];
  assign nl_MultLoop_acc_1603_nl = ({(MultLoop_acc_1604_nl) , (z_out_1160_29_7[10:0])})
      + (z_out_986_29_7[21:0]);
  assign MultLoop_acc_1603_nl = nl_MultLoop_acc_1603_nl[21:0];
  assign AccumDotWidth_mux1h_1226_nl = MUX1HOT_v_22_8_2((AccumDotWidth_acc_2630_nl),
      z_out_244, z_out_527, z_out_258, (AccumDotWidth_acc_2636_nl), (AccumDotWidth_acc_2637_nl),
      (AccumDotWidth_acc_2640_nl), (MultLoop_acc_1603_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2646_nl = z_out_525 + z_out_544;
  assign AccumDotWidth_acc_2646_nl = nl_AccumDotWidth_acc_2646_nl[21:0];
  assign nl_AccumDotWidth_acc_2647_nl = conv_s2s_21_22(z_out_1072_29_7[22:2]) + conv_s2s_21_22(z_out_856_29_7[22:2])
      + conv_s2s_21_22(z_out_884_29_7[22:2]) + conv_s2s_21_22(z_out_1032_29_9);
  assign AccumDotWidth_acc_2647_nl = nl_AccumDotWidth_acc_2647_nl[21:0];
  assign AccumDotWidth_mux1h_1227_nl = MUX1HOT_v_22_8_2(z_out_558, AccumDotWidth_acc_1218_itm,
      z_out_525, z_out_247, (AccumDotWidth_acc_2646_nl), (AccumDotWidth_acc_2647_nl),
      z_out_849, z_out_309, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_564 = (AccumDotWidth_mux1h_1226_nl) + (AccumDotWidth_mux1h_1227_nl);
  assign z_out_564 = nl_z_out_564[21:0];
  assign nl_MultLoop_acc_1606_nl = (z_out_664_28_7[21:11]) + conv_s2s_8_11(InitAccum_io_read_b4_rsc_cse_sva[7:0]);
  assign MultLoop_acc_1606_nl = nl_MultLoop_acc_1606_nl[10:0];
  assign nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[7:0]));
  assign MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1605_nl = ({(MultLoop_acc_1606_nl) , (z_out_664_28_7[10:0])})
      + (readslicef_29_22_7((MultLoop_1_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1605_nl = nl_MultLoop_acc_1605_nl[21:0];
  assign AccumDotWidth_mux1h_1228_nl = MUX1HOT_v_22_7_2(z_out_372, z_out_235, z_out_251,
      z_out_257, z_out_850, z_out_259, (MultLoop_acc_1605_nl), {(fsm_output[1]) ,
      (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) , (fsm_output[6]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[15:8]));
  assign MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[23:16]));
  assign MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1607_nl = (readslicef_29_22_7((MultLoop_2_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + (readslicef_29_22_7((MultLoop_3_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1607_nl = nl_MultLoop_acc_1607_nl[21:0];
  assign AccumDotWidth_mux1h_1229_nl = MUX1HOT_v_22_8_2(z_out_371, AccumDotWidth_acc_1235_itm,
      z_out_256, z_out_257, z_out_260, z_out_848, z_out_310, (MultLoop_acc_1607_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_565 = (AccumDotWidth_mux1h_1228_nl) + (AccumDotWidth_mux1h_1229_nl);
  assign z_out_565 = nl_z_out_565[21:0];
  assign nl_AccumDotWidth_acc_2655_nl = (z_out_1065_29_9[20:11]) + conv_s2s_8_10(b2_rsci_idat_mxwt[47:40]);
  assign AccumDotWidth_acc_2655_nl = nl_AccumDotWidth_acc_2655_nl[9:0];
  assign nl_AccumDotWidth_acc_2650_nl = conv_s2s_21_22({(AccumDotWidth_acc_2655_nl)
      , (z_out_1065_29_9[10:0])}) + conv_s2s_21_22(z_out_925_29_7[22:2]) + conv_s2s_21_22(z_out_607_29_7[22:2])
      + conv_s2s_21_22(z_out_609_29_7[22:2]) + conv_s2s_21_22(z_out_614_29_7[22:2])
      + conv_s2s_21_22(z_out_616_29_7[22:2]);
  assign AccumDotWidth_acc_2650_nl = nl_AccumDotWidth_acc_2650_nl[21:0];
  assign nl_AccumDotWidth_acc_2660_nl = conv_s2s_21_22(z_out_1088_29_7[22:2]) + conv_s2s_21_22(z_out_860_29_7[22:2])
      + conv_s2s_21_22(z_out_1003_29_9) + conv_s2s_21_22(z_out_611_29_7[22:2]);
  assign AccumDotWidth_acc_2660_nl = nl_AccumDotWidth_acc_2660_nl[21:0];
  assign nl_AccumDotWidth_acc_2656_nl = (AccumDotWidth_acc_2660_nl) + conv_s2s_21_22(z_out_1154_29_7[22:2])
      + conv_s2s_21_22(z_out_947_29_7[22:2]) + conv_s2s_21_22(z_out_1135_29_9) +
      conv_s2s_21_22(z_out_1170_29_7[22:2]);
  assign AccumDotWidth_acc_2656_nl = nl_AccumDotWidth_acc_2656_nl[21:0];
  assign nl_AccumDotWidth_acc_2668_nl = (z_out_1156_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2668_nl = nl_AccumDotWidth_acc_2668_nl[9:0];
  assign nl_AccumDotWidth_acc_2663_nl = conv_s2s_21_22({(AccumDotWidth_acc_2668_nl)
      , (z_out_1156_29_7[12:2])}) + conv_s2s_21_22(z_out_1102_29_7[22:2]) + conv_s2s_21_22(z_out_622_29_7[22:2])
      + conv_s2s_21_22(z_out_1119_29_7[22:2]) + conv_s2s_21_22(z_out_585_29_7[22:2])
      + conv_s2s_21_22(z_out_610_29_7[22:2]);
  assign AccumDotWidth_acc_2663_nl = nl_AccumDotWidth_acc_2663_nl[21:0];
  assign AccumDotWidth_mux1h_1230_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2650_nl),
      z_out_245, z_out_249, (AccumDotWidth_acc_2656_nl), z_out_849, (AccumDotWidth_acc_2663_nl),
      z_out_851, {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2673_nl = conv_s2s_21_22(z_out_1035_29_7[22:2]) + conv_s2s_21_22(z_out_1114_29_7[22:2])
      + conv_s2s_21_22(z_out_1078_29_7[22:2]) + conv_s2s_21_22(z_out_589_29_7[22:2]);
  assign AccumDotWidth_acc_2673_nl = nl_AccumDotWidth_acc_2673_nl[21:0];
  assign nl_AccumDotWidth_acc_2669_nl = (AccumDotWidth_acc_2673_nl) + conv_s2s_21_22(z_out_630_29_7[22:2])
      + conv_s2s_21_22(z_out_970_29_7[22:2]) + conv_s2s_21_22(z_out_917_29_7[22:2])
      + conv_s2s_21_22(z_out_1136_29_9);
  assign AccumDotWidth_acc_2669_nl = nl_AccumDotWidth_acc_2669_nl[21:0];
  assign nl_MultLoop_acc_1608_nl = (z_out_576_29_7[21:0]) + MultLoop_1107_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1608_nl = nl_MultLoop_acc_1608_nl[21:0];
  assign AccumDotWidth_mux1h_1231_nl = MUX1HOT_v_22_8_2(z_out_807, AccumDotWidth_acc_1201_itm,
      z_out_247, z_out_328, (AccumDotWidth_acc_2669_nl), z_out_335, z_out_545, (MultLoop_acc_1608_nl),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_566 = (AccumDotWidth_mux1h_1230_nl) + (AccumDotWidth_mux1h_1231_nl);
  assign z_out_566 = nl_z_out_566[21:0];
  assign nl_AccumDotWidth_acc_2676_nl = conv_s2s_21_22(z_out_1010_29_7[22:2]) + conv_s2s_21_22(z_out_607_29_7[22:2]);
  assign AccumDotWidth_acc_2676_nl = nl_AccumDotWidth_acc_2676_nl[21:0];
  assign AccumDotWidth_mux1h_1232_nl = MUX1HOT_v_22_5_2(z_out_379, z_out_700, z_out_690,
      (AccumDotWidth_acc_2676_nl), z_out_736, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_AccumDotWidth_acc_2677_nl = conv_s2s_21_22(z_out_882_29_7[22:2]) + conv_s2s_21_22(z_out_1022_29_7[22:2]);
  assign AccumDotWidth_acc_2677_nl = nl_AccumDotWidth_acc_2677_nl[21:0];
  assign AccumDotWidth_mux1h_1233_nl = MUX1HOT_v_22_5_2(z_out_743, z_out_699, z_out_712,
      (AccumDotWidth_acc_2677_nl), z_out_369, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_z_out_567 = (AccumDotWidth_mux1h_1232_nl) + (AccumDotWidth_mux1h_1233_nl);
  assign z_out_567 = nl_z_out_567[21:0];
  assign ConvFiltWidth_else_mux1h_805_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (w2_rsci_idat_mxwt[1071:1064]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (MultLoop_io_read_w4_rsc_cse_sva[1503:1496]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_806_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_160_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_805_nl)) *
      $signed((ConvFiltWidth_else_mux1h_806_nl)));
  assign z_out_568_29_7 = readslicef_30_23_7((mul_160_nl));
  assign ConvFiltWidth_else_mux1h_807_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]), (MultLoop_io_read_w4_rsc_cse_sva[1495:1488]),
      {MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_808_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_46_cse , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_161_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_807_nl)) *
      $signed((ConvFiltWidth_else_mux1h_808_nl)));
  assign z_out_569_29_7 = readslicef_30_23_7((mul_161_nl));
  assign ConvFiltWidth_else_mux1h_809_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]), (MultLoop_io_read_w4_rsc_cse_sva[5895:5888]),
      {(fsm_output[2]) , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_810_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_162_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_809_nl)) *
      $signed((ConvFiltWidth_else_mux1h_810_nl)));
  assign z_out_570_29_7 = readslicef_30_23_7((mul_162_nl));
  assign ConvFiltWidth_else_mux1h_811_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]), (MultLoop_io_read_w4_rsc_cse_sva[1487:1480]),
      {MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_812_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_46_cse , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_163_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_811_nl)) *
      $signed((ConvFiltWidth_else_mux1h_812_nl)));
  assign z_out_571_29_7 = readslicef_30_23_7((mul_163_nl));
  assign ConvFiltWidth_else_mux1h_813_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (MultLoop_io_read_w4_rsc_cse_sva[1479:1472]),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_36_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_164_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_813_nl)) *
      $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_36_nl)));
  assign z_out_572_29_7 = readslicef_30_23_7((mul_164_nl));
  assign ConvFiltWidth_else_mux1h_814_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[39:32]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]), (MultLoop_io_read_w4_rsc_cse_sva[8839:8832]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_815_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_165_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_814_nl)) *
      $signed((ConvFiltWidth_else_mux1h_815_nl)));
  assign z_out_573_29_7 = readslicef_30_23_7((mul_165_nl));
  assign ConvFiltWidth_else_mux1h_816_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]),
      (w2_rsci_idat_mxwt[175:168]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (MultLoop_io_read_w4_rsc_cse_sva[1471:1464]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_817_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_166_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_816_nl)) *
      $signed((ConvFiltWidth_else_mux1h_817_nl)));
  assign z_out_574_29_7 = readslicef_30_23_7((mul_166_nl));
  assign ConvFiltWidth_else_mux1h_818_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (w2_rsci_idat_mxwt[879:872]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (MultLoop_io_read_w4_rsc_cse_sva[1047:1040]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_819_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_167_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_818_nl)) *
      $signed((ConvFiltWidth_else_mux1h_819_nl)));
  assign z_out_575_29_7 = readslicef_30_23_7((mul_167_nl));
  assign ConvFiltWidth_else_mux1h_820_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (w2_rsci_idat_mxwt[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]),
      (MultLoop_io_read_w4_rsc_cse_sva[8847:8840]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_821_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_168_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_820_nl)) *
      $signed((ConvFiltWidth_else_mux1h_821_nl)));
  assign z_out_576_29_7 = readslicef_30_23_7((mul_168_nl));
  assign ConvFiltWidth_else_mux1h_822_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (w2_rsci_idat_mxwt[231:224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]),
      (MultLoop_io_read_w4_rsc_cse_sva[1031:1024]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_823_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_169_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_822_nl)) *
      $signed((ConvFiltWidth_else_mux1h_823_nl)));
  assign z_out_577_29_7 = readslicef_30_23_7((mul_169_nl));
  assign ConvFiltWidth_else_mux1h_824_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[423:416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (MultLoop_io_read_w4_rsc_cse_sva[2711:2704]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_825_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_170_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_824_nl)) *
      $signed((ConvFiltWidth_else_mux1h_825_nl)));
  assign z_out_578_29_7 = readslicef_30_23_7((mul_170_nl));
  assign ConvFiltWidth_else_mux1h_826_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (w2_rsci_idat_mxwt[687:680]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (MultLoop_io_read_w4_rsc_cse_sva[2719:2712]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_827_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_171_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_826_nl)) *
      $signed((ConvFiltWidth_else_mux1h_827_nl)));
  assign z_out_579_29_7 = readslicef_30_23_7((mul_171_nl));
  assign ConvFiltWidth_else_mux1h_828_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (w2_rsci_idat_mxwt[495:488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (MultLoop_io_read_w4_rsc_cse_sva[2695:2688]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_829_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_172_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_828_nl)) *
      $signed((ConvFiltWidth_else_mux1h_829_nl)));
  assign z_out_580_29_7 = readslicef_30_23_7((mul_172_nl));
  assign ConvFiltWidth_else_mux1h_830_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (w2_rsci_idat_mxwt[615:608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (MultLoop_io_read_w4_rsc_cse_sva[2703:2696]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_831_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_173_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_830_nl)) *
      $signed((ConvFiltWidth_else_mux1h_831_nl)));
  assign z_out_581_29_7 = readslicef_30_23_7((mul_173_nl));
  assign ConvFiltWidth_else_mux1h_832_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]), (MultLoop_io_read_w4_rsc_cse_sva[2727:2720]),
      {MultLoop_or_93_cse , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_833_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}), {(fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_174_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_832_nl)) *
      $signed((ConvFiltWidth_else_mux1h_833_nl)));
  assign z_out_582_29_7 = readslicef_30_23_7((mul_174_nl));
  assign ConvFiltWidth_else_mux1h_834_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]),
      (w2_rsci_idat_mxwt[63:56]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]), (MultLoop_io_read_w4_rsc_cse_sva[1039:1032]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_835_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[549:528]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_175_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_834_nl)) *
      $signed((ConvFiltWidth_else_mux1h_835_nl)));
  assign z_out_583_29_7 = readslicef_30_23_7((mul_175_nl));
  assign ConvFiltWidth_else_mux1h_836_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[71:64]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (MultLoop_io_read_w4_rsc_cse_sva[2735:2728]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_837_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}), {(fsm_output[1]) , (fsm_output[2])
      , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_176_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_836_nl)) *
      $signed((ConvFiltWidth_else_mux1h_837_nl)));
  assign z_out_584_29_7 = readslicef_30_23_7((mul_176_nl));
  assign ConvFiltWidth_else_mux1h_838_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (w2_rsci_idat_mxwt[959:952]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]), (MultLoop_io_read_w4_rsc_cse_sva[2743:2736]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_839_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[8])});
  assign mul_177_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_838_nl)) *
      $signed((ConvFiltWidth_else_mux1h_839_nl)));
  assign z_out_585_29_7 = readslicef_30_23_7((mul_177_nl));
  assign ConvFiltWidth_else_mux1h_840_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (w2_rsci_idat_mxwt[135:128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]),
      (MultLoop_io_read_w4_rsc_cse_sva[2751:2744]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_841_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , (fsm_output[8])});
  assign mul_178_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_840_nl)) *
      $signed((ConvFiltWidth_else_mux1h_841_nl)));
  assign z_out_586_29_7 = readslicef_30_23_7((mul_178_nl));
  assign ConvFiltWidth_else_mux1h_842_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (w2_rsci_idat_mxwt[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]), (MultLoop_io_read_w4_rsc_cse_sva[2759:2752]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_843_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_179_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_842_nl)) *
      $signed((ConvFiltWidth_else_mux1h_843_nl)));
  assign z_out_587_29_7 = readslicef_30_23_7((mul_179_nl));
  assign ConvFiltWidth_else_mux1h_844_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (w2_rsci_idat_mxwt[263:256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (MultLoop_io_read_w4_rsc_cse_sva[2767:2760]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_845_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_180_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_844_nl)) *
      $signed((ConvFiltWidth_else_mux1h_845_nl)));
  assign z_out_588_29_7 = readslicef_30_23_7((mul_180_nl));
  assign ConvFiltWidth_else_mux1h_846_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[71:64]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (MultLoop_io_read_w4_rsc_cse_sva[2775:2768]), {(fsm_output[1]) , MultLoop_or_22_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_847_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_181_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_846_nl)) *
      $signed((ConvFiltWidth_else_mux1h_847_nl)));
  assign z_out_589_29_7 = readslicef_30_23_7((mul_181_nl));
  assign ConvFiltWidth_else_mux1h_848_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]),
      (w2_rsci_idat_mxwt[1031:1024]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]),
      (MultLoop_io_read_w4_rsc_cse_sva[4703:4696]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_849_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_182_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_848_nl)) *
      $signed((ConvFiltWidth_else_mux1h_849_nl)));
  assign z_out_590_29_7 = readslicef_30_23_7((mul_182_nl));
  assign ConvFiltWidth_else_mux1h_850_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (w2_rsci_idat_mxwt[255:248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]),
      (MultLoop_io_read_w4_rsc_cse_sva[4711:4704]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_851_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_183_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_850_nl)) *
      $signed((ConvFiltWidth_else_mux1h_851_nl)));
  assign z_out_591_29_7 = readslicef_30_23_7((mul_183_nl));
  assign ConvFiltWidth_else_mux1h_852_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (MultLoop_io_read_w4_rsc_cse_sva[4719:4712]), {(fsm_output[1]) , MultLoop_or_22_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_853_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_184_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_852_nl)) *
      $signed((ConvFiltWidth_else_mux1h_853_nl)));
  assign z_out_592_29_7 = readslicef_30_23_7((mul_184_nl));
  assign ConvFiltWidth_else_mux1h_854_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (w2_rsci_idat_mxwt[647:640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (MultLoop_io_read_w4_rsc_cse_sva[4631:4624]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_855_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_185_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_854_nl)) *
      $signed((ConvFiltWidth_else_mux1h_855_nl)));
  assign z_out_593_29_7 = readslicef_30_23_7((mul_185_nl));
  assign ConvFiltWidth_else_mux1h_856_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[455:448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]), (MultLoop_io_read_w4_rsc_cse_sva[4727:4720]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_857_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_186_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_856_nl)) *
      $signed((ConvFiltWidth_else_mux1h_857_nl)));
  assign z_out_594_29_7 = readslicef_30_23_7((mul_186_nl));
  assign ConvFiltWidth_else_or_730_cse = (fsm_output[6:3]!=4'b0000);
  assign ConvFiltWidth_else_mux1h_858_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]), (w2_rsci_idat_mxwt[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]),
      (MultLoop_io_read_w4_rsc_cse_sva[4735:4728]), {(fsm_output[3]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_859_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (input_1_rsci_idat_mxwt[1033:1012]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_730_cse , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[1]) , (fsm_output[8])});
  assign mul_187_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_858_nl)) *
      $signed((ConvFiltWidth_else_mux1h_859_nl)));
  assign z_out_595_29_7 = readslicef_30_23_7((mul_187_nl));
  assign ConvFiltWidth_else_mux1h_860_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (w2_rsci_idat_mxwt[135:128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (MultLoop_io_read_w4_rsc_cse_sva[4743:4736]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_861_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_188_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_860_nl)) *
      $signed((ConvFiltWidth_else_mux1h_861_nl)));
  assign z_out_596_29_7 = readslicef_30_23_7((mul_188_nl));
  assign ConvFiltWidth_else_mux1h_862_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]),
      (w2_rsci_idat_mxwt[335:328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]),
      (MultLoop_io_read_w4_rsc_cse_sva[4751:4744]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_863_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_189_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_862_nl)) *
      $signed((ConvFiltWidth_else_mux1h_863_nl)));
  assign z_out_597_29_7 = readslicef_30_23_7((mul_189_nl));
  assign ConvFiltWidth_else_mux1h_864_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]),
      (w2_rsci_idat_mxwt[647:640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (MultLoop_io_read_w4_rsc_cse_sva[4623:4616]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_865_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , AccumDotWidth_or_38_cse , (fsm_output[8])});
  assign mul_190_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_864_nl)) *
      $signed((ConvFiltWidth_else_mux1h_865_nl)));
  assign z_out_598_29_7 = readslicef_30_23_7((mul_190_nl));
  assign ConvFiltWidth_else_mux1h_866_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (w2_rsci_idat_mxwt[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (MultLoop_io_read_w4_rsc_cse_sva[4759:4752]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_867_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_191_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_866_nl)) *
      $signed((ConvFiltWidth_else_mux1h_867_nl)));
  assign z_out_599_29_7 = readslicef_30_23_7((mul_191_nl));
  assign ConvFiltWidth_else_mux1h_868_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]),
      (w2_rsci_idat_mxwt[263:256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]),
      (MultLoop_io_read_w4_rsc_cse_sva[4767:4760]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_869_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_192_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_868_nl)) *
      $signed((ConvFiltWidth_else_mux1h_869_nl)));
  assign z_out_600_29_7 = readslicef_30_23_7((mul_192_nl));
  assign ConvFiltWidth_else_mux1h_870_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]),
      (w2_rsci_idat_mxwt[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (MultLoop_io_read_w4_rsc_cse_sva[2511:2504]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_871_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_193_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_870_nl)) *
      $signed((ConvFiltWidth_else_mux1h_871_nl)));
  assign z_out_601_29_7 = readslicef_30_23_7((mul_193_nl));
  assign ConvFiltWidth_else_mux1h_872_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]), (MultLoop_io_read_w4_rsc_cse_sva[2519:2512]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_873_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[8])});
  assign mul_194_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_872_nl)) *
      $signed((ConvFiltWidth_else_mux1h_873_nl)));
  assign z_out_602_29_7 = readslicef_30_23_7((mul_194_nl));
  assign ConvFiltWidth_else_mux1h_874_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[143:136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]),
      (MultLoop_io_read_w4_rsc_cse_sva[2527:2520]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_875_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_195_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_874_nl)) *
      $signed((ConvFiltWidth_else_mux1h_875_nl)));
  assign z_out_603_29_7 = readslicef_30_23_7((mul_195_nl));
  assign ConvFiltWidth_else_mux1h_876_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]), (MultLoop_io_read_w4_rsc_cse_sva[2495:2488]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_877_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[8])});
  assign mul_196_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_876_nl)) *
      $signed((ConvFiltWidth_else_mux1h_877_nl)));
  assign z_out_604_29_7 = readslicef_30_23_7((mul_196_nl));
  assign ConvFiltWidth_else_or_751_cse = (fsm_output[3]) | (fsm_output[5]) | (fsm_output[6]);
  assign ConvFiltWidth_else_mux1h_878_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]),
      (w2_rsci_idat_mxwt[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]),
      (MultLoop_io_read_w4_rsc_cse_sva[8015:8008]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_879_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , ConvFiltWidth_else_or_751_cse , (fsm_output[8])});
  assign mul_197_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_878_nl)) *
      $signed((ConvFiltWidth_else_mux1h_879_nl)));
  assign z_out_605_29_7 = readslicef_30_23_7((mul_197_nl));
  assign ConvFiltWidth_else_or_752_cse = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_880_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (MultLoop_io_read_w4_rsc_cse_sva[2503:2496]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_881_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_198_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_880_nl)) *
      $signed((ConvFiltWidth_else_mux1h_881_nl)));
  assign z_out_606_29_7 = readslicef_30_23_7((mul_198_nl));
  assign ConvFiltWidth_else_mux1h_882_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (w2_rsci_idat_mxwt[367:360]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (MultLoop_io_read_w4_rsc_cse_sva[2055:2048]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_883_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , (fsm_output[8])});
  assign mul_199_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_882_nl)) *
      $signed((ConvFiltWidth_else_mux1h_883_nl)));
  assign z_out_607_29_7 = readslicef_30_23_7((mul_199_nl));
  assign ConvFiltWidth_else_mux1h_884_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (w2_rsci_idat_mxwt[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (MultLoop_io_read_w4_rsc_cse_sva[8023:8016]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_885_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , AccumDotWidth_or_139_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_200_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_884_nl)) *
      $signed((ConvFiltWidth_else_mux1h_885_nl)));
  assign z_out_608_29_7 = readslicef_30_23_7((mul_200_nl));
  assign ConvFiltWidth_else_mux1h_886_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (w2_rsci_idat_mxwt[559:552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (MultLoop_io_read_w4_rsc_cse_sva[2071:2064]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_887_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_201_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_886_nl)) *
      $signed((ConvFiltWidth_else_mux1h_887_nl)));
  assign z_out_609_29_7 = readslicef_30_23_7((mul_201_nl));
  assign ConvFiltWidth_else_mux1h_888_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]),
      (MultLoop_io_read_w4_rsc_cse_sva[5927:5920]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse , (fsm_output[6])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_889_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_87_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_202_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_888_nl)) *
      $signed((ConvFiltWidth_else_mux1h_889_nl)));
  assign z_out_610_29_7 = readslicef_30_23_7((mul_202_nl));
  assign ConvFiltWidth_else_mux1h_890_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]), (w2_rsci_idat_mxwt[359:352]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]),
      (MultLoop_io_read_w4_rsc_cse_sva[5935:5928]), {(fsm_output[2]) , MultLoop_or_22_cse
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_891_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), (input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , MultLoop_or_46_cse
      , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[8])});
  assign mul_203_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_890_nl)) *
      $signed((ConvFiltWidth_else_mux1h_891_nl)));
  assign z_out_611_29_7 = readslicef_30_23_7((mul_203_nl));
  assign ConvFiltWidth_else_mux1h_892_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[543:536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]), (MultLoop_io_read_w4_rsc_cse_sva[5943:5936]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_893_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_751_cse , (fsm_output[8])});
  assign mul_204_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_892_nl)) *
      $signed((ConvFiltWidth_else_mux1h_893_nl)));
  assign z_out_612_29_7 = readslicef_30_23_7((mul_204_nl));
  assign ConvFiltWidth_else_mux1h_894_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[351:344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]), (MultLoop_io_read_w4_rsc_cse_sva[5951:5944]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_895_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_205_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_894_nl)) *
      $signed((ConvFiltWidth_else_mux1h_895_nl)));
  assign z_out_613_29_7 = readslicef_30_23_7((mul_205_nl));
  assign ConvFiltWidth_else_mux1h_896_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]),
      (w2_rsci_idat_mxwt[751:744]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]), (MultLoop_io_read_w4_rsc_cse_sva[5959:5952]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[6]) ,
      (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_897_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , AccumDotWidth_or_157_cse
      , (fsm_output[8])});
  assign mul_206_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_896_nl)) *
      $signed((ConvFiltWidth_else_mux1h_897_nl)));
  assign z_out_614_29_7 = readslicef_30_23_7((mul_206_nl));
  assign ConvFiltWidth_else_mux1h_898_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (w2_rsci_idat_mxwt[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]),
      (MultLoop_io_read_w4_rsc_cse_sva[5903:5896]), {(fsm_output[2]) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_899_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , AccumDotWidth_or_139_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_207_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_898_nl)) *
      $signed((ConvFiltWidth_else_mux1h_899_nl)));
  assign z_out_615_29_7 = readslicef_30_23_7((mul_207_nl));
  assign ConvFiltWidth_else_mux1h_900_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (w2_rsci_idat_mxwt[943:936]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]), (MultLoop_io_read_w4_rsc_cse_sva[2063:2056]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_145_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_901_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_208_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_900_nl)) *
      $signed((ConvFiltWidth_else_mux1h_901_nl)));
  assign z_out_616_29_7 = readslicef_30_23_7((mul_208_nl));
  assign ConvFiltWidth_else_mux1h_902_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]),
      (MultLoop_io_read_w4_rsc_cse_sva[5879:5872]), {(fsm_output[2]) , AccumDotWidth_or_157_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_903_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_209_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_902_nl)) *
      $signed((ConvFiltWidth_else_mux1h_903_nl)));
  assign z_out_617_29_7 = readslicef_30_23_7((mul_209_nl));
  assign ConvFiltWidth_else_mux1h_904_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]),
      (MultLoop_io_read_w4_rsc_cse_sva[5871:5864]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_37_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_210_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_904_nl)) *
      $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_37_nl)));
  assign z_out_618_29_7 = readslicef_30_23_7((mul_210_nl));
  assign ConvFiltWidth_else_mux1h_905_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]),
      (w2_rsci_idat_mxwt[631:624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]),
      (MultLoop_io_read_w4_rsc_cse_sva[5887:5880]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_906_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_29_cse , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_211_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_905_nl)) *
      $signed((ConvFiltWidth_else_mux1h_906_nl)));
  assign z_out_619_29_7 = readslicef_30_23_7((mul_211_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_53_cse = (fsm_output[2])
      | (fsm_output[3]) | (fsm_output[5]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_574_nl = MUX1HOT_v_8_7_2((MultLoop_io_read_w4_rsc_cse_sva[7311:7304]),
      (MultLoop_io_read_w4_rsc_cse_sva[9359:9352]), (w2_rsci_idat_mxwt[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]), (MultLoop_io_read_w4_rsc_cse_sva[143:136]),
      {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_52_nl = (fsm_output[4])
      | (fsm_output[6]) | (fsm_output[8]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_575_nl = MUX1HOT_v_22_3_2(({1'b0
      , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm}),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      {(nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_52_nl) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_53_cse});
  assign mul_212_nl = conv_u2u_30_30($signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_574_nl))
      * $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_575_nl)));
  assign z_out_620_29_7 = readslicef_30_23_7((mul_212_nl));
  assign ConvFiltWidth_else_mux1h_907_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]),
      (MultLoop_io_read_w4_rsc_cse_sva[9863:9856]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_38_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_213_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_907_nl)) *
      $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_38_nl)));
  assign z_out_621_29_7 = readslicef_30_23_7((mul_213_nl));
  assign ConvFiltWidth_else_mux1h_908_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]),
      (MultLoop_io_read_w4_rsc_cse_sva[9823:9816]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_39_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_214_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_908_nl)) *
      $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_39_nl)));
  assign z_out_622_29_7 = readslicef_30_23_7((mul_214_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse = (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_576_nl = MUX1HOT_v_8_8_2((MultLoop_io_read_w4_rsc_cse_sva[8415:8408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]), (w2_rsci_idat_mxwt[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (MultLoop_io_read_w4_rsc_cse_sva[223:216]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_577_nl = MUX1HOT_v_22_4_2(({1'b0
      , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm}),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), (input_1_rsci_idat_mxwt[1055:1034]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_38_cse
      , (fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse});
  assign mul_215_nl = conv_u2u_30_30($signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_576_nl))
      * $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_577_nl)));
  assign z_out_623_29_7 = readslicef_30_23_7((mul_215_nl));
  assign ConvFiltWidth_else_or_787_cse = (fsm_output[7:4]!=4'b0000);
  assign ConvFiltWidth_else_mux1h_909_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]),
      (w2_rsci_idat_mxwt[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (MultLoop_io_read_w4_rsc_cse_sva[9751:9744]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_910_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_787_cse , (fsm_output[8])});
  assign mul_216_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_909_nl)) *
      $signed((ConvFiltWidth_else_mux1h_910_nl)));
  assign z_out_624_29_7 = readslicef_30_23_7((mul_216_nl));
  assign ConvFiltWidth_else_mux1h_911_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]),
      (w2_rsci_idat_mxwt[911:904]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]), (MultLoop_io_read_w4_rsc_cse_sva[9743:9736]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_912_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_787_cse , (fsm_output[8])});
  assign mul_217_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_911_nl)) *
      $signed((ConvFiltWidth_else_mux1h_912_nl)));
  assign z_out_625_29_7 = readslicef_30_23_7((mul_217_nl));
  assign ConvFiltWidth_else_mux1h_913_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]),
      (w2_rsci_idat_mxwt[55:48]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (MultLoop_io_read_w4_rsc_cse_sva[9735:9728]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_914_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[681:660]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_218_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_913_nl)) *
      $signed((ConvFiltWidth_else_mux1h_914_nl)));
  assign z_out_626_29_7 = readslicef_30_23_7((mul_218_nl));
  assign ConvFiltWidth_else_mux1h_915_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]),
      (w2_rsci_idat_mxwt[919:912]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (MultLoop_io_read_w4_rsc_cse_sva[9727:9720]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_916_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse
      , (fsm_output[8])});
  assign mul_219_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_915_nl)) *
      $signed((ConvFiltWidth_else_mux1h_916_nl)));
  assign z_out_627_29_7 = readslicef_30_23_7((mul_219_nl));
  assign ConvFiltWidth_else_mux1h_917_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]),
      (w2_rsci_idat_mxwt[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]), (MultLoop_io_read_w4_rsc_cse_sva[9719:9712]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_918_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse
      , (fsm_output[8])});
  assign mul_220_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_917_nl)) *
      $signed((ConvFiltWidth_else_mux1h_918_nl)));
  assign z_out_628_29_7 = readslicef_30_23_7((mul_220_nl));
  assign ConvFiltWidth_else_mux1h_919_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[247:240]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]),
      (MultLoop_io_read_w4_rsc_cse_sva[9711:9704]), {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_920_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_787_cse , (fsm_output[8])});
  assign mul_221_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_919_nl)) *
      $signed((ConvFiltWidth_else_mux1h_920_nl)));
  assign z_out_629_29_7 = readslicef_30_23_7((mul_221_nl));
  assign ConvFiltWidth_else_mux1h_921_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]),
      (MultLoop_io_read_w4_rsc_cse_sva[6311:6304]), (w2_rsci_idat_mxwt[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (MultLoop_io_read_w4_rsc_cse_sva[167:160]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_922_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm}),
      (input_1_rsci_idat_mxwt[1055:1034]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_53_cse
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse , (fsm_output[1])});
  assign mul_222_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_921_nl)) *
      $signed((ConvFiltWidth_else_mux1h_922_nl)));
  assign z_out_630_29_7 = readslicef_30_23_7((mul_222_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_578_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[7719:7712]),
      (MultLoop_io_read_w4_rsc_cse_sva[3655:3648]), (MultLoop_io_read_w4_rsc_cse_sva[9231:9224]),
      (w4_rsci_idat_mxwt[8167:8160]), (MultLoop_io_read_w4_rsc_cse_sva[9071:9064]),
      (MultLoop_io_read_w4_rsc_cse_sva[6319:6312]), {(fsm_output[5]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_579_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm, nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_mul_223_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_578_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_579_nl));
  assign mul_223_nl = nl_mul_223_nl[28:0];
  assign z_out_631_28_7 = readslicef_29_22_7((mul_223_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_580_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[3039:3032]),
      (MultLoop_io_read_w4_rsc_cse_sva[3615:3608]), (MultLoop_io_read_w4_rsc_cse_sva[4143:4136]),
      (MultLoop_io_read_w4_rsc_cse_sva[8231:8224]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_581_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_5_if_exu_pmx_20_0_lpi_1_dfm, {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_224_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_580_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_581_nl));
  assign mul_224_nl = nl_mul_224_nl[28:0];
  assign z_out_632_28_7 = readslicef_29_22_7((mul_224_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_582_nl = MUX1HOT_v_8_6_2((MultLoop_io_read_w4_rsc_cse_sva[3119:3112]),
      (MultLoop_io_read_w4_rsc_cse_sva[2591:2584]), (w4_rsci_idat_mxwt[967:960]),
      (MultLoop_io_read_w4_rsc_cse_sva[9239:9232]), (MultLoop_io_read_w4_rsc_cse_sva[9079:9072]),
      (MultLoop_io_read_w4_rsc_cse_sva[7743:7736]), {(fsm_output[4]) , (fsm_output[3])
      , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_583_nl = MUX1HOT_v_21_6_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm, nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5])});
  assign nl_mul_225_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_582_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_583_nl));
  assign mul_225_nl = nl_mul_225_nl[28:0];
  assign z_out_633_28_7 = readslicef_29_22_7((mul_225_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_584_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[3023:3016]),
      (MultLoop_io_read_w4_rsc_cse_sva[4295:4288]), (MultLoop_io_read_w4_rsc_cse_sva[3639:3632]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_585_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_226_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_584_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_585_nl));
  assign mul_226_nl = nl_mul_226_nl[28:0];
  assign z_out_634_28_7 = readslicef_29_22_7((mul_226_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_135_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[3663:3656]),
      (w4_rsci_idat_mxwt[975:968]), fsm_output[1]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_136_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[1]);
  assign nl_mul_227_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_135_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_136_nl));
  assign mul_227_nl = nl_mul_227_nl[28:0];
  assign z_out_635_28_7 = readslicef_29_22_7((mul_227_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_586_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1199:1192]),
      (w4_rsci_idat_mxwt[991:984]), (MultLoop_io_read_w4_rsc_cse_sva[4695:4688]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_587_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_228_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_586_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_587_nl));
  assign mul_228_nl = nl_mul_228_nl[28:0];
  assign z_out_636_28_7 = readslicef_29_22_7((mul_228_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_588_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7727:7720]),
      (MultLoop_io_read_w4_rsc_cse_sva[1255:1248]), (w4_rsci_idat_mxwt[1007:1000]),
      (MultLoop_io_read_w4_rsc_cse_sva[4687:4680]), {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_589_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_229_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_588_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_589_nl));
  assign mul_229_nl = nl_mul_229_nl[28:0];
  assign z_out_637_28_7 = readslicef_29_22_7((mul_229_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_590_nl = MUX1HOT_v_8_4_2((w4_rsci_idat_mxwt[8159:8152]),
      (MultLoop_io_read_w4_rsc_cse_sva[4679:4672]), (MultLoop_io_read_w4_rsc_cse_sva[5167:5160]),
      (MultLoop_io_read_w4_rsc_cse_sva[7391:7384]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_591_nl = MUX1HOT_v_21_4_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign nl_mul_230_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_590_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_591_nl));
  assign mul_230_nl = nl_mul_230_nl[28:0];
  assign z_out_638_28_7 = readslicef_29_22_7((mul_230_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_137_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[3031:3024]),
      (MultLoop_io_read_w4_rsc_cse_sva[1607:1600]), fsm_output[3]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_138_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[3]);
  assign nl_mul_231_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_137_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_138_nl));
  assign mul_231_nl = nl_mul_231_nl[28:0];
  assign z_out_639_28_7 = readslicef_29_22_7((mul_231_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_139_nl = MUX_v_8_2_2((w4_rsci_idat_mxwt[3063:3056]),
      (MultLoop_io_read_w4_rsc_cse_sva[1615:1608]), fsm_output[3]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_140_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[3]);
  assign nl_mul_232_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_139_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_140_nl));
  assign mul_232_nl = nl_mul_232_nl[28:0];
  assign z_out_640_28_7 = readslicef_29_22_7((mul_232_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_592_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[1015:1008]),
      (MultLoop_io_read_w4_rsc_cse_sva[1071:1064]), (MultLoop_io_read_w4_rsc_cse_sva[2623:2616]),
      (MultLoop_io_read_w4_rsc_cse_sva[9063:9056]), (MultLoop_io_read_w4_rsc_cse_sva[7415:7408]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_593_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_233_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_592_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_593_nl));
  assign mul_233_nl = nl_mul_233_nl[28:0];
  assign z_out_641_28_7 = readslicef_29_22_7((mul_233_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_594_nl = MUX1HOT_v_8_5_2((w4_rsci_idat_mxwt[7159:7152]),
      (MultLoop_io_read_w4_rsc_cse_sva[6367:6360]), (MultLoop_io_read_w4_rsc_cse_sva[2647:2640]),
      (MultLoop_io_read_w4_rsc_cse_sva[9055:9048]), (MultLoop_io_read_w4_rsc_cse_sva[7407:7400]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_595_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_mul_234_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_594_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_595_nl));
  assign mul_234_nl = nl_mul_234_nl[28:0];
  assign z_out_642_28_7 = readslicef_29_22_7((mul_234_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_596_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[4047:4040]),
      (MultLoop_io_read_w4_rsc_cse_sva[4319:4312]), (MultLoop_io_read_w4_rsc_cse_sva[5663:5656]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_597_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_235_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_596_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_597_nl));
  assign mul_235_nl = nl_mul_235_nl[28:0];
  assign z_out_643_28_7 = readslicef_29_22_7((mul_235_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_598_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[4039:4032]),
      (MultLoop_io_read_w4_rsc_cse_sva[5671:5664]), (MultLoop_io_read_w4_rsc_cse_sva[6191:6184]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_599_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_236_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_598_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_599_nl));
  assign mul_236_nl = nl_mul_236_nl[28:0];
  assign z_out_644_28_7 = readslicef_29_22_7((mul_236_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_600_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[4311:4304]),
      (w4_rsci_idat_mxwt[7111:7104]), (MultLoop_io_read_w4_rsc_cse_sva[5679:5672]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_601_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_237_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_600_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_601_nl));
  assign mul_237_nl = nl_mul_237_nl[28:0];
  assign z_out_645_28_7 = readslicef_29_22_7((mul_237_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_602_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1231:1224]),
      (w4_rsci_idat_mxwt[7119:7112]), (MultLoop_io_read_w4_rsc_cse_sva[5687:5680]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_603_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_238_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_602_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_603_nl));
  assign mul_238_nl = nl_mul_238_nl[28:0];
  assign z_out_646_28_7 = readslicef_29_22_7((mul_238_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_604_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[7127:7120]),
      (MultLoop_io_read_w4_rsc_cse_sva[5335:5328]), (MultLoop_io_read_w4_rsc_cse_sva[5695:5688]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_605_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_239_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_604_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_605_nl));
  assign mul_239_nl = nl_mul_239_nl[28:0];
  assign z_out_647_28_7 = readslicef_29_22_7((mul_239_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_606_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[10095:10088]),
      (w4_rsci_idat_mxwt[8135:8128]), (MultLoop_io_read_w4_rsc_cse_sva[2223:2216]),
      (MultLoop_io_read_w4_rsc_cse_sva[5703:5696]), (MultLoop_io_read_w4_rsc_cse_sva[8239:8232]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_607_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_110_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_22_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_6_if_exu_pmx_20_0_lpi_1_dfm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_240_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_606_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_607_nl));
  assign mul_240_nl = nl_mul_240_nl[28:0];
  assign z_out_648_28_7 = readslicef_29_22_7((mul_240_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_608_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[983:976]),
      (MultLoop_io_read_w4_rsc_cse_sva[5343:5336]), (MultLoop_io_read_w4_rsc_cse_sva[5711:5704]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_609_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_123_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_241_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_608_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_609_nl));
  assign mul_241_nl = nl_mul_241_nl[28:0];
  assign z_out_649_28_7 = readslicef_29_22_7((mul_241_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_610_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[7135:7128]),
      (MultLoop_io_read_w4_rsc_cse_sva[5719:5712]), (MultLoop_io_read_w4_rsc_cse_sva[7215:7208]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_611_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_124_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_mul_242_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_610_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_611_nl));
  assign mul_242_nl = nl_mul_242_nl[28:0];
  assign z_out_650_28_7 = readslicef_29_22_7((mul_242_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_612_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1239:1232]),
      (w4_rsci_idat_mxwt[7143:7136]), (MultLoop_io_read_w4_rsc_cse_sva[4639:4632]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_613_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_243_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_612_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_613_nl));
  assign mul_243_nl = nl_mul_243_nl[28:0];
  assign z_out_651_28_7 = readslicef_29_22_7((mul_243_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_614_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[3055:3048]),
      (MultLoop_io_read_w4_rsc_cse_sva[5327:5320]), (MultLoop_io_read_w4_rsc_cse_sva[4647:4640]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_615_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_244_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_614_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_615_nl));
  assign mul_244_nl = nl_mul_244_nl[28:0];
  assign z_out_652_28_7 = readslicef_29_22_7((mul_244_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_141_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[3671:3664]),
      (w4_rsci_idat_mxwt[3015:3008]), fsm_output[1]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_142_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[1]);
  assign nl_mul_245_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_141_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_142_nl));
  assign mul_245_nl = nl_mul_245_nl[28:0];
  assign z_out_653_28_7 = readslicef_29_22_7((mul_245_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_143_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[2615:2608]),
      (w4_rsci_idat_mxwt[6135:6128]), fsm_output[1]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_144_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      fsm_output[1]);
  assign nl_mul_246_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_143_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_144_nl));
  assign mul_246_nl = nl_mul_246_nl[28:0];
  assign z_out_654_28_7 = readslicef_29_22_7((mul_246_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_616_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[10079:10072]),
      (w4_rsci_idat_mxwt[8143:8136]), (MultLoop_io_read_w4_rsc_cse_sva[6359:6352]),
      (MultLoop_io_read_w4_rsc_cse_sva[2639:2632]), (MultLoop_io_read_w4_rsc_cse_sva[7399:7392]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_617_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_nnet_relu_layer2_t_layer3_t_relu_config3_for_and_107_cse,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_122_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_27_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_29_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_247_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_616_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_617_nl));
  assign mul_247_nl = nl_mul_247_nl[28:0];
  assign z_out_655_28_7 = readslicef_29_22_7((mul_247_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_618_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[10087:10080]),
      (w4_rsci_idat_mxwt[4087:4080]), (MultLoop_io_read_w4_rsc_cse_sva[6351:6344]),
      (MultLoop_io_read_w4_rsc_cse_sva[2631:2624]), (MultLoop_io_read_w4_rsc_cse_sva[8247:8240]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_619_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_109_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_7_if_exu_pmx_20_0_lpi_1_dfm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_248_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_618_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_619_nl));
  assign mul_248_nl = nl_mul_248_nl[28:0];
  assign z_out_656_28_7 = readslicef_29_22_7((mul_248_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_620_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1271:1264]),
      (w4_rsci_idat_mxwt[7151:7144]), (MultLoop_io_read_w4_rsc_cse_sva[1567:1560]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_621_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_31_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_249_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_620_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_621_nl));
  assign mul_249_nl = nl_mul_249_nl[28:0];
  assign z_out_657_28_7 = readslicef_29_22_7((mul_249_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_622_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1263:1256]),
      (w4_rsci_idat_mxwt[4071:4064]), (MultLoop_io_read_w4_rsc_cse_sva[1591:1584]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_623_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_30_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_250_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_622_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_623_nl));
  assign mul_250_nl = nl_mul_250_nl[28:0];
  assign z_out_658_28_7 = readslicef_29_22_7((mul_250_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_624_nl = MUX1HOT_v_8_3_2((w4_rsci_idat_mxwt[999:992]),
      (MultLoop_io_read_w4_rsc_cse_sva[4303:4296]), (MultLoop_io_read_w4_rsc_cse_sva[4655:4648]),
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_625_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_26_if_exu_pmx_20_0_lpi_1_dfm_mx0w2,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_mul_251_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_624_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_625_nl));
  assign mul_251_nl = nl_mul_251_nl[28:0];
  assign z_out_659_28_7 = readslicef_29_22_7((mul_251_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_626_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1223:1216]),
      (w4_rsci_idat_mxwt[3047:3040]), (MultLoop_io_read_w4_rsc_cse_sva[1583:1576]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_627_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_252_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_626_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_627_nl));
  assign mul_252_nl = nl_mul_252_nl[28:0];
  assign z_out_660_28_7 = readslicef_29_22_7((mul_252_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_628_nl = MUX1HOT_v_8_5_2((MultLoop_io_read_w4_rsc_cse_sva[10103:10096]),
      (w4_rsci_idat_mxwt[4079:4072]), (MultLoop_io_read_w4_rsc_cse_sva[6343:6336]),
      (MultLoop_io_read_w4_rsc_cse_sva[1623:1616]), (MultLoop_io_read_w4_rsc_cse_sva[8223:8216]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_629_nl = MUX1HOT_v_21_5_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_111_if_exu_pmx_20_0_lpi_1_dfm_1,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_4_if_exu_pmx_20_0_lpi_1_dfm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_mul_253_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_628_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_629_nl));
  assign mul_253_nl = nl_mul_253_nl[28:0];
  assign z_out_661_28_7 = readslicef_29_22_7((mul_253_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_630_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[1247:1240]),
      (w4_rsci_idat_mxwt[8183:8176]), (MultLoop_io_read_w4_rsc_cse_sva[4663:4656]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_631_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_28_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_127_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_254_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_630_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_631_nl));
  assign mul_254_nl = nl_mul_254_nl[28:0];
  assign z_out_662_28_7 = readslicef_29_22_7((mul_254_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_632_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[5319:5312]),
      (w4_rsci_idat_mxwt[8175:8168]), (MultLoop_io_read_w4_rsc_cse_sva[1575:1568]),
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_633_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_25_if_exu_pmx_20_0_lpi_1_dfm_mx0w3,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_126_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm_mx0w0,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[3])});
  assign nl_mul_255_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_632_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_633_nl));
  assign mul_255_nl = nl_mul_255_nl[28:0];
  assign z_out_663_28_7 = readslicef_29_22_7((mul_255_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse = (fsm_output[2])
      | (fsm_output[8]);
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_634_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7431:7424]),
      (MultLoop_io_read_w4_rsc_cse_sva[9159:9152]), (MultLoop_io_read_w4_rsc_cse_sva[6263:6256]),
      (MultLoop_io_read_w4_rsc_cse_sva[1023:1016]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_635_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_33_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[5]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse
      , (fsm_output[4])});
  assign nl_mul_256_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_634_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_635_nl));
  assign mul_256_nl = nl_mul_256_nl[28:0];
  assign z_out_664_28_7 = readslicef_29_22_7((mul_256_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_636_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7447:7440]),
      (MultLoop_io_read_w4_rsc_cse_sva[9103:9096]), (MultLoop_io_read_w4_rsc_cse_sva[6295:6288]),
      (MultLoop_io_read_w4_rsc_cse_sva[151:144]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_637_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_35_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[5]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse});
  assign nl_mul_257_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_636_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_637_nl));
  assign mul_257_nl = nl_mul_257_nl[28:0];
  assign z_out_665_28_7 = readslicef_29_22_7((mul_257_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_638_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7455:7448]),
      (MultLoop_io_read_w4_rsc_cse_sva[9111:9104]), (MultLoop_io_read_w4_rsc_cse_sva[6303:6296]),
      (MultLoop_io_read_w4_rsc_cse_sva[159:152]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_639_nl = MUX1HOT_v_21_3_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_36_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm,
      {(fsm_output[5]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse});
  assign nl_mul_258_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_638_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_639_nl));
  assign mul_258_nl = nl_mul_258_nl[28:0];
  assign z_out_666_28_7 = readslicef_29_22_7((mul_258_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_640_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7319:7312]),
      (MultLoop_io_read_w4_rsc_cse_sva[9087:9080]), (MultLoop_io_read_w4_rsc_cse_sva[8343:8336]),
      (MultLoop_io_read_w4_rsc_cse_sva[807:800]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_145_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_19_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse);
  assign nl_mul_259_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_640_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_145_nl));
  assign mul_259_nl = nl_mul_259_nl[28:0];
  assign z_out_667_28_7 = readslicef_29_22_7((mul_259_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_641_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7327:7320]),
      (MultLoop_io_read_w4_rsc_cse_sva[9095:9088]), (MultLoop_io_read_w4_rsc_cse_sva[8351:8344]),
      (MultLoop_io_read_w4_rsc_cse_sva[815:808]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_146_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_20_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse);
  assign nl_mul_260_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_641_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_146_nl));
  assign mul_260_nl = nl_mul_260_nl[28:0];
  assign z_out_668_28_7 = readslicef_29_22_7((mul_260_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_642_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[7335:7328]),
      (MultLoop_io_read_w4_rsc_cse_sva[8359:8352]), (MultLoop_io_read_w4_rsc_cse_sva[10111:10104]),
      (MultLoop_io_read_w4_rsc_cse_sva[10023:10016]), {(fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_147_nl = MUX_v_21_2_2(nnet_relu_layer2_t_layer3_t_relu_config3_for_21_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse);
  assign nl_mul_261_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_642_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_147_nl));
  assign mul_261_nl = nl_mul_261_nl[28:0];
  assign z_out_669_28_7 = readslicef_29_22_7((mul_261_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_643_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9391:9384]),
      (MultLoop_io_read_w4_rsc_cse_sva[9119:9112]), (MultLoop_io_read_w4_rsc_cse_sva[8367:8360]),
      (MultLoop_io_read_w4_rsc_cse_sva[175:168]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_8_nl
      = MUX_v_21_2_2(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[2]);
  assign nl_mul_262_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_643_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_8_nl));
  assign mul_262_nl = nl_mul_262_nl[28:0];
  assign z_out_670_28_7 = readslicef_29_22_7((mul_262_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_644_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9399:9392]),
      (MultLoop_io_read_w4_rsc_cse_sva[9127:9120]), (MultLoop_io_read_w4_rsc_cse_sva[8375:8368]),
      (MultLoop_io_read_w4_rsc_cse_sva[183:176]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_9_nl
      = MUX_v_21_2_2(ConvOutHeight_1_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[2]);
  assign nl_mul_263_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_644_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_9_nl));
  assign mul_263_nl = nl_mul_263_nl[28:0];
  assign z_out_671_28_7 = readslicef_29_22_7((mul_263_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_645_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9407:9400]),
      (MultLoop_io_read_w4_rsc_cse_sva[8383:8376]), (MultLoop_io_read_w4_rsc_cse_sva[191:184]),
      {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_264_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_645_nl))
      * $signed(conv_u2s_21_22(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_1_ConvFiltHeight_2_ConvFiltWidth_1_else_slc_29_9_itm));
  assign mul_264_nl = nl_mul_264_nl[28:0];
  assign z_out_672_28_7 = readslicef_29_22_7((mul_264_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_646_nl = MUX1HOT_v_8_3_2((MultLoop_io_read_w4_rsc_cse_sva[9415:9408]),
      (MultLoop_io_read_w4_rsc_cse_sva[8391:8384]), (MultLoop_io_read_w4_rsc_cse_sva[199:192]),
      {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[8])});
  assign nl_mul_265_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_646_nl))
      * $signed(conv_u2s_21_22(ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm));
  assign mul_265_nl = nl_mul_265_nl[28:0];
  assign z_out_673_28_7 = readslicef_29_22_7((mul_265_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_647_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9423:9416]),
      (MultLoop_io_read_w4_rsc_cse_sva[9135:9128]), (MultLoop_io_read_w4_rsc_cse_sva[8399:8392]),
      (MultLoop_io_read_w4_rsc_cse_sva[207:200]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[5]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_10_nl
      = MUX_v_21_2_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[2]);
  assign nl_mul_266_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_647_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_10_nl));
  assign mul_266_nl = nl_mul_266_nl[28:0];
  assign z_out_674_28_7 = readslicef_29_22_7((mul_266_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_648_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[9431:9424]),
      (MultLoop_io_read_w4_rsc_cse_sva[8407:8400]), (MultLoop_io_read_w4_rsc_cse_sva[10183:10176]),
      (MultLoop_io_read_w4_rsc_cse_sva[215:208]), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_11_nl
      = MUX_v_21_2_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm,
      fsm_output[2]);
  assign nl_mul_267_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_648_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_11_nl));
  assign mul_267_nl = nl_mul_267_nl[28:0];
  assign z_out_675_28_7 = readslicef_29_22_7((mul_267_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_649_nl = MUX1HOT_v_8_4_2((MultLoop_io_read_w4_rsc_cse_sva[8335:8328]),
      (MultLoop_io_read_w4_rsc_cse_sva[10119:10112]), (MultLoop_io_read_w4_rsc_cse_sva[6287:6280]),
      (MultLoop_io_read_w4_rsc_cse_sva[10031:10024]), {(fsm_output[5]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[8])});
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_12_nl
      = MUX_v_21_2_2(ConvOutHeight_3_ConvOutWidth_1_ConvFilt_7_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm,
      nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm,
      nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse);
  assign nl_mul_268_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux1h_649_nl))
      * $signed(conv_u2s_21_22(nnet_product_layer3_t_config4_weight_t_config4_accum_t_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_12_nl));
  assign mul_268_nl = nl_mul_268_nl[28:0];
  assign z_out_676_28_7 = readslicef_29_22_7((mul_268_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_148_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7231:7224]),
      (MultLoop_io_read_w4_rsc_cse_sva[63:56]), fsm_output[8]);
  assign nl_mul_269_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_148_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_8_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_269_nl = nl_mul_269_nl[28:0];
  assign z_out_677_28_7 = readslicef_29_22_7((mul_269_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_149_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7239:7232]),
      (MultLoop_io_read_w4_rsc_cse_sva[71:64]), fsm_output[8]);
  assign nl_mul_270_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_149_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_9_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_270_nl = nl_mul_270_nl[28:0];
  assign z_out_678_28_7 = readslicef_29_22_7((mul_270_nl));
  assign nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_150_nl = MUX_v_8_2_2((MultLoop_io_read_w4_rsc_cse_sva[7287:7280]),
      (MultLoop_io_read_w4_rsc_cse_sva[119:112]), fsm_output[8]);
  assign nl_mul_271_nl = $signed((nnet_product_layer3_t_config4_weight_t_config4_accum_t_mux_150_nl))
      * $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_125_if_exu_pmx_20_0_lpi_1_dfm));
  assign mul_271_nl = nl_mul_271_nl[28:0];
  assign z_out_679_28_7 = readslicef_29_22_7((mul_271_nl));
  assign nl_AccumDotWidth_acc_2678_nl = (z_out_623_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2678_nl = nl_AccumDotWidth_acc_2678_nl[9:0];
  assign AccumDotWidth_mux1h_1234_nl = MUX1HOT_v_21_7_2((z_out_1037_29_7[22:2]),
      (z_out_924_29_7[22:2]), z_out_989_29_9, ({(AccumDotWidth_acc_2678_nl) , (z_out_623_29_7[12:2])}),
      (z_out_1050_29_7[22:2]), (z_out_1053_29_7[22:2]), (z_out_1096_29_7[22:2]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1235_nl = MUX1HOT_v_21_7_2((z_out_1038_29_7[22:2]),
      (z_out_938_29_7[22:2]), (z_out_919_29_7[22:2]), (z_out_985_29_7[22:2]), (z_out_1145_29_7[22:2]),
      (z_out_945_29_7[22:2]), (z_out_1146_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_680 = conv_s2u_21_22(AccumDotWidth_mux1h_1234_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1235_nl);
  assign z_out_680 = nl_z_out_680[21:0];
  assign nl_AccumDotWidth_acc_2679_nl = (z_out_627_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]);
  assign AccumDotWidth_acc_2679_nl = nl_AccumDotWidth_acc_2679_nl[9:0];
  assign nl_AccumDotWidth_acc_2680_nl = (z_out_623_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[23:16]);
  assign AccumDotWidth_acc_2680_nl = nl_AccumDotWidth_acc_2680_nl[9:0];
  assign AccumDotWidth_mux1h_1236_nl = MUX1HOT_v_21_7_2((z_out_572_29_7[22:2]), (z_out_947_29_7[22:2]),
      ({(AccumDotWidth_acc_2679_nl) , (z_out_627_29_7[12:2])}), ({(AccumDotWidth_acc_2680_nl)
      , (z_out_623_29_7[12:2])}), (z_out_955_29_7[22:2]), (z_out_936_29_7[22:2]),
      (z_out_570_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1237_nl = MUX1HOT_v_21_6_2((z_out_875_29_7[22:2]), (z_out_941_29_7[22:2]),
      z_out_993_29_9, (z_out_602_29_7[22:2]), (z_out_596_29_7[22:2]), (z_out_938_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6])});
  assign nl_z_out_681 = conv_s2u_21_22(AccumDotWidth_mux1h_1236_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1237_nl);
  assign z_out_681 = nl_z_out_681[21:0];
  assign AccumDotWidth_mux1h_1238_nl = MUX1HOT_v_21_6_2((z_out_999_29_7[22:2]), (z_out_943_29_7[22:2]),
      (z_out_1157_29_7[22:2]), (z_out_1160_29_7[22:2]), (z_out_1169_29_7[22:2]),
      (z_out_1162_29_7[22:2]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1239_nl = MUX1HOT_v_21_7_2((z_out_1009_29_7[22:2]),
      (z_out_940_29_7[22:2]), (z_out_949_29_7[22:2]), (z_out_995_29_7[22:2]), (z_out_926_29_7[22:2]),
      (z_out_1084_29_7[22:2]), (z_out_857_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_682 = conv_s2u_21_22(AccumDotWidth_mux1h_1238_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1239_nl);
  assign z_out_682 = nl_z_out_682[21:0];
  assign nl_AccumDotWidth_acc_2681_nl = (z_out_1027_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2681_nl = nl_AccumDotWidth_acc_2681_nl[9:0];
  assign nl_AccumDotWidth_acc_2682_nl = (z_out_896_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[7:0]);
  assign AccumDotWidth_acc_2682_nl = nl_AccumDotWidth_acc_2682_nl[9:0];
  assign AccumDotWidth_mux1h_1240_nl = MUX1HOT_v_10_6_2((z_out_1106_29_7[22:13]),
      z_out_25, (AccumDotWidth_acc_2681_nl), (z_out_958_29_7[22:13]), (z_out_1153_29_7[22:13]),
      (AccumDotWidth_acc_2682_nl), {(fsm_output[2]) , AccumDotWidth_or_132_cse_1
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1241_nl = MUX1HOT_v_11_7_2((z_out_1106_29_7[12:2]),
      (z_out_628_29_7[12:2]), (z_out_1027_29_7[12:2]), (z_out_627_29_7[12:2]), (z_out_958_29_7[12:2]),
      (z_out_1153_29_7[12:2]), (z_out_896_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1242_nl = MUX1HOT_v_21_7_2((z_out_976_29_7[22:2]), (z_out_626_29_7[22:2]),
      (z_out_576_29_7[22:2]), (z_out_897_29_7[22:2]), (z_out_599_29_7[22:2]), (z_out_947_29_7[22:2]),
      (z_out_1108_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_683 = conv_s2u_21_22({(AccumDotWidth_mux1h_1240_nl) , (AccumDotWidth_mux1h_1241_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_1242_nl);
  assign z_out_683 = nl_z_out_683[21:0];
  assign nl_AccumDotWidth_acc_2683_nl = (z_out_1032_29_9[20:11]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2683_nl = nl_AccumDotWidth_acc_2683_nl[9:0];
  assign nl_AccumDotWidth_acc_2684_nl = (z_out_622_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[15:8]);
  assign AccumDotWidth_acc_2684_nl = nl_AccumDotWidth_acc_2684_nl[9:0];
  assign AccumDotWidth_mux1h_1243_nl = MUX1HOT_v_21_7_2((z_out_944_29_7[22:2]), (z_out_1035_29_7[22:2]),
      ({(AccumDotWidth_acc_2683_nl) , (z_out_1032_29_9[10:0])}), ({(AccumDotWidth_acc_2684_nl)
      , (z_out_622_29_7[12:2])}), z_out_1134_29_9, (z_out_1110_29_7[22:2]), (z_out_1097_29_7[22:2]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1244_nl = MUX1HOT_v_21_7_2((z_out_953_29_7[22:2]), (z_out_1055_29_7[22:2]),
      (z_out_577_29_7[22:2]), (z_out_600_29_7[22:2]), (z_out_1016_29_7[22:2]), (z_out_1147_29_7[22:2]),
      z_out_904_29_9, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_684 = conv_s2u_21_22(AccumDotWidth_mux1h_1243_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1244_nl);
  assign z_out_684 = nl_z_out_684[21:0];
  assign AccumDotWidth_mux1h_754_nl = MUX1HOT_v_10_3_2((z_out_620_29_7[22:13]), (z_out_628_29_7[22:13]),
      (z_out_625_29_7[22:13]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])});
  assign AccumDotWidth_AccumDotWidth_mux_17_nl = MUX_v_8_2_2((b2_rsci_idat_mxwt[47:40]),
      (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[39:32]),
      MultLoop_or_46_cse);
  assign nl_AccumDotWidth_acc_2730_nl = (AccumDotWidth_mux1h_754_nl) + conv_s2u_8_10(AccumDotWidth_AccumDotWidth_mux_17_nl);
  assign AccumDotWidth_acc_2730_nl = nl_AccumDotWidth_acc_2730_nl[9:0];
  assign nl_AccumDotWidth_acc_2685_nl = (z_out_933_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[55:48]);
  assign AccumDotWidth_acc_2685_nl = nl_AccumDotWidth_acc_2685_nl[9:0];
  assign AccumDotWidth_or_209_nl = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]);
  assign AccumDotWidth_mux1h_1245_nl = MUX1HOT_v_10_5_2((z_out_954_29_7[22:13]),
      (AccumDotWidth_acc_2730_nl), (z_out_956_29_7[22:13]), (z_out_855_29_7[22:13]),
      (AccumDotWidth_acc_2685_nl), {(fsm_output[2]) , (AccumDotWidth_or_209_nl) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1246_nl = MUX1HOT_v_11_7_2((z_out_954_29_7[12:2]), (z_out_620_29_7[12:2]),
      (z_out_628_29_7[12:2]), (z_out_625_29_7[12:2]), (z_out_956_29_7[12:2]), (z_out_855_29_7[12:2]),
      (z_out_933_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1247_nl = MUX1HOT_v_21_6_2(z_out_1142_29_9, (z_out_1167_29_7[22:2]),
      (z_out_980_29_7[22:2]), (z_out_601_29_7[22:2]), (z_out_877_29_7[22:2]), (z_out_1128_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_685 = conv_s2u_21_22({(AccumDotWidth_mux1h_1245_nl) , (AccumDotWidth_mux1h_1246_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_1247_nl);
  assign z_out_685 = nl_z_out_685[21:0];
  assign nl_AccumDotWidth_acc_2686_nl = (z_out_890_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2686_nl = nl_AccumDotWidth_acc_2686_nl[9:0];
  assign nl_AccumDotWidth_acc_2687_nl = (z_out_936_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[63:56]);
  assign AccumDotWidth_acc_2687_nl = nl_AccumDotWidth_acc_2687_nl[9:0];
  assign AccumDotWidth_mux1h_1248_nl = MUX1HOT_v_10_6_2((z_out_1024_29_7[22:13]),
      z_out_28, (AccumDotWidth_acc_2686_nl), (z_out_957_29_7[22:13]), (z_out_1155_29_7[22:13]),
      (AccumDotWidth_acc_2687_nl), {(fsm_output[2]) , AccumDotWidth_or_132_cse_1
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1249_nl = MUX1HOT_v_11_7_2((z_out_1024_29_7[12:2]),
      (z_out_630_29_7[12:2]), (z_out_890_29_7[12:2]), (z_out_629_29_7[12:2]), (z_out_957_29_7[12:2]),
      (z_out_1155_29_7[12:2]), (z_out_936_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1250_nl = MUX1HOT_v_21_6_2((z_out_1000_29_7[22:2]),
      (z_out_1160_29_7[22:2]), (z_out_575_29_7[22:2]), (z_out_604_29_7[22:2]), (z_out_943_29_7[22:2]),
      (z_out_1124_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , AccumDotWidth_or_38_cse , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_686 = conv_s2u_21_22({(AccumDotWidth_mux1h_1248_nl) , (AccumDotWidth_mux1h_1249_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_1250_nl);
  assign z_out_686 = nl_z_out_686[21:0];
  assign AccumDotWidth_mux_79_nl = MUX_v_10_2_2((z_out_627_29_7[22:13]), (z_out_624_29_7[22:13]),
      fsm_output[4]);
  assign AccumDotWidth_mux_80_nl = MUX_v_8_2_2((b2_rsci_idat_mxwt[23:16]), (nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[31:24]),
      fsm_output[4]);
  assign nl_AccumDotWidth_acc_2728_nl = (AccumDotWidth_mux_79_nl) + conv_s2u_8_10(AccumDotWidth_mux_80_nl);
  assign AccumDotWidth_acc_2728_nl = nl_AccumDotWidth_acc_2728_nl[9:0];
  assign nl_AccumDotWidth_acc_2688_nl = (z_out_931_29_7[22:13]) + conv_s2s_8_10(nnet_conv_2d_input_t_layer2_t_config2_for_for_for_io_read_b2_rsc_cse_sva[47:40]);
  assign AccumDotWidth_acc_2688_nl = nl_AccumDotWidth_acc_2688_nl[9:0];
  assign AccumDotWidth_mux1h_1251_nl = MUX1HOT_v_10_6_2((z_out_991_29_7[22:13]),
      (AccumDotWidth_acc_2728_nl), z_out_28, (z_out_1056_29_7[22:13]), (z_out_1170_29_7[22:13]),
      (AccumDotWidth_acc_2688_nl), {(fsm_output[2]) , AccumDotWidth_or_132_cse_1
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1252_nl = MUX1HOT_v_11_7_2((z_out_991_29_7[12:2]), (z_out_627_29_7[12:2]),
      (z_out_622_29_7[12:2]), (z_out_624_29_7[12:2]), (z_out_1056_29_7[12:2]), (z_out_1170_29_7[12:2]),
      (z_out_931_29_7[12:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1253_nl = MUX1HOT_v_21_7_2((z_out_574_29_7[22:2]), (z_out_1173_29_7[22:2]),
      (z_out_982_29_7[22:2]), (z_out_596_29_7[22:2]), (z_out_1148_29_7[22:2]), (z_out_913_29_7[22:2]),
      (z_out_1127_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_687 = conv_s2u_21_22({(AccumDotWidth_mux1h_1251_nl) , (AccumDotWidth_mux1h_1252_nl)})
      + conv_s2u_21_22(AccumDotWidth_mux1h_1253_nl);
  assign z_out_687 = nl_z_out_687[21:0];
  assign AccumDotWidth_mux1h_1254_nl = MUX1HOT_v_21_7_2((z_out_596_29_7[22:2]), ({z_out_27
      , (z_out_623_29_7[12:2])}), ({z_out_32 , (z_out_621_29_7[12:2])}), ({z_out_33
      , (z_out_628_29_7[12:2])}), (z_out_1057_29_7[22:2]), (z_out_1173_29_7[22:2]),
      ({z_out_30 , (z_out_929_29_7[12:2])}), {(fsm_output[2]) , (fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1255_nl = MUX1HOT_v_21_7_2((z_out_1156_29_7[22:2]),
      (z_out_1172_29_7[22:2]), (z_out_981_29_7[22:2]), (z_out_603_29_7[22:2]), (z_out_1152_29_7[22:2]),
      (z_out_914_29_7[22:2]), (z_out_1109_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_688 = conv_s2u_21_22(AccumDotWidth_mux1h_1254_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1255_nl);
  assign z_out_688 = nl_z_out_688[21:0];
  assign AccumDotWidth_mux1h_1256_nl = MUX1HOT_v_21_7_2((z_out_1084_29_7[22:2]),
      (z_out_954_29_7[22:2]), (z_out_1147_29_7[22:2]), (z_out_1076_29_7[22:2]), (z_out_572_29_7[22:2]),
      (z_out_944_29_7[22:2]), (z_out_1095_29_7[22:2]), {(fsm_output[4]) , (fsm_output[3])
      , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1257_nl = MUX1HOT_v_21_7_2((z_out_854_29_7[22:2]), z_out_904_29_9,
      (z_out_1130_29_7[22:2]), (z_out_1079_29_7[22:2]), (z_out_994_29_7[22:2]), (z_out_1124_29_7[22:2]),
      (z_out_1147_29_7[22:2]), {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_689 = conv_s2u_21_22(AccumDotWidth_mux1h_1256_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1257_nl);
  assign z_out_689 = nl_z_out_689[21:0];
  assign AccumDotWidth_mux1h_1258_nl = MUX1HOT_v_21_7_2((z_out_1115_29_7[22:2]),
      (z_out_1074_29_7[22:2]), (z_out_1118_29_7[22:2]), (z_out_1163_29_7[22:2]),
      (z_out_1077_29_7[22:2]), (z_out_623_29_7[22:2]), (z_out_926_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1259_nl = MUX1HOT_v_21_7_2((z_out_1154_29_7[22:2]),
      (z_out_1073_29_7[22:2]), (z_out_1157_29_7[22:2]), (z_out_1174_29_7[22:2]),
      (z_out_1007_29_7[22:2]), (z_out_899_29_7[22:2]), (z_out_605_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_690 = conv_s2u_21_22(AccumDotWidth_mux1h_1258_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1259_nl);
  assign z_out_690 = nl_z_out_690[21:0];
  assign AccumDotWidth_mux1h_1260_nl = MUX1HOT_v_21_7_2((z_out_1173_29_7[22:2]),
      (z_out_1075_29_7[22:2]), (z_out_1117_29_7[22:2]), (z_out_975_29_7[22:2]), (z_out_1094_29_7[22:2]),
      (z_out_871_29_7[22:2]), (z_out_569_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1261_nl = MUX1HOT_v_21_7_2((z_out_854_29_7[22:2]), z_out_1063_29_9,
      (z_out_912_29_7[22:2]), (z_out_1180_29_7[22:2]), (z_out_950_29_7[22:2]), (z_out_1097_29_7[22:2]),
      (z_out_986_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_691 = conv_s2u_21_22(AccumDotWidth_mux1h_1260_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1261_nl);
  assign z_out_691 = nl_z_out_691[21:0];
  assign AccumDotWidth_mux1h_1262_nl = MUX1HOT_v_21_7_2((z_out_945_29_7[22:2]), (z_out_1069_29_7[22:2]),
      (z_out_944_29_7[22:2]), (z_out_1158_29_7[22:2]), (z_out_868_29_7[22:2]), (z_out_621_29_7[22:2]),
      (z_out_1173_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1263_nl = MUX1HOT_v_21_7_2((z_out_1108_29_7[22:2]),
      (z_out_1068_29_7[22:2]), (z_out_854_29_7[22:2]), (z_out_1125_29_7[22:2]), (z_out_886_29_7[22:2]),
      (z_out_895_29_7[22:2]), (z_out_915_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_692 = conv_s2u_21_22(AccumDotWidth_mux1h_1262_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1263_nl);
  assign z_out_692 = nl_z_out_692[21:0];
  assign AccumDotWidth_mux1h_1264_nl = MUX1HOT_v_21_7_2(z_out_904_29_9, (z_out_1071_29_7[22:2]),
      (z_out_1186_29_7[22:2]), (z_out_998_29_7[22:2]), (z_out_1112_29_7[22:2]), (z_out_1096_29_7[22:2]),
      (z_out_927_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1265_nl = MUX1HOT_v_21_7_2((z_out_1152_29_7[22:2]),
      (z_out_1070_29_7[22:2]), (z_out_891_29_7[22:2]), (z_out_896_29_7[22:2]), (z_out_931_29_7[22:2]),
      (z_out_1160_29_7[22:2]), (z_out_611_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_693 = conv_s2u_21_22(AccumDotWidth_mux1h_1264_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1265_nl);
  assign z_out_693 = nl_z_out_693[21:0];
  assign AccumDotWidth_mux1h_1266_nl = MUX1HOT_v_21_7_2((z_out_1028_29_7[22:2]),
      z_out_1062_29_9, (z_out_956_29_7[22:2]), (z_out_1092_29_7[22:2]), (z_out_1044_29_7[22:2]),
      (z_out_628_29_7[22:2]), (z_out_923_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1267_nl = MUX1HOT_v_21_7_2((z_out_1013_29_7[22:2]),
      (z_out_896_29_7[22:2]), (z_out_599_29_7[22:2]), z_out_1136_29_9, (z_out_859_29_7[22:2]),
      (z_out_898_29_7[22:2]), (z_out_607_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_694 = conv_s2u_21_22(AccumDotWidth_mux1h_1266_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1267_nl);
  assign z_out_694 = nl_z_out_694[21:0];
  assign AccumDotWidth_mux1h_1268_nl = MUX1HOT_v_21_7_2((z_out_1160_29_7[22:2]),
      (z_out_861_29_7[22:2]), (z_out_943_29_7[22:2]), (z_out_1035_29_7[22:2]), (z_out_944_29_7[22:2]),
      (z_out_867_29_7[22:2]), (z_out_1170_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1269_nl = MUX1HOT_v_21_7_2((z_out_855_29_7[22:2]), (z_out_858_29_7[22:2]),
      (z_out_860_29_7[22:2]), (z_out_1076_29_7[22:2]), (z_out_1162_29_7[22:2]), (z_out_1092_29_7[22:2]),
      (z_out_1080_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_695 = conv_s2u_21_22(AccumDotWidth_mux1h_1268_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1269_nl);
  assign z_out_695 = nl_z_out_695[21:0];
  assign AccumDotWidth_mux1h_1270_nl = MUX1HOT_v_21_7_2((z_out_1151_29_7[22:2]),
      (z_out_853_29_7[22:2]), (z_out_1000_29_7[22:2]), (z_out_991_29_7[22:2]), (z_out_922_29_7[22:2]),
      z_out_1004_29_9, (z_out_865_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1271_nl = MUX1HOT_v_21_7_2((z_out_1125_29_7[22:2]),
      (z_out_854_29_7[22:2]), (z_out_1169_29_7[22:2]), (z_out_1072_29_7[22:2]), (z_out_1087_29_7[22:2]),
      (z_out_1100_29_7[22:2]), (z_out_967_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_696 = conv_s2u_21_22(AccumDotWidth_mux1h_1270_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1271_nl);
  assign z_out_696 = nl_z_out_696[21:0];
  assign AccumDotWidth_mux1h_1272_nl = MUX1HOT_v_21_7_2(z_out_1047_29_9, (z_out_857_29_7[22:2]),
      (z_out_619_29_7[22:2]), (z_out_909_29_7[22:2]), (z_out_1027_29_7[22:2]), (z_out_629_29_7[22:2]),
      (z_out_1145_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1273_nl = MUX1HOT_v_21_7_2((z_out_907_29_7[22:2]), (z_out_859_29_7[22:2]),
      (z_out_1043_29_7[22:2]), (z_out_1075_29_7[22:2]), (z_out_621_29_7[22:2]), (z_out_905_29_7[22:2]),
      (z_out_941_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_697 = conv_s2u_21_22(AccumDotWidth_mux1h_1272_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1273_nl);
  assign z_out_697 = nl_z_out_697[21:0];
  assign AccumDotWidth_mux1h_1274_nl = MUX1HOT_v_21_7_2((z_out_1116_29_7[22:2]),
      (z_out_1078_29_7[22:2]), (z_out_951_29_7[22:2]), (z_out_997_29_7[22:2]), (z_out_1174_29_7[22:2]),
      (z_out_619_29_7[22:2]), (z_out_998_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1275_nl = MUX1HOT_v_21_7_2((z_out_1149_29_7[22:2]),
      (z_out_1072_29_7[22:2]), (z_out_1074_29_7[22:2]), (z_out_905_29_7[22:2]), (z_out_930_29_7[22:2]),
      (z_out_900_29_7[22:2]), (z_out_1069_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_698 = conv_s2u_21_22(AccumDotWidth_mux1h_1274_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1275_nl);
  assign z_out_698 = nl_z_out_698[21:0];
  assign AccumDotWidth_mux1h_1276_nl = MUX1HOT_v_21_6_2((z_out_947_29_7[22:2]), (z_out_865_29_7[22:2]),
      (z_out_966_29_7[22:2]), (z_out_955_29_7[22:2]), (z_out_914_29_7[22:2]), (z_out_870_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , AccumDotWidth_or_140_cse});
  assign AccumDotWidth_mux1h_1277_nl = MUX1HOT_v_21_6_2((z_out_1128_29_7[22:2]),
      (z_out_860_29_7[22:2]), (z_out_1078_29_7[22:2]), (z_out_1110_29_7[22:2]), (z_out_1081_29_7[22:2]),
      (z_out_1028_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , AccumDotWidth_or_140_cse});
  assign nl_z_out_699 = conv_s2u_21_22(AccumDotWidth_mux1h_1276_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1277_nl);
  assign z_out_699 = nl_z_out_699[21:0];
  assign AccumDotWidth_mux1h_1278_nl = MUX1HOT_v_21_7_2((z_out_1035_29_7[22:2]),
      (z_out_1185_29_7[22:2]), (z_out_626_29_7[22:2]), (z_out_911_29_7[22:2]), (z_out_946_29_7[22:2]),
      (z_out_872_29_7[22:2]), z_out_1047_29_9, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1279_nl = MUX1HOT_v_21_7_2((z_out_952_29_7[22:2]), (z_out_1019_29_7[22:2]),
      (z_out_914_29_7[22:2]), (z_out_859_29_7[22:2]), (z_out_1171_29_7[22:2]), (z_out_1022_29_7[22:2]),
      (z_out_872_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_700 = conv_s2u_21_22(AccumDotWidth_mux1h_1278_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1279_nl);
  assign z_out_700 = nl_z_out_700[21:0];
  assign AccumDotWidth_mux1h_1280_nl = MUX1HOT_v_21_7_2((z_out_1103_29_7[22:2]),
      (z_out_929_29_7[22:2]), z_out_1142_29_9, (z_out_1152_29_7[22:2]), z_out_1020_29_9,
      (z_out_934_29_7[22:2]), (z_out_597_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1281_nl = MUX1HOT_v_21_7_2((z_out_967_29_7[22:2]), (z_out_580_29_7[22:2]),
      (z_out_583_29_7[22:2]), z_out_1137_29_9, (z_out_612_29_7[22:2]), (z_out_966_29_7[22:2]),
      z_out_1017_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_701 = conv_s2u_21_22(AccumDotWidth_mux1h_1280_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1281_nl);
  assign z_out_701 = nl_z_out_701[21:0];
  assign AccumDotWidth_mux1h_1282_nl = MUX1HOT_v_21_7_2((z_out_1114_29_7[22:2]),
      (z_out_915_29_7[22:2]), (z_out_592_29_7[22:2]), (z_out_961_29_7[22:2]), (z_out_975_29_7[22:2]),
      (z_out_974_29_7[22:2]), (z_out_571_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1283_nl = MUX1HOT_v_21_7_2((z_out_1145_29_7[22:2]),
      (z_out_913_29_7[22:2]), (z_out_607_29_7[22:2]), (z_out_1120_29_7[22:2]), (z_out_966_29_7[22:2]),
      (z_out_937_29_7[22:2]), (z_out_982_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_702 = conv_s2u_21_22(AccumDotWidth_mux1h_1282_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1283_nl);
  assign z_out_702 = nl_z_out_702[21:0];
  assign AccumDotWidth_mux1h_1284_nl = MUX1HOT_v_21_7_2((z_out_990_29_7[22:2]), (z_out_857_29_7[22:2]),
      (z_out_1155_29_7[22:2]), z_out_1003_29_9, (z_out_1023_29_7[22:2]), (z_out_574_29_7[22:2]),
      (z_out_1167_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1285_nl = MUX1HOT_v_21_7_2((z_out_1019_29_7[22:2]),
      (z_out_591_29_7[22:2]), (z_out_935_29_7[22:2]), (z_out_908_29_7[22:2]), (z_out_619_29_7[22:2]),
      (z_out_1159_29_7[22:2]), (z_out_1091_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_703 = conv_s2u_21_22(AccumDotWidth_mux1h_1284_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1285_nl);
  assign z_out_703 = nl_z_out_703[21:0];
  assign AccumDotWidth_mux1h_1286_nl = MUX1HOT_v_21_7_2(z_out_993_29_9, (z_out_577_29_7[22:2]),
      z_out_962_29_9, (z_out_1104_29_7[22:2]), (z_out_610_29_7[22:2]), (z_out_1105_29_7[22:2]),
      (z_out_1019_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1287_nl = MUX1HOT_v_21_7_2((z_out_630_29_7[22:2]), (z_out_578_29_7[22:2]),
      (z_out_897_29_7[22:2]), (z_out_1181_29_7[22:2]), (z_out_1041_29_7[22:2]), (z_out_1152_29_7[22:2]),
      (z_out_1050_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_704 = conv_s2u_21_22(AccumDotWidth_mux1h_1286_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1287_nl);
  assign z_out_704 = nl_z_out_704[21:0];
  assign AccumDotWidth_mux1h_1288_nl = MUX1HOT_v_21_7_2((z_out_1005_29_7[22:2]),
      z_out_1144_29_9, (z_out_589_29_7[22:2]), (z_out_964_29_7[22:2]), (z_out_921_29_7[22:2]),
      (z_out_1164_29_7[22:2]), (z_out_1052_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1289_nl = MUX1HOT_v_21_7_2((z_out_1021_29_7[22:2]),
      (z_out_1088_29_7[22:2]), (z_out_605_29_7[22:2]), (z_out_1071_29_7[22:2]), (z_out_1084_29_7[22:2]),
      (z_out_1081_29_7[22:2]), (z_out_596_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_705 = conv_s2u_21_22(AccumDotWidth_mux1h_1288_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1289_nl);
  assign z_out_705 = nl_z_out_705[21:0];
  assign AccumDotWidth_mux1h_1290_nl = MUX1HOT_v_21_7_2((z_out_1167_29_7[22:2]),
      (z_out_579_29_7[22:2]), (z_out_888_29_7[22:2]), (z_out_960_29_7[22:2]), (z_out_889_29_7[22:2]),
      z_out_1188_29_9, (z_out_574_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1291_nl = MUX1HOT_v_21_7_2((z_out_1090_29_7[22:2]),
      (z_out_575_29_7[22:2]), (z_out_927_29_7[22:2]), (z_out_1117_29_7[22:2]), z_out_1032_29_9,
      (z_out_1013_29_7[22:2]), z_out_992_29_9, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_706 = conv_s2u_21_22(AccumDotWidth_mux1h_1290_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1291_nl);
  assign z_out_706 = nl_z_out_706[21:0];
  assign AccumDotWidth_mux1h_1292_nl = MUX1HOT_v_21_7_2((z_out_920_29_7[22:2]), (z_out_581_29_7[22:2]),
      (z_out_1001_29_7[22:2]), (z_out_1148_29_7[22:2]), (z_out_580_29_7[22:2]), (z_out_929_29_7[22:2]),
      (z_out_855_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1293_nl = MUX1HOT_v_21_7_2((z_out_577_29_7[22:2]), (z_out_576_29_7[22:2]),
      (z_out_964_29_7[22:2]), (z_out_1109_29_7[22:2]), (z_out_996_29_7[22:2]), (z_out_903_29_7[22:2]),
      (z_out_893_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_707 = conv_s2u_21_22(AccumDotWidth_mux1h_1292_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1293_nl);
  assign z_out_707 = nl_z_out_707[21:0];
  assign AccumDotWidth_mux1h_1294_nl = MUX1HOT_v_21_6_2((z_out_1045_29_7[22:2]),
      (z_out_597_29_7[22:2]), (z_out_972_29_7[22:2]), (z_out_910_29_7[22:2]), (z_out_872_29_7[22:2]),
      z_out_1136_29_9, {AccumDotWidth_or_149_cse , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1295_nl = MUX1HOT_v_21_7_2((z_out_1049_29_7[22:2]),
      (z_out_1072_29_7[22:2]), (z_out_950_29_7[22:2]), (z_out_857_29_7[22:2]), (z_out_888_29_7[22:2]),
      (z_out_952_29_7[22:2]), (z_out_1152_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_708 = conv_s2u_21_22(AccumDotWidth_mux1h_1294_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1295_nl);
  assign z_out_708 = nl_z_out_708[21:0];
  assign AccumDotWidth_mux1h_1296_nl = MUX1HOT_v_21_7_2((z_out_1092_29_7[22:2]),
      (z_out_1007_29_7[22:2]), (z_out_969_29_7[22:2]), (z_out_1001_29_7[22:2]), (z_out_910_29_7[22:2]),
      (z_out_1056_29_7[22:2]), (z_out_987_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1297_nl = MUX1HOT_v_21_6_2((z_out_1103_29_7[22:2]),
      (z_out_1050_29_7[22:2]), (z_out_866_29_7[22:2]), (z_out_894_29_7[22:2]), (z_out_1086_29_7[22:2]),
      (z_out_1183_29_7[22:2]), {AccumDotWidth_or_153_cse , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign nl_z_out_709 = conv_s2u_21_22(AccumDotWidth_mux1h_1296_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1297_nl);
  assign z_out_709 = nl_z_out_709[21:0];
  assign AccumDotWidth_mux1h_1298_nl = MUX1HOT_v_21_7_2((z_out_853_29_7[22:2]), z_out_1067_29_9,
      (z_out_994_29_7[22:2]), (z_out_1093_29_7[22:2]), (z_out_1101_29_7[22:2]), (z_out_887_29_7[22:2]),
      z_out_963_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1299_nl = MUX1HOT_v_21_7_2(z_out_992_29_9, z_out_1059_29_9,
      (z_out_1035_29_7[22:2]), (z_out_1186_29_7[22:2]), (z_out_1161_29_7[22:2]),
      z_out_1066_29_9, (z_out_1184_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_710 = conv_s2u_21_22(AccumDotWidth_mux1h_1298_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1299_nl);
  assign z_out_710 = nl_z_out_710[21:0];
  assign AccumDotWidth_mux1h_1300_nl = MUX1HOT_v_21_7_2(z_out_1065_29_9, (z_out_568_29_7[22:2]),
      (z_out_975_29_7[22:2]), (z_out_952_29_7[22:2]), (z_out_573_29_7[22:2]), z_out_993_29_9,
      z_out_1140_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1301_nl = MUX1HOT_v_21_7_2((z_out_889_29_7[22:2]), (z_out_574_29_7[22:2]),
      (z_out_868_29_7[22:2]), (z_out_1073_29_7[22:2]), (z_out_997_29_7[22:2]), z_out_1006_29_9,
      z_out_978_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_711 = conv_s2u_21_22(AccumDotWidth_mux1h_1300_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1301_nl);
  assign z_out_711 = nl_z_out_711[21:0];
  assign AccumDotWidth_mux1h_1302_nl = MUX1HOT_v_21_7_2((z_out_971_29_7[22:2]), z_out_1144_29_9,
      (z_out_1167_29_7[22:2]), (z_out_934_29_7[22:2]), (z_out_871_29_7[22:2]), (z_out_935_29_7[22:2]),
      (z_out_1162_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1303_nl = MUX1HOT_v_21_7_2((z_out_901_29_7[22:2]), (z_out_1130_29_7[22:2]),
      (z_out_1093_29_7[22:2]), (z_out_938_29_7[22:2]), (z_out_968_29_7[22:2]), (z_out_613_29_7[22:2]),
      (z_out_1082_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_712 = conv_s2u_21_22(AccumDotWidth_mux1h_1302_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1303_nl);
  assign z_out_712 = nl_z_out_712[21:0];
  assign AccumDotWidth_mux1h_1304_nl = MUX1HOT_v_21_7_2((z_out_982_29_7[22:2]), (z_out_1165_29_7[22:2]),
      (z_out_937_29_7[22:2]), (z_out_872_29_7[22:2]), (z_out_1106_29_7[22:2]), (z_out_956_29_7[22:2]),
      (z_out_624_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1305_nl = MUX1HOT_v_21_7_2((z_out_624_29_7[22:2]), (z_out_1163_29_7[22:2]),
      (z_out_1073_29_7[22:2]), (z_out_1027_29_7[22:2]), (z_out_1119_29_7[22:2]),
      (z_out_987_29_7[22:2]), z_out_1046_29_9, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_713 = conv_s2u_21_22(AccumDotWidth_mux1h_1304_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1305_nl);
  assign z_out_713 = nl_z_out_713[21:0];
  assign AccumDotWidth_mux1h_1306_nl = MUX1HOT_v_21_7_2((z_out_941_29_7[22:2]), z_out_1142_29_9,
      (z_out_955_29_7[22:2]), (z_out_1166_29_7[22:2]), (z_out_877_29_7[22:2]), (z_out_1157_29_7[22:2]),
      (z_out_869_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1307_nl = MUX1HOT_v_21_7_2(z_out_1135_29_9, (z_out_914_29_7[22:2]),
      (z_out_1105_29_7[22:2]), (z_out_1169_29_7[22:2]), (z_out_928_29_7[22:2]), (z_out_949_29_7[22:2]),
      z_out_1033_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_714 = conv_s2u_21_22(AccumDotWidth_mux1h_1306_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1307_nl);
  assign z_out_714 = nl_z_out_714[21:0];
  assign AccumDotWidth_mux1h_1308_nl = MUX1HOT_v_21_7_2(z_out_1031_29_9, (z_out_1105_29_7[22:2]),
      (z_out_1119_29_7[22:2]), (z_out_868_29_7[22:2]), (z_out_1130_29_7[22:2]), (z_out_1171_29_7[22:2]),
      z_out_1142_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1309_nl = MUX1HOT_v_21_7_2(z_out_1020_29_9, (z_out_1107_29_7[22:2]),
      (z_out_911_29_7[22:2]), (z_out_1030_29_7[22:2]), (z_out_990_29_7[22:2]), (z_out_921_29_7[22:2]),
      (z_out_1154_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_715 = conv_s2u_21_22(AccumDotWidth_mux1h_1308_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1309_nl);
  assign z_out_715 = nl_z_out_715[21:0];
  assign AccumDotWidth_mux1h_1310_nl = MUX1HOT_v_21_7_2((z_out_884_29_7[22:2]), (z_out_1095_29_7[22:2]),
      (z_out_940_29_7[22:2]), (z_out_928_29_7[22:2]), z_out_1132_29_9, (z_out_1151_29_7[22:2]),
      (z_out_1105_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1311_nl = MUX1HOT_v_21_7_2((z_out_615_29_7[22:2]), z_out_1143_29_9,
      (z_out_855_29_7[22:2]), (z_out_918_29_7[22:2]), (z_out_1121_29_7[22:2]), (z_out_953_29_7[22:2]),
      (z_out_1158_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_716 = conv_s2u_21_22(AccumDotWidth_mux1h_1310_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1311_nl);
  assign z_out_716 = nl_z_out_716[21:0];
  assign AccumDotWidth_mux1h_1312_nl = MUX1HOT_v_21_6_2((z_out_1026_29_7[22:2]),
      (z_out_1131_29_7[22:2]), (z_out_1182_29_7[22:2]), (z_out_595_29_7[22:2]), (z_out_1166_29_7[22:2]),
      (z_out_1000_29_7[22:2]), {(fsm_output[2]) , AccumDotWidth_or_132_cse_1 , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1313_nl = MUX1HOT_v_21_7_2(z_out_1018_29_9, (z_out_1077_29_7[22:2]),
      (z_out_1159_29_7[22:2]), (z_out_1009_29_7[22:2]), (z_out_1116_29_7[22:2]),
      (z_out_919_29_7[22:2]), (z_out_1078_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_717 = conv_s2u_21_22(AccumDotWidth_mux1h_1312_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1313_nl);
  assign z_out_717 = nl_z_out_717[21:0];
  assign AccumDotWidth_mux1h_1314_nl = MUX1HOT_v_21_7_2((z_out_1040_29_7[22:2]),
      z_out_1132_29_9, (z_out_620_29_7[22:2]), (z_out_871_29_7[22:2]), (z_out_1129_29_7[22:2]),
      (z_out_874_29_7[22:2]), (z_out_861_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1315_nl = MUX1HOT_v_21_7_2((z_out_905_29_7[22:2]), (z_out_1106_29_7[22:2]),
      z_out_1048_29_9, (z_out_1029_29_7[22:2]), (z_out_1011_29_7[22:2]), (z_out_617_29_7[22:2]),
      (z_out_918_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_718 = conv_s2u_21_22(AccumDotWidth_mux1h_1314_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1315_nl);
  assign z_out_718 = nl_z_out_718[21:0];
  assign AccumDotWidth_mux1h_1316_nl = MUX1HOT_v_21_7_2((z_out_1036_29_7[22:2]),
      (z_out_601_29_7[22:2]), (z_out_920_29_7[22:2]), (z_out_1172_29_7[22:2]), (z_out_867_29_7[22:2]),
      (z_out_860_29_7[22:2]), (z_out_858_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1317_nl = MUX1HOT_v_21_7_2((z_out_899_29_7[22:2]), (z_out_596_29_7[22:2]),
      (z_out_1068_29_7[22:2]), z_out_1065_29_9, (z_out_883_29_7[22:2]), (z_out_977_29_7[22:2]),
      (z_out_920_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_719 = conv_s2u_21_22(AccumDotWidth_mux1h_1316_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1317_nl);
  assign z_out_719 = nl_z_out_719[21:0];
  assign AccumDotWidth_mux1h_1318_nl = MUX1HOT_v_21_7_2((z_out_1039_29_7[22:2]),
      (z_out_599_29_7[22:2]), (z_out_958_29_7[22:2]), (z_out_936_29_7[22:2]), (z_out_1070_29_7[22:2]),
      (z_out_902_29_7[22:2]), (z_out_1175_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1319_nl = MUX1HOT_v_21_7_2((z_out_576_29_7[22:2]), (z_out_589_29_7[22:2]),
      z_out_1132_29_9, (z_out_917_29_7[22:2]), (z_out_1178_29_7[22:2]), (z_out_1077_29_7[22:2]),
      (z_out_1079_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_720 = conv_s2u_21_22(AccumDotWidth_mux1h_1318_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1319_nl);
  assign z_out_720 = nl_z_out_720[21:0];
  assign AccumDotWidth_mux1h_1320_nl = MUX1HOT_v_21_7_2((z_out_872_29_7[22:2]), (z_out_600_29_7[22:2]),
      (z_out_1120_29_7[22:2]), (z_out_1077_29_7[22:2]), (z_out_1098_29_7[22:2]),
      (z_out_892_29_7[22:2]), (z_out_1055_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1321_nl = MUX1HOT_v_21_7_2((z_out_923_29_7[22:2]), (z_out_598_29_7[22:2]),
      (z_out_916_29_7[22:2]), (z_out_1011_29_7[22:2]), (z_out_624_29_7[22:2]), (z_out_579_29_7[22:2]),
      (z_out_1026_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_721 = conv_s2u_21_22(AccumDotWidth_mux1h_1320_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1321_nl);
  assign z_out_721 = nl_z_out_721[21:0];
  assign AccumDotWidth_mux1h_1322_nl = MUX1HOT_v_21_7_2((z_out_1094_29_7[22:2]),
      (z_out_918_29_7[22:2]), (z_out_946_29_7[22:2]), (z_out_1105_29_7[22:2]), (z_out_1058_29_7[22:2]),
      (z_out_890_29_7[22:2]), (z_out_1001_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1323_nl = MUX1HOT_v_21_7_2((z_out_1099_29_7[22:2]),
      z_out_1059_29_9, (z_out_859_29_7[22:2]), (z_out_1014_29_7[22:2]), (z_out_954_29_7[22:2]),
      (z_out_1026_29_7[22:2]), (z_out_606_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_722 = conv_s2u_21_22(AccumDotWidth_mux1h_1322_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1323_nl);
  assign z_out_722 = nl_z_out_722[21:0];
  assign AccumDotWidth_mux1h_1324_nl = MUX1HOT_v_21_7_2((z_out_983_29_7[22:2]), (z_out_629_29_7[22:2]),
      (z_out_896_29_7[22:2]), (z_out_922_29_7[22:2]), (z_out_602_29_7[22:2]), (z_out_893_29_7[22:2]),
      (z_out_907_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1325_nl = MUX1HOT_v_21_7_2((z_out_625_29_7[22:2]), (z_out_619_29_7[22:2]),
      (z_out_1158_29_7[22:2]), (z_out_853_29_7[22:2]), (z_out_1115_29_7[22:2]), z_out_1140_29_9,
      (z_out_589_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_723 = conv_s2u_21_22(AccumDotWidth_mux1h_1324_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1325_nl);
  assign z_out_723 = nl_z_out_723[21:0];
  assign AccumDotWidth_mux1h_1326_nl = MUX1HOT_v_21_7_2((z_out_903_29_7[22:2]), (z_out_1094_29_7[22:2]),
      z_out_1141_29_9, (z_out_1002_29_7[22:2]), (z_out_1055_29_7[22:2]), (z_out_1079_29_7[22:2]),
      (z_out_619_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1327_nl = MUX1HOT_v_21_7_2((z_out_951_29_7[22:2]), (z_out_902_29_7[22:2]),
      (z_out_593_29_7[22:2]), (z_out_863_29_7[22:2]), z_out_963_29_9, (z_out_1074_29_7[22:2]),
      (z_out_1044_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_724 = conv_s2u_21_22(AccumDotWidth_mux1h_1326_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1327_nl);
  assign z_out_724 = nl_z_out_724[21:0];
  assign AccumDotWidth_mux1h_1328_nl = MUX1HOT_v_21_7_2(z_out_1048_29_9, (z_out_1170_29_7[22:2]),
      z_out_1138_29_9, (z_out_987_29_7[22:2]), (z_out_1036_29_7[22:2]), (z_out_1182_29_7[22:2]),
      (z_out_966_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1329_nl = MUX1HOT_v_21_7_2((z_out_1042_29_7[22:2]),
      (z_out_1081_29_7[22:2]), (z_out_1187_29_7[22:2]), (z_out_1041_29_7[22:2]),
      (z_out_927_29_7[22:2]), z_out_1018_29_9, (z_out_1130_29_7[22:2]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_725 = conv_s2u_21_22(AccumDotWidth_mux1h_1328_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1329_nl);
  assign z_out_725 = nl_z_out_725[21:0];
  assign AccumDotWidth_mux1h_1330_nl = MUX1HOT_v_21_7_2((z_out_1178_29_7[22:2]),
      (z_out_909_29_7[22:2]), (z_out_1161_29_7[22:2]), (z_out_883_29_7[22:2]), (z_out_576_29_7[22:2]),
      (z_out_858_29_7[22:2]), (z_out_901_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1331_nl = MUX1HOT_v_21_7_2((z_out_916_29_7[22:2]), (z_out_922_29_7[22:2]),
      (z_out_1185_29_7[22:2]), (z_out_1026_29_7[22:2]), z_out_965_29_9, (z_out_970_29_7[22:2]),
      (z_out_582_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_726 = conv_s2u_21_22(AccumDotWidth_mux1h_1330_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1331_nl);
  assign z_out_726 = nl_z_out_726[21:0];
  assign AccumDotWidth_mux1h_1332_nl = MUX1HOT_v_21_6_2((z_out_1101_29_7[22:2]),
      (z_out_1164_29_7[22:2]), (z_out_1038_29_7[22:2]), (z_out_1015_29_7[22:2]),
      z_out_1137_29_9, (z_out_991_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , AccumDotWidth_or_140_cse});
  assign AccumDotWidth_mux1h_1333_nl = MUX1HOT_v_21_7_2((z_out_966_29_7[22:2]), (z_out_1166_29_7[22:2]),
      (z_out_938_29_7[22:2]), (z_out_1086_29_7[22:2]), (z_out_1120_29_7[22:2]), (z_out_883_29_7[22:2]),
      (z_out_1038_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_727 = conv_s2u_21_22(AccumDotWidth_mux1h_1332_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1333_nl);
  assign z_out_727 = nl_z_out_727[21:0];
  assign AccumDotWidth_mux1h_1334_nl = MUX1HOT_v_21_7_2((z_out_863_29_7[22:2]), (z_out_1168_29_7[22:2]),
      z_out_992_29_9, (z_out_1074_29_7[22:2]), (z_out_577_29_7[22:2]), (z_out_1117_29_7[22:2]),
      (z_out_889_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1335_nl = MUX1HOT_v_21_7_2((z_out_887_29_7[22:2]), (z_out_911_29_7[22:2]),
      (z_out_602_29_7[22:2]), (z_out_583_29_7[22:2]), z_out_962_29_9, (z_out_1126_29_7[22:2]),
      (z_out_1029_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_728 = conv_s2u_21_22(AccumDotWidth_mux1h_1334_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1335_nl);
  assign z_out_728 = nl_z_out_728[21:0];
  assign AccumDotWidth_mux1h_1336_nl = MUX1HOT_v_21_7_2((z_out_606_29_7[22:2]), (z_out_910_29_7[22:2]),
      z_out_1065_29_9, (z_out_1019_29_7[22:2]), (z_out_973_29_7[22:2]), (z_out_997_29_7[22:2]),
      (z_out_1072_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1337_nl = MUX1HOT_v_21_7_2((z_out_1078_29_7[22:2]),
      (z_out_921_29_7[22:2]), (z_out_924_29_7[22:2]), (z_out_976_29_7[22:2]), (z_out_879_29_7[22:2]),
      (z_out_915_29_7[22:2]), (z_out_1110_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_729 = conv_s2u_21_22(AccumDotWidth_mux1h_1336_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1337_nl);
  assign z_out_729 = nl_z_out_729[21:0];
  assign AccumDotWidth_mux1h_1338_nl = MUX1HOT_v_21_7_2((z_out_859_29_7[22:2]), (z_out_1171_29_7[22:2]),
      (z_out_945_29_7[22:2]), (z_out_920_29_7[22:2]), (z_out_1040_29_7[22:2]), (z_out_625_29_7[22:2]),
      (z_out_890_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1339_nl = MUX1HOT_v_21_7_2((z_out_587_29_7[22:2]), (z_out_1170_29_7[22:2]),
      (z_out_857_29_7[22:2]), (z_out_1179_29_7[22:2]), (z_out_1051_29_7[22:2]), (z_out_1043_29_7[22:2]),
      (z_out_1024_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_730 = conv_s2u_21_22(AccumDotWidth_mux1h_1338_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1339_nl);
  assign z_out_730 = nl_z_out_730[21:0];
  assign AccumDotWidth_mux1h_1340_nl = MUX1HOT_v_21_7_2((z_out_1043_29_7[22:2]),
      (z_out_595_29_7[22:2]), (z_out_599_29_7[22:2]), (z_out_1165_29_7[22:2]), (z_out_1092_29_7[22:2]),
      z_out_1061_29_9, (z_out_1115_29_7[22:2]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1341_nl = MUX1HOT_v_21_7_2((z_out_1036_29_7[22:2]),
      (z_out_1053_29_7[22:2]), (z_out_892_29_7[22:2]), (z_out_971_29_7[22:2]), (z_out_951_29_7[22:2]),
      (z_out_1094_29_7[22:2]), (z_out_977_29_7[22:2]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_731 = conv_s2u_21_22(AccumDotWidth_mux1h_1340_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1341_nl);
  assign z_out_731 = nl_z_out_731[21:0];
  assign AccumDotWidth_mux1h_1342_nl = MUX1HOT_v_21_7_2((z_out_1044_29_7[22:2]),
      (z_out_1098_29_7[22:2]), (z_out_1153_29_7[22:2]), (z_out_1145_29_7[22:2]),
      (z_out_571_29_7[22:2]), (z_out_570_29_7[22:2]), (z_out_1166_29_7[22:2]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1343_nl = MUX1HOT_v_21_7_2(z_out_1047_29_9, (z_out_1181_29_7[22:2]),
      (z_out_929_29_7[22:2]), z_out_1139_29_9, (z_out_1000_29_7[22:2]), (z_out_1156_29_7[22:2]),
      (z_out_912_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_732 = conv_s2u_21_22(AccumDotWidth_mux1h_1342_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1343_nl);
  assign z_out_732 = nl_z_out_732[21:0];
  assign AccumDotWidth_mux1h_1344_nl = MUX1HOT_v_21_7_2((z_out_885_29_7[22:2]), (z_out_1023_29_7[22:2]),
      (z_out_1008_29_7[22:2]), (z_out_972_29_7[22:2]), (z_out_1105_29_7[22:2]), (z_out_1106_29_7[22:2]),
      (z_out_1161_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1345_nl = MUX1HOT_v_21_7_2((z_out_886_29_7[22:2]), (z_out_1183_29_7[22:2]),
      (z_out_871_29_7[22:2]), (z_out_1184_29_7[22:2]), (z_out_1049_29_7[22:2]), z_out_978_29_9,
      (z_out_922_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_733 = conv_s2u_21_22(AccumDotWidth_mux1h_1344_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1345_nl);
  assign z_out_733 = nl_z_out_733[21:0];
  assign AccumDotWidth_mux1h_1346_nl = MUX1HOT_v_21_7_2((z_out_887_29_7[22:2]), (z_out_958_29_7[22:2]),
      (z_out_1154_29_7[22:2]), (z_out_1085_29_7[22:2]), z_out_1047_29_9, (z_out_1176_29_7[22:2]),
      (z_out_1149_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1347_nl = MUX1HOT_v_21_7_2((z_out_883_29_7[22:2]), (z_out_906_29_7[22:2]),
      (z_out_990_29_7[22:2]), (z_out_860_29_7[22:2]), (z_out_866_29_7[22:2]), (z_out_1016_29_7[22:2]),
      (z_out_943_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_734 = conv_s2u_21_22(AccumDotWidth_mux1h_1346_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1347_nl);
  assign z_out_734 = nl_z_out_734[21:0];
  assign AccumDotWidth_mux1h_1348_nl = MUX1HOT_v_21_6_2((z_out_1040_29_7[22:2]),
      (z_out_1150_29_7[22:2]), z_out_1004_29_9, (z_out_1021_29_7[22:2]), (z_out_1167_29_7[22:2]),
      (z_out_1157_29_7[22:2]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1349_nl = MUX1HOT_v_21_5_2((z_out_1039_29_7[22:2]),
      (z_out_953_29_7[22:2]), (z_out_864_29_7[22:2]), (z_out_1058_29_7[22:2]), (z_out_1089_29_7[22:2]),
      {(fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[2]) ,
      (fsm_output[6])});
  assign nl_z_out_735 = conv_s2u_21_22(AccumDotWidth_mux1h_1348_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1349_nl);
  assign z_out_735 = nl_z_out_735[21:0];
  assign AccumDotWidth_mux1h_1350_nl = MUX1HOT_v_21_7_2((z_out_882_29_7[22:2]), (z_out_964_29_7[22:2]),
      (z_out_582_29_7[22:2]), z_out_965_29_9, (z_out_1042_29_7[22:2]), (z_out_1095_29_7[22:2]),
      (z_out_629_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1351_nl = MUX1HOT_v_21_7_2((z_out_881_29_7[22:2]), (z_out_579_29_7[22:2]),
      (z_out_611_29_7[22:2]), (z_out_1121_29_7[22:2]), (z_out_1054_29_7[22:2]), (z_out_976_29_7[22:2]),
      (z_out_1043_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_736 = conv_s2u_21_22(AccumDotWidth_mux1h_1350_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1351_nl);
  assign z_out_736 = nl_z_out_736[21:0];
  assign AccumDotWidth_mux1h_1352_nl = MUX1HOT_v_21_7_2((z_out_889_29_7[22:2]), z_out_963_29_9,
      (z_out_973_29_7[22:2]), (z_out_1128_29_7[22:2]), (z_out_1156_29_7[22:2]), (z_out_569_29_7[22:2]),
      (z_out_1148_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1353_nl = MUX1HOT_v_21_7_2((z_out_890_29_7[22:2]), (z_out_894_29_7[22:2]),
      (z_out_1034_29_7[22:2]), (z_out_912_29_7[22:2]), (z_out_925_29_7[22:2]), (z_out_1187_29_7[22:2]),
      (z_out_946_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_737 = conv_s2u_21_22(AccumDotWidth_mux1h_1352_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1353_nl);
  assign z_out_737 = nl_z_out_737[21:0];
  assign AccumDotWidth_mux1h_1354_nl = MUX1HOT_v_21_7_2((z_out_880_29_7[22:2]), (z_out_602_29_7[22:2]),
      (z_out_997_29_7[22:2]), (z_out_999_29_7[22:2]), (z_out_1111_29_7[22:2]), (z_out_1050_29_7[22:2]),
      (z_out_1160_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1355_nl = MUX1HOT_v_21_6_2((z_out_888_29_7[22:2]), (z_out_1091_29_7[22:2]),
      z_out_1006_29_9, z_out_1138_29_9, (z_out_1102_29_7[22:2]), (z_out_916_29_7[22:2]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_738 = conv_s2u_21_22(AccumDotWidth_mux1h_1354_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1355_nl);
  assign z_out_738 = nl_z_out_738[21:0];
  assign AccumDotWidth_mux1h_1356_nl = MUX1HOT_v_21_6_2((z_out_884_29_7[22:2]), (z_out_1100_29_7[22:2]),
      z_out_1047_29_9, (z_out_1146_29_7[22:2]), (z_out_931_29_7[22:2]), (z_out_955_29_7[22:2]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1357_nl = MUX1HOT_v_21_6_2((z_out_1158_29_7[22:2]),
      (z_out_1184_29_7[22:2]), (z_out_1022_29_7[22:2]), (z_out_946_29_7[22:2]), (z_out_950_29_7[22:2]),
      (z_out_1180_29_7[22:2]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_739 = conv_s2u_21_22(AccumDotWidth_mux1h_1356_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1357_nl);
  assign z_out_739 = nl_z_out_739[21:0];
  assign AccumDotWidth_mux1h_1358_nl = MUX1HOT_v_21_6_2((z_out_1005_29_7[22:2]),
      z_out_1133_29_9, (z_out_999_29_7[22:2]), (z_out_915_29_7[22:2]), (z_out_1168_29_7[22:2]),
      (z_out_1040_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1359_nl = MUX1HOT_v_21_6_2((z_out_580_29_7[22:2]), (z_out_1129_29_7[22:2]),
      (z_out_1049_29_7[22:2]), (z_out_858_29_7[22:2]), (z_out_1091_29_7[22:2]), (z_out_876_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_740 = conv_s2u_21_22(AccumDotWidth_mux1h_1358_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1359_nl);
  assign z_out_740 = nl_z_out_740[21:0];
  assign AccumDotWidth_mux1h_1360_nl = MUX1HOT_v_21_6_2((z_out_1002_29_7[22:2]),
      (z_out_1109_29_7[22:2]), (z_out_998_29_7[22:2]), (z_out_990_29_7[22:2]), (z_out_994_29_7[22:2]),
      (z_out_1039_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1361_nl = MUX1HOT_v_21_6_2((z_out_879_29_7[22:2]), (z_out_1122_29_7[22:2]),
      (z_out_863_29_7[22:2]), (z_out_1068_29_7[22:2]), (z_out_880_29_7[22:2]), (z_out_1002_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_741 = conv_s2u_21_22(AccumDotWidth_mux1h_1360_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1361_nl);
  assign z_out_741 = nl_z_out_741[21:0];
  assign AccumDotWidth_mux1h_1362_nl = MUX1HOT_v_21_6_2((z_out_1171_29_7[22:2]),
      (z_out_856_29_7[22:2]), (z_out_947_29_7[22:2]), (z_out_1049_29_7[22:2]), (z_out_909_29_7[22:2]),
      (z_out_954_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1363_nl = MUX1HOT_v_21_6_2((z_out_1030_29_7[22:2]),
      (z_out_855_29_7[22:2]), (z_out_861_29_7[22:2]), (z_out_1079_29_7[22:2]), (z_out_891_29_7[22:2]),
      (z_out_1185_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_742 = conv_s2u_21_22(AccumDotWidth_mux1h_1362_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1363_nl);
  assign z_out_742 = nl_z_out_742[21:0];
  assign AccumDotWidth_mux1h_1364_nl = MUX1HOT_v_21_6_2((z_out_1164_29_7[22:2]),
      (z_out_588_29_7[22:2]), z_out_1004_29_9, (z_out_1094_29_7[22:2]), z_out_1144_29_9,
      (z_out_1049_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1365_nl = MUX1HOT_v_21_6_2((z_out_1025_29_7[22:2]),
      (z_out_594_29_7[22:2]), (z_out_1165_29_7[22:2]), z_out_1188_29_9, (z_out_1045_29_7[22:2]),
      z_out_1067_29_9, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_743 = conv_s2u_21_22(AccumDotWidth_mux1h_1364_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1365_nl);
  assign z_out_743 = nl_z_out_743[21:0];
  assign AccumDotWidth_mux1h_1366_nl = MUX1HOT_v_21_6_2((z_out_885_29_7[22:2]), (z_out_590_29_7[22:2]),
      (z_out_1168_29_7[22:2]), (z_out_996_29_7[22:2]), (z_out_1169_29_7[22:2]), (z_out_1036_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1367_nl = MUX1HOT_v_21_6_2((z_out_616_29_7[22:2]), (z_out_586_29_7[22:2]),
      (z_out_1019_29_7[22:2]), (z_out_626_29_7[22:2]), (z_out_930_29_7[22:2]), (z_out_873_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_744 = conv_s2u_21_22(AccumDotWidth_mux1h_1366_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1367_nl);
  assign z_out_744 = nl_z_out_744[21:0];
  assign AccumDotWidth_mux1h_1368_nl = MUX1HOT_v_21_6_2((z_out_1161_29_7[22:2]),
      z_out_1134_29_9, (z_out_917_29_7[22:2]), (z_out_921_29_7[22:2]), (z_out_1146_29_7[22:2]),
      (z_out_595_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1369_nl = MUX1HOT_v_21_6_2((z_out_1029_29_7[22:2]),
      (z_out_1127_29_7[22:2]), (z_out_1069_29_7[22:2]), (z_out_855_29_7[22:2]), (z_out_1175_29_7[22:2]),
      (z_out_1015_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_745 = conv_s2u_21_22(AccumDotWidth_mux1h_1368_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1369_nl);
  assign z_out_745 = nl_z_out_745[21:0];
  assign AccumDotWidth_mux1h_1370_nl = MUX1HOT_v_21_6_2((z_out_1155_29_7[22:2]),
      (z_out_1123_29_7[22:2]), (z_out_915_29_7[22:2]), (z_out_1007_29_7[22:2]), (z_out_568_29_7[22:2]),
      (z_out_1064_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1371_nl = MUX1HOT_v_21_6_2(z_out_1140_29_9, (z_out_1128_29_7[22:2]),
      (z_out_858_29_7[22:2]), (z_out_1078_29_7[22:2]), (z_out_995_29_7[22:2]), (z_out_1051_29_7[22:2]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign nl_z_out_746 = conv_s2u_21_22(AccumDotWidth_mux1h_1370_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1371_nl);
  assign z_out_746 = nl_z_out_746[21:0];
  assign AccumDotWidth_mux1h_1372_nl = MUX1HOT_v_21_5_2(z_out_1003_29_9, (z_out_1108_29_7[22:2]),
      (z_out_1097_29_7[22:2]), (z_out_972_29_7[22:2]), (z_out_604_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1373_nl = MUX1HOT_v_21_5_2((z_out_878_29_7[22:2]), z_out_1140_29_9,
      (z_out_1185_29_7[22:2]), z_out_942_29_9, (z_out_1011_29_7[22:2]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_747 = conv_s2u_21_22(AccumDotWidth_mux1h_1372_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1373_nl);
  assign z_out_747 = nl_z_out_747[21:0];
  assign AccumDotWidth_mux1h_1374_nl = MUX1HOT_v_21_4_2((z_out_1148_29_7[22:2]),
      (z_out_593_29_7[22:2]), (z_out_1036_29_7[22:2]), z_out_962_29_9, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[7])});
  assign AccumDotWidth_mux1h_1375_nl = MUX1HOT_v_21_4_2((z_out_588_29_7[22:2]), (z_out_587_29_7[22:2]),
      (z_out_908_29_7[22:2]), (z_out_1179_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_748 = conv_s2u_21_22(AccumDotWidth_mux1h_1374_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1375_nl);
  assign z_out_748 = nl_z_out_748[21:0];
  assign AccumDotWidth_mux1h_1376_nl = MUX1HOT_v_21_3_2((z_out_1153_29_7[22:2]),
      (z_out_591_29_7[22:2]), (z_out_1098_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1377_nl = MUX1HOT_v_21_3_2((z_out_585_29_7[22:2]), (z_out_1126_29_7[22:2]),
      (z_out_627_29_7[22:2]), {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6])});
  assign nl_z_out_749 = conv_s2u_21_22(AccumDotWidth_mux1h_1376_nl) + conv_s2u_21_22(AccumDotWidth_mux1h_1377_nl);
  assign z_out_749 = nl_z_out_749[21:0];
  assign AccumDotWidth_mux_143_nl = MUX_v_21_2_2((z_out_1044_29_7[22:2]), (z_out_1122_29_7[22:2]),
      fsm_output[6]);
  assign AccumDotWidth_mux_144_nl = MUX_v_21_2_2((z_out_581_29_7[22:2]), (z_out_1009_29_7[22:2]),
      fsm_output[6]);
  assign nl_z_out_750 = conv_s2u_21_22(AccumDotWidth_mux_143_nl) + conv_s2u_21_22(AccumDotWidth_mux_144_nl);
  assign z_out_750 = nl_z_out_750[21:0];
  assign AccumDotWidth_mux1h_1378_nl = MUX1HOT_v_22_7_2(z_out_237, z_out_471, z_out_269,
      z_out_543, z_out_826, z_out_565, z_out_274, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1379_nl = MUX1HOT_v_22_7_2(z_out_320, z_out_469, z_out_519,
      z_out_237, z_out_319, z_out_513, z_out_273, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_751 = (AccumDotWidth_mux1h_1378_nl) + (AccumDotWidth_mux1h_1379_nl);
  assign z_out_751 = nl_z_out_751[21:0];
  assign nl_MultLoop_acc_1611_nl = (z_out_889_29_7[21:0]) + (z_out_890_29_7[21:0]);
  assign MultLoop_acc_1611_nl = nl_MultLoop_acc_1611_nl[21:0];
  assign nl_MultLoop_acc_1612_nl = (z_out_879_29_7[21:0]) + (z_out_911_29_7[21:0]);
  assign MultLoop_acc_1612_nl = nl_MultLoop_acc_1612_nl[21:0];
  assign nl_MultLoop_acc_1610_nl = (MultLoop_acc_1611_nl) + (MultLoop_acc_1612_nl);
  assign MultLoop_acc_1610_nl = nl_MultLoop_acc_1610_nl[21:0];
  assign nl_MultLoop_acc_1609_nl = (MultLoop_acc_1610_nl) + z_out_517;
  assign MultLoop_acc_1609_nl = nl_MultLoop_acc_1609_nl[21:0];
  assign AccumDotWidth_mux1h_1380_nl = MUX1HOT_v_22_6_2(z_out_317, z_out_535, z_out_460,
      z_out_453, z_out_325, (MultLoop_acc_1609_nl), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1613_nl = z_out_516 + z_out_515;
  assign MultLoop_acc_1613_nl = nl_MultLoop_acc_1613_nl[21:0];
  assign AccumDotWidth_mux1h_1381_nl = MUX1HOT_v_22_6_2(z_out_318, z_out_534, z_out_285,
      z_out_565, z_out_238, (MultLoop_acc_1613_nl), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_752 = (AccumDotWidth_mux1h_1380_nl) + (AccumDotWidth_mux1h_1381_nl);
  assign z_out_752 = nl_z_out_752[21:0];
  assign MultLoop_mux1h_507_nl = MUX1HOT_v_22_3_2(z_out_448, z_out_44_28_7, z_out_127_28_7,
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign MultLoop_mux1h_508_nl = MUX1HOT_v_22_3_2(z_out_449, z_out_34_28_7, z_out_76_28_7,
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_753 = (MultLoop_mux1h_507_nl) + (MultLoop_mux1h_508_nl);
  assign z_out_753 = nl_z_out_753[21:0];
  assign nl_MultLoop_acc_1616_nl = (z_out_1183_29_7[21:0]) + MultLoop_193_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1616_nl = nl_MultLoop_acc_1616_nl[21:0];
  assign nl_MultLoop_acc_1617_nl = (z_out_1181_29_7[21:0]) + (z_out_1171_29_7[21:0]);
  assign MultLoop_acc_1617_nl = nl_MultLoop_acc_1617_nl[21:0];
  assign nl_MultLoop_acc_1614_nl = MultLoop_acc_89_itm + (MultLoop_acc_1616_nl) +
      (MultLoop_acc_1617_nl);
  assign MultLoop_acc_1614_nl = nl_MultLoop_acc_1614_nl[21:0];
  assign AccumDotWidth_mux1h_1382_nl = MUX1HOT_v_22_3_2(z_out_529, z_out_458, (MultLoop_acc_1614_nl),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1383_nl = MUX1HOT_v_22_3_2(z_out_531, z_out_511, MultLoop_acc_113_itm,
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_754 = (AccumDotWidth_mux1h_1382_nl) + (AccumDotWidth_mux1h_1383_nl);
  assign z_out_754 = nl_z_out_754[21:0];
  assign nl_MultLoop_acc_1620_nl = z_out_192_28_7 + z_out_191_28_7;
  assign MultLoop_acc_1620_nl = nl_MultLoop_acc_1620_nl[21:0];
  assign nl_MultLoop_acc_1621_nl = z_out_190_28_7 + z_out_189_28_7;
  assign MultLoop_acc_1621_nl = nl_MultLoop_acc_1621_nl[21:0];
  assign nl_MultLoop_acc_1619_nl = (MultLoop_acc_1620_nl) + (MultLoop_acc_1621_nl);
  assign MultLoop_acc_1619_nl = nl_MultLoop_acc_1619_nl[21:0];
  assign nl_MultLoop_acc_1618_nl = z_out_565 + (MultLoop_acc_1619_nl);
  assign MultLoop_acc_1618_nl = nl_MultLoop_acc_1618_nl[21:0];
  assign AccumDotWidth_mux1h_1384_nl = MUX1HOT_v_22_6_2(z_out_536, z_out_269, z_out_540,
      z_out_519, z_out_463, (MultLoop_acc_1618_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1624_nl = z_out_677_28_7 + z_out_678_28_7;
  assign MultLoop_acc_1624_nl = nl_MultLoop_acc_1624_nl[21:0];
  assign nl_MultLoop_acc_1625_nl = z_out_166_28_7 + z_out_167_28_7;
  assign MultLoop_acc_1625_nl = nl_MultLoop_acc_1625_nl[21:0];
  assign nl_MultLoop_acc_1627_nl = z_out_158_28_7 + z_out_159_28_7;
  assign MultLoop_acc_1627_nl = nl_MultLoop_acc_1627_nl[21:0];
  assign nl_MultLoop_acc_1628_nl = z_out_156_28_7 + z_out_679_28_7;
  assign MultLoop_acc_1628_nl = nl_MultLoop_acc_1628_nl[21:0];
  assign nl_MultLoop_acc_1622_nl = (MultLoop_acc_1624_nl) + (MultLoop_acc_1625_nl)
      + (MultLoop_acc_1627_nl) + (MultLoop_acc_1628_nl);
  assign MultLoop_acc_1622_nl = nl_MultLoop_acc_1622_nl[21:0];
  assign AccumDotWidth_mux1h_1385_nl = MUX1HOT_v_22_6_2(z_out_527, z_out_270, z_out_518,
      z_out_522, z_out_464, (MultLoop_acc_1622_nl), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_755 = (AccumDotWidth_mux1h_1384_nl) + (AccumDotWidth_mux1h_1385_nl);
  assign z_out_755 = nl_z_out_755[21:0];
  assign AccumDotWidth_mux1h_1386_nl = MUX1HOT_v_22_7_2(z_out_530, z_out_263, z_out_264,
      z_out_539, z_out_456, z_out_518, MultLoop_acc_562_itm, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1631_nl = (z_out_972_29_7[21:0]) + (z_out_1096_29_7[21:0]);
  assign MultLoop_acc_1631_nl = nl_MultLoop_acc_1631_nl[21:0];
  assign nl_MultLoop_acc_1632_nl = (z_out_1019_29_7[21:0]) + (z_out_1005_29_7[21:0]);
  assign MultLoop_acc_1632_nl = nl_MultLoop_acc_1632_nl[21:0];
  assign nl_MultLoop_acc_1634_nl = (z_out_991_29_7[21:0]) + (z_out_967_29_7[21:0]);
  assign MultLoop_acc_1634_nl = nl_MultLoop_acc_1634_nl[21:0];
  assign nl_MultLoop_acc_1635_nl = (z_out_1007_29_7[21:0]) + (z_out_1021_29_7[21:0]);
  assign MultLoop_acc_1635_nl = nl_MultLoop_acc_1635_nl[21:0];
  assign nl_MultLoop_acc_1629_nl = (MultLoop_acc_1631_nl) + (MultLoop_acc_1632_nl)
      + (MultLoop_acc_1634_nl) + (MultLoop_acc_1635_nl);
  assign MultLoop_acc_1629_nl = nl_MultLoop_acc_1629_nl[21:0];
  assign AccumDotWidth_mux1h_1387_nl = MUX1HOT_v_22_7_2(z_out_533, z_out_528, z_out_564,
      z_out_330, z_out_510, z_out_844, (MultLoop_acc_1629_nl), {(fsm_output[1]) ,
      (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_756 = (AccumDotWidth_mux1h_1386_nl) + (AccumDotWidth_mux1h_1387_nl);
  assign z_out_756 = nl_z_out_756[21:0];
  assign MultLoop_mux1h_509_nl = MUX1HOT_v_22_3_2(MultLoop_acc_128_itm, z_out_123_28_7,
      z_out_829, {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_510_nl = MUX1HOT_v_22_3_2(z_out_437, z_out_131_28_7, z_out_827,
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_757 = (MultLoop_mux1h_509_nl) + (MultLoop_mux1h_510_nl);
  assign z_out_757 = nl_z_out_757[21:0];
  assign AccumDotWidth_mux1h_1388_nl = MUX1HOT_v_22_3_2(z_out_265, z_out_537, z_out_836,
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1389_nl = MUX1HOT_v_22_3_2(z_out_275, z_out_320, MultLoop_acc_756_itm,
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_758 = (AccumDotWidth_mux1h_1388_nl) + (AccumDotWidth_mux1h_1389_nl);
  assign z_out_758 = nl_z_out_758[21:0];
  assign nl_MultLoop_acc_1636_nl = z_out_563 + MultLoop_acc_867_itm;
  assign MultLoop_acc_1636_nl = nl_MultLoop_acc_1636_nl[21:0];
  assign AccumDotWidth_mux1h_1390_nl = MUX1HOT_v_22_7_2(z_out_835, z_out_524, z_out_270,
      z_out_323, z_out_540, z_out_519, (MultLoop_acc_1636_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1391_nl = MUX1HOT_v_22_7_2(z_out_836, z_out_525, z_out_566,
      z_out_236, z_out_508, AccumDotWidth_acc_1945_itm, MultLoop_acc_883_itm, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_759 = (AccumDotWidth_mux1h_1390_nl) + (AccumDotWidth_mux1h_1391_nl);
  assign z_out_759 = nl_z_out_759[21:0];
  assign AccumDotWidth_mux_145_nl = MUX_v_22_2_2(z_out_837, z_out_474, fsm_output[8]);
  assign AccumDotWidth_mux_146_nl = MUX_v_22_2_2(z_out_838, MultLoop_acc_377_itm,
      fsm_output[8]);
  assign nl_z_out_760 = (AccumDotWidth_mux_145_nl) + (AccumDotWidth_mux_146_nl);
  assign z_out_760 = nl_z_out_760[21:0];
  assign MultLoop_mux1h_511_nl = MUX1HOT_v_22_3_2(z_out_839, z_out_138_28_7, z_out_76_28_7,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign MultLoop_mux1h_512_nl = MUX1HOT_v_22_3_2(z_out_840, z_out_118_28_7, z_out_136_28_7,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_z_out_761 = (MultLoop_mux1h_511_nl) + (MultLoop_mux1h_512_nl);
  assign z_out_761 = nl_z_out_761[21:0];
  assign AccumDotWidth_mux1h_1392_nl = MUX1HOT_v_22_4_2(z_out_267, z_out_533, z_out_541,
      z_out_826, {(fsm_output[2]) , AccumDotWidth_or_157_cse , (fsm_output[4]) ,
      (fsm_output[8])});
  assign AccumDotWidth_mux1h_1393_nl = MUX1HOT_v_22_5_2(z_out_266, z_out_530, z_out_243,
      z_out_317, MultLoop_acc_1010_itm, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_762 = (AccumDotWidth_mux1h_1392_nl) + (AccumDotWidth_mux1h_1393_nl);
  assign z_out_762 = nl_z_out_762[21:0];
  assign AccumDotWidth_mux_147_nl = MUX_v_22_2_2(z_out_847, z_out_815, fsm_output[8]);
  assign AccumDotWidth_mux_148_nl = MUX_v_22_2_2(z_out_264, MultLoop_acc_1139_itm,
      fsm_output[8]);
  assign nl_z_out_763 = (AccumDotWidth_mux_147_nl) + (AccumDotWidth_mux_148_nl);
  assign z_out_763 = nl_z_out_763[21:0];
  assign MultLoop_mux_99_nl = MUX_v_22_2_2(z_out_455, z_out_517, fsm_output[2]);
  assign MultLoop_mux_100_nl = MUX_v_22_2_2(z_out_446, z_out_526, fsm_output[2]);
  assign nl_z_out_764 = (MultLoop_mux_99_nl) + (MultLoop_mux_100_nl);
  assign z_out_764 = nl_z_out_764[21:0];
  assign AccumDotWidth_mux1h_1394_nl = MUX1HOT_v_22_4_2(z_out_527, z_out_36_28_7,
      z_out_830, z_out_142_28_7, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign AccumDotWidth_mux1h_1395_nl = MUX1HOT_v_22_4_2(z_out_516, z_out_35_28_7,
      z_out_845, z_out_144_28_7, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[4])});
  assign nl_z_out_765 = (AccumDotWidth_mux1h_1394_nl) + (AccumDotWidth_mux1h_1395_nl);
  assign z_out_765 = nl_z_out_765[21:0];
  assign AccumDotWidth_mux1h_1396_nl = MUX1HOT_v_22_4_2(z_out_453, MultLoop_acc_628_itm,
      z_out_71_28_7, z_out_272, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[3])
      , (fsm_output[5])});
  assign AccumDotWidth_mux1h_1397_nl = MUX1HOT_v_22_4_2(z_out_454, z_out_439, z_out_70_28_7,
      z_out_277, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_766 = (AccumDotWidth_mux1h_1396_nl) + (AccumDotWidth_mux1h_1397_nl);
  assign z_out_766 = nl_z_out_766[21:0];
  assign MultLoop_mux1h_513_nl = MUX1HOT_v_22_7_2(z_out_288, z_out_449, MultLoop_acc_88_itm,
      z_out_197, z_out_220, z_out_293, z_out_224, {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_514_nl = MUX1HOT_v_22_7_2(z_out_289, z_out_218, z_out_214,
      z_out_507, z_out_495, z_out_291, z_out_219, {(fsm_output[1]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[2]) , (fsm_output[7]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_767 = (MultLoop_mux1h_513_nl) + (MultLoop_mux1h_514_nl);
  assign z_out_767 = nl_z_out_767[21:0];
  assign MultLoop_mux1h_515_nl = MUX1HOT_v_22_4_2(z_out_118_28_7, z_out_228, z_out_63_28_7,
      z_out_121_28_7, {(fsm_output[3]) , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[4])});
  assign MultLoop_mux1h_516_nl = MUX1HOT_v_22_4_2(z_out_122_28_7, z_out_227, z_out_74_28_7,
      z_out_129_28_7, {(fsm_output[3]) , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[4])});
  assign nl_z_out_768 = (MultLoop_mux1h_515_nl) + (MultLoop_mux1h_516_nl);
  assign z_out_768 = nl_z_out_768[21:0];
  assign MultLoop_mux1h_517_nl = MUX1HOT_v_22_5_2(z_out_123_28_7, z_out_456, z_out_96_28_7,
      z_out_40_28_7, z_out_134_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_518_nl = MUX1HOT_v_22_5_2(z_out_124_28_7, z_out_533, z_out_103_28_7,
      z_out_43_28_7, z_out_143_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out_769 = (MultLoop_mux1h_517_nl) + (MultLoop_mux1h_518_nl);
  assign z_out_769 = nl_z_out_769[21:0];
  assign MultLoop_mux1h_519_nl = MUX1HOT_v_22_5_2(z_out_213, z_out_773, z_out_220,
      z_out_224, z_out_764, {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[2])});
  assign MultLoop_mux1h_520_nl = MUX1HOT_v_22_5_2(z_out_214, z_out_769, z_out_448,
      z_out_225, z_out_754, {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[2])});
  assign nl_z_out_770 = (MultLoop_mux1h_519_nl) + (MultLoop_mux1h_520_nl);
  assign z_out_770 = nl_z_out_770[21:0];
  assign MultLoop_mux1h_521_nl = MUX1HOT_v_22_5_2(z_out_216, z_out_497, z_out_292,
      z_out_495, z_out_222, {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[2]) , AccumDotWidth_or_38_cse});
  assign nl_MultLoop_acc_1637_nl = z_out_505 + z_out_485;
  assign MultLoop_acc_1637_nl = nl_MultLoop_acc_1637_nl[21:0];
  assign MultLoop_mux1h_522_nl = MUX1HOT_v_22_5_2(z_out_217, z_out_465, z_out_289,
      z_out_468, (MultLoop_acc_1637_nl), {MultLoop_or_81_cse , (fsm_output[3]) ,
      (fsm_output[6]) , (fsm_output[2]) , (fsm_output[4])});
  assign nl_z_out_771 = (MultLoop_mux1h_521_nl) + (MultLoop_mux1h_522_nl);
  assign z_out_771 = nl_z_out_771[21:0];
  assign AccumDotWidth_mux1h_1398_nl = MUX1HOT_v_22_5_2(z_out_751, z_out_226, z_out_495,
      MultLoop_acc_308_itm, z_out_230, {(fsm_output[2]) , MultLoop_or_81_cse , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[4])});
  assign AccumDotWidth_mux1h_1399_nl = MUX1HOT_v_22_6_2(z_out_752, z_out_222, z_out_468,
      AccumDotWidth_acc_1274_itm, z_out_216, z_out_232, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_772 = (AccumDotWidth_mux1h_1398_nl) + (AccumDotWidth_mux1h_1399_nl);
  assign z_out_772 = nl_z_out_772[21:0];
  assign MultLoop_mux1h_523_nl = MUX1HOT_v_22_5_2(z_out_133_28_7, z_out_126_28_7,
      z_out_91_28_7, z_out_759, z_out_144_28_7, {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign MultLoop_mux1h_524_nl = MUX1HOT_v_22_5_2(z_out_134_28_7, z_out_136_28_7,
      z_out_86_28_7, z_out_760, z_out_140_28_7, {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_z_out_773 = (MultLoop_mux1h_523_nl) + (MultLoop_mux1h_524_nl);
  assign z_out_773 = nl_z_out_773[21:0];
  assign MultLoop_mux1h_525_nl = MUX1HOT_v_22_5_2(z_out_224, z_out_464, z_out_290,
      z_out_440, z_out_216, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[3]) , (fsm_output[4])});
  assign MultLoop_mux1h_526_nl = MUX1HOT_v_22_4_2(z_out_219, z_out_271, z_out_302,
      z_out_439, {AccumDotWidth_or_132_cse_1 , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[3])});
  assign nl_z_out_774 = (MultLoop_mux1h_525_nl) + (MultLoop_mux1h_526_nl);
  assign z_out_774 = nl_z_out_774[21:0];
  assign AccumDotWidth_mux1h_1400_nl = MUX1HOT_v_22_4_2(z_out_525, z_out_288, z_out_298,
      z_out_438, {(fsm_output[2]) , (fsm_output[4]) , MultLoop_or_81_cse , (fsm_output[3])});
  assign AccumDotWidth_mux1h_1401_nl = MUX1HOT_v_22_5_2(z_out_530, z_out_212, z_out_288,
      z_out_303, z_out_437, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[3])});
  assign nl_z_out_775 = (AccumDotWidth_mux1h_1400_nl) + (AccumDotWidth_mux1h_1401_nl);
  assign z_out_775 = nl_z_out_775[21:0];
  assign MultLoop_mux1h_527_nl = MUX1HOT_v_22_5_2(z_out_303, z_out_294, z_out_442,
      z_out_439, MultLoop_acc_499_itm, {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[2]) , AccumDotWidth_or_145_cse});
  assign MultLoop_mux1h_528_nl = MUX1HOT_v_22_6_2(z_out_225, z_out_290, z_out_449,
      z_out_438, MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_298, {(fsm_output[5]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[2])
      , (fsm_output[6]) , (fsm_output[4])});
  assign nl_z_out_776 = (MultLoop_mux1h_527_nl) + (MultLoop_mux1h_528_nl);
  assign z_out_776 = nl_z_out_776[21:0];
  assign MultLoop_mux1h_529_nl = MUX1HOT_v_22_6_2(z_out_298, z_out_465, z_out_452,
      z_out_221, z_out_442, z_out_840, {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_530_nl = MUX1HOT_v_22_5_2(z_out_303, z_out_496, z_out_457,
      z_out_233, z_out_441, {(fsm_output[6]) , (fsm_output[1]) , MultLoop_or_93_cse
      , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out_777 = (MultLoop_mux1h_529_nl) + (MultLoop_mux1h_530_nl);
  assign z_out_777 = nl_z_out_777[21:0];
  assign AccumDotWidth_mux1h_1402_nl = MUX1HOT_v_22_6_2(z_out_704, z_out_388, z_out_358,
      z_out_347, z_out_717, (z_out_1086_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1403_nl = MUX1HOT_v_22_6_2(z_out_707, z_out_380, z_out_353,
      z_out_350, z_out_714, (z_out_1089_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_778 = (AccumDotWidth_mux1h_1402_nl) + (AccumDotWidth_mux1h_1403_nl);
  assign z_out_778 = nl_z_out_778[21:0];
  assign MultLoop_or_113_nl = (fsm_output[4]) | or_tmp_4503;
  assign MultLoop_mux1h_531_nl = MUX1HOT_v_22_4_2(MultLoop_acc_1007_itm, z_out_298,
      z_out_214, z_out_290, {(MultLoop_or_113_nl) , (fsm_output[3]) , (fsm_output[1])
      , (fsm_output[7])});
  assign MultLoop_mux1h_532_nl = MUX1HOT_v_22_5_2(z_out_447, z_out_290, z_out_292,
      z_out_214, MultLoop_acc_1000_itm, {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[1])
      , (fsm_output[7]) , or_tmp_4503});
  assign nl_z_out_779 = (MultLoop_mux1h_531_nl) + (MultLoop_mux1h_532_nl);
  assign z_out_779 = nl_z_out_779[21:0];
  assign AccumDotWidth_mux_149_nl = MUX_v_22_2_2(AccumDotWidth_acc_1181_itm, (z_out_867_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_150_nl = MUX_v_22_2_2(z_out_428, (z_out_866_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_780 = (AccumDotWidth_mux_149_nl) + (AccumDotWidth_mux_150_nl);
  assign z_out_780 = nl_z_out_780[21:0];
  assign MultLoop_mux1h_533_nl = MUX1HOT_v_22_5_2(z_out_299, z_out_458, z_out_292,
      z_out_225, z_out_39_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[3])});
  assign MultLoop_mux1h_534_nl = MUX1HOT_v_22_5_2(z_out_297, z_out_450, z_out_294,
      z_out_296, z_out_38_28_7, {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])
      , (fsm_output[1]) , (fsm_output[3])});
  assign nl_z_out_781 = (MultLoop_mux1h_533_nl) + (MultLoop_mux1h_534_nl);
  assign z_out_781 = nl_z_out_781[21:0];
  assign MultLoop_mux1h_535_nl = MUX1HOT_v_22_4_2(z_out_230, z_out_453, z_out_293,
      z_out_755, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[2])});
  assign nl_MultLoop_acc_1638_nl = z_out_834 + z_out_438;
  assign MultLoop_acc_1638_nl = nl_MultLoop_acc_1638_nl[21:0];
  assign MultLoop_mux1h_536_nl = MUX1HOT_v_22_4_2(z_out_212, (MultLoop_acc_1638_nl),
      z_out_296, z_out_758, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2])});
  assign nl_z_out_782 = (MultLoop_mux1h_535_nl) + (MultLoop_mux1h_536_nl);
  assign z_out_782 = nl_z_out_782[21:0];
  assign MultLoop_or_114_nl = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[2]);
  assign MultLoop_mux1h_537_nl = MUX1HOT_v_22_5_2(z_out_438, MultLoop_acc_102_itm,
      z_out_764, z_out_786, z_out_294, {(fsm_output[7]) , (MultLoop_or_114_nl) ,
      (fsm_output[5]) , (fsm_output[1]) , (fsm_output[3])});
  assign MultLoop_mux1h_538_nl = MUX1HOT_v_22_6_2(z_out_499, z_out_303, z_out_752,
      z_out_232, MultLoop_acc_1089_itm, MultLoop_acc_1010_itm, {(fsm_output[7]) ,
      MultLoop_or_46_cse , (fsm_output[5]) , (fsm_output[1]) , (fsm_output[6]) ,
      (fsm_output[2])});
  assign nl_z_out_783 = (MultLoop_mux1h_537_nl) + (MultLoop_mux1h_538_nl);
  assign z_out_783 = nl_z_out_783[21:0];
  assign MultLoop_mux1h_539_nl = MUX1HOT_v_22_4_2(z_out_477, MultLoop_acc_243_itm,
      z_out_763, z_out_773, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[2])
      , (fsm_output[5])});
  assign MultLoop_mux1h_540_nl = MUX1HOT_v_22_4_2(z_out_482, z_out_443, z_out_756,
      z_out_769, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[5])});
  assign nl_z_out_784 = (MultLoop_mux1h_539_nl) + (MultLoop_mux1h_540_nl);
  assign z_out_784 = nl_z_out_784[21:0];
  assign MultLoop_mux1h_541_nl = MUX1HOT_v_22_3_2(z_out_291, z_out_302, z_out_304,
      {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])});
  assign MultLoop_MultLoop_mux_15_nl = MUX_v_22_2_2(z_out_295, z_out_226, fsm_output[4]);
  assign nl_z_out_785 = (MultLoop_mux1h_541_nl) + (MultLoop_MultLoop_mux_15_nl);
  assign z_out_785 = nl_z_out_785[21:0];
  assign nl_MultLoop_acc_1639_nl = z_out_655_28_7 + z_out_656_28_7;
  assign MultLoop_acc_1639_nl = nl_MultLoop_acc_1639_nl[21:0];
  assign nl_MultLoop_acc_1640_nl = z_out_84_28_7 + z_out_89_28_7;
  assign MultLoop_acc_1640_nl = nl_MultLoop_acc_1640_nl[21:0];
  assign MultLoop_mux1h_542_nl = MUX1HOT_v_22_5_2((MultLoop_acc_1639_nl), z_out_505,
      z_out_452, MultLoop_acc_626_itm, (MultLoop_acc_1640_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_145_cse , (fsm_output[5])});
  assign nl_MultLoop_acc_1641_nl = z_out_78_28_7 + z_out_68_28_7;
  assign MultLoop_acc_1641_nl = nl_MultLoop_acc_1641_nl[21:0];
  assign MultLoop_mux1h_543_nl = MUX1HOT_v_22_6_2(z_out_442, z_out_221, z_out_457,
      AccumDotWidth_acc_1167_itm, (MultLoop_acc_1641_nl), z_out_436, {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_786 = (MultLoop_mux1h_542_nl) + (MultLoop_mux1h_543_nl);
  assign z_out_786 = nl_z_out_786[21:0];
  assign MultLoop_mux1h_544_nl = MUX1HOT_v_22_3_2(z_out_296, z_out_297, z_out_215,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign MultLoop_mux1h_545_nl = MUX1HOT_v_22_3_2(z_out_213, z_out_293, z_out_212,
      {(fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])});
  assign nl_z_out_787 = (MultLoop_mux1h_544_nl) + (MultLoop_mux1h_545_nl);
  assign z_out_787 = nl_z_out_787[21:0];
  assign MultLoop_mux1h_546_nl = MUX1HOT_v_22_6_2(z_out_213, z_out_304, z_out_277,
      MultLoop_acc_372_itm, z_out_289, z_out_786, {(fsm_output[7]) , (fsm_output[1])
      , (fsm_output[2]) , AccumDotWidth_or_145_cse , (fsm_output[3]) , (fsm_output[5])});
  assign MultLoop_mux1h_547_nl = MUX1HOT_v_22_7_2(z_out_292, z_out_218, z_out_284,
      MultLoop_acc_113_itm, z_out_295, z_out_777, z_out_446, {(fsm_output[7]) , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_788 = (MultLoop_mux1h_546_nl) + (MultLoop_mux1h_547_nl);
  assign z_out_788 = nl_z_out_788[21:0];
  assign MultLoop_mux1h_548_nl = MUX1HOT_v_22_3_2(z_out_297, z_out_293, z_out_302,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])});
  assign MultLoop_mux1h_549_nl = MUX1HOT_v_22_3_2(z_out_291, z_out_215, z_out_299,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1])});
  assign nl_z_out_789 = (MultLoop_mux1h_548_nl) + (MultLoop_mux1h_549_nl);
  assign z_out_789 = nl_z_out_789[21:0];
  assign MultLoop_mux1h_550_nl = MUX1HOT_v_22_3_2(z_out_213, z_out_289, MultLoop_acc_483_itm,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign MultLoop_mux1h_551_nl = MUX1HOT_v_22_3_2(z_out_215, z_out_299, z_out_290,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[4])});
  assign nl_z_out_790 = (MultLoop_mux1h_550_nl) + (MultLoop_mux1h_551_nl);
  assign z_out_790 = nl_z_out_790[21:0];
  assign AccumDotWidth_mux_151_nl = MUX_v_22_2_2(AccumDotWidth_acc_1326_itm, (z_out_1187_29_7[21:0]),
      fsm_output[8]);
  assign AccumDotWidth_mux_152_nl = MUX_v_22_2_2(z_out_426, (z_out_892_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_791 = (AccumDotWidth_mux_151_nl) + (AccumDotWidth_mux_152_nl);
  assign z_out_791 = nl_z_out_791[21:0];
  assign MultLoop_mux_101_nl = MUX_v_22_2_2(MultLoop_acc_356_itm, z_out_73_28_7,
      fsm_output[3]);
  assign MultLoop_mux_102_nl = MUX_v_22_2_2(z_out_292, z_out_72_28_7, fsm_output[3]);
  assign nl_z_out_792 = (MultLoop_mux_101_nl) + (MultLoop_mux_102_nl);
  assign z_out_792 = nl_z_out_792[21:0];
  assign AccumDotWidth_mux1h_1404_nl = MUX1HOT_v_22_3_2(z_out_708, z_out_697, (z_out_1083_29_7[21:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1405_nl = MUX1HOT_v_22_3_2(z_out_703, z_out_692, (z_out_1082_29_7[21:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_793 = (AccumDotWidth_mux1h_1404_nl) + (AccumDotWidth_mux1h_1405_nl);
  assign z_out_793 = nl_z_out_793[21:0];
  assign MultLoop_mux1h_552_nl = MUX1HOT_v_22_7_2(AccumDotWidth_acc_1378_itm, z_out_422,
      z_out_360, z_out_424, z_out_414, AccumDotWidth_acc_1871_itm, (z_out_1009_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign MultLoop_mux1h_553_nl = MUX1HOT_v_22_7_2(MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_423, z_out_361, z_out_431, z_out_417, z_out_740, (z_out_922_29_7[21:0]),
      {(fsm_output[6]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_794 = (MultLoop_mux1h_552_nl) + (MultLoop_mux1h_553_nl);
  assign z_out_794 = nl_z_out_794[21:0];
  assign AccumDotWidth_mux1h_1406_nl = MUX1HOT_v_22_7_2(z_out_461, z_out_395, z_out_385,
      z_out_372, z_out_402, z_out_739, (z_out_930_29_7[21:0]), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1407_nl = MUX1HOT_v_22_6_2(z_out_462, z_out_399, z_out_382,
      z_out_699, z_out_385, (z_out_924_29_7[21:0]), {(fsm_output[2]) , (fsm_output[1])
      , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_795 = (AccumDotWidth_mux1h_1406_nl) + (AccumDotWidth_mux1h_1407_nl);
  assign z_out_795 = nl_z_out_795[21:0];
  assign MultLoop_mux1h_554_nl = MUX1HOT_v_22_6_2(z_out_292, z_out_284, z_out_777,
      MultLoop_acc_229_itm, z_out_289, z_out_218, {(fsm_output[3]) , (fsm_output[6])
      , (fsm_output[1]) , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[7])
      , (fsm_output[5])});
  assign MultLoop_mux1h_555_nl = MUX1HOT_v_22_7_2(z_out_288, z_out_276, z_out_784,
      z_out_289, MultLoop_acc_1089_itm, MultLoop_acc_968_itm, z_out_232, {(fsm_output[3])
      , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[2]) , (fsm_output[7])
      , (fsm_output[5])});
  assign nl_z_out_796 = (MultLoop_mux1h_554_nl) + (MultLoop_mux1h_555_nl);
  assign z_out_796 = nl_z_out_796[21:0];
  assign nl_AccumDotWidth_acc_2689_nl = conv_s2s_21_22(z_out_597_29_7[22:2]) + conv_s2s_21_22(z_out_1052_29_7[22:2]);
  assign AccumDotWidth_acc_2689_nl = nl_AccumDotWidth_acc_2689_nl[21:0];
  assign nl_AccumDotWidth_acc_2690_nl = conv_s2s_21_22(z_out_1073_29_7[22:2]) + conv_s2s_21_22(z_out_929_29_7[22:2]);
  assign AccumDotWidth_acc_2690_nl = nl_AccumDotWidth_acc_2690_nl[21:0];
  assign AccumDotWidth_mux1h_1408_nl = MUX1HOT_v_22_4_2((AccumDotWidth_acc_2689_nl),
      (AccumDotWidth_acc_2690_nl), z_out_745, (z_out_1093_29_7[21:0]), {(fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2691_nl = conv_s2s_21_22(z_out_1151_29_7[22:2]) + conv_s2s_21_22(z_out_1103_29_7[22:2]);
  assign AccumDotWidth_acc_2691_nl = nl_AccumDotWidth_acc_2691_nl[21:0];
  assign nl_AccumDotWidth_acc_2692_nl = conv_s2s_21_22(z_out_1133_29_9) + conv_s2s_21_22(z_out_1013_29_7[22:2]);
  assign AccumDotWidth_acc_2692_nl = nl_AccumDotWidth_acc_2692_nl[21:0];
  assign AccumDotWidth_mux1h_1409_nl = MUX1HOT_v_22_4_2((AccumDotWidth_acc_2691_nl),
      (AccumDotWidth_acc_2692_nl), z_out_744, (z_out_1090_29_7[21:0]), {(fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_797 = (AccumDotWidth_mux1h_1408_nl) + (AccumDotWidth_mux1h_1409_nl);
  assign z_out_797 = nl_z_out_797[21:0];
  assign MultLoop_mux_103_nl = MUX_v_22_2_2(z_out_291, z_out_124_28_7, fsm_output[3]);
  assign MultLoop_mux_104_nl = MUX_v_22_2_2(z_out_217, z_out_129_28_7, fsm_output[3]);
  assign nl_z_out_798 = (MultLoop_mux_103_nl) + (MultLoop_mux_104_nl);
  assign z_out_798 = nl_z_out_798[21:0];
  assign nl_AccumDotWidth_acc_2693_nl = conv_s2s_21_22(z_out_1167_29_7[22:2]) + conv_s2s_21_22(z_out_862_29_7[22:2]);
  assign AccumDotWidth_acc_2693_nl = nl_AccumDotWidth_acc_2693_nl[21:0];
  assign nl_AccumDotWidth_acc_2694_nl = conv_s2s_21_22(z_out_876_29_7[22:2]) + conv_s2s_21_22(z_out_884_29_7[22:2]);
  assign AccumDotWidth_acc_2694_nl = nl_AccumDotWidth_acc_2694_nl[21:0];
  assign AccumDotWidth_mux1h_1410_nl = MUX1HOT_v_22_6_2(z_out_746, z_out_714, (AccumDotWidth_acc_2693_nl),
      (AccumDotWidth_acc_2694_nl), z_out_748, (z_out_1172_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2695_nl = conv_s2s_21_22(z_out_930_29_7[22:2]) + conv_s2s_21_22(z_out_903_29_7[22:2]);
  assign AccumDotWidth_acc_2695_nl = nl_AccumDotWidth_acc_2695_nl[21:0];
  assign nl_AccumDotWidth_acc_2696_nl = conv_s2s_21_22(z_out_1029_29_7[22:2]) + conv_s2s_21_22(z_out_618_29_7[22:2]);
  assign AccumDotWidth_acc_2696_nl = nl_AccumDotWidth_acc_2696_nl[21:0];
  assign AccumDotWidth_mux1h_1411_nl = MUX1HOT_v_22_6_2(z_out_747, z_out_715, (AccumDotWidth_acc_2695_nl),
      (AccumDotWidth_acc_2696_nl), z_out_746, (z_out_1156_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_799 = (AccumDotWidth_mux1h_1410_nl) + (AccumDotWidth_mux1h_1411_nl);
  assign z_out_799 = nl_z_out_799[21:0];
  assign MultLoop_mux_105_nl = MUX_v_22_2_2(z_out_304, z_out_75_28_7, fsm_output[3]);
  assign MultLoop_mux_106_nl = MUX_v_22_2_2(z_out_214, z_out_69_28_7, fsm_output[3]);
  assign nl_z_out_800 = (MultLoop_mux_105_nl) + (MultLoop_mux_106_nl);
  assign z_out_800 = nl_z_out_800[21:0];
  assign nl_AccumDotWidth_acc_2697_nl = conv_s2s_21_22(z_out_1104_29_7[22:2]) + conv_s2s_21_22(z_out_967_29_7[22:2]);
  assign AccumDotWidth_acc_2697_nl = nl_AccumDotWidth_acc_2697_nl[21:0];
  assign AccumDotWidth_mux_153_nl = MUX_v_22_2_2((AccumDotWidth_acc_2697_nl), (z_out_1170_29_7[21:0]),
      fsm_output[8]);
  assign nl_AccumDotWidth_acc_2698_nl = conv_s2s_21_22(z_out_1131_29_7[22:2]) + conv_s2s_21_22(z_out_1021_29_7[22:2]);
  assign AccumDotWidth_acc_2698_nl = nl_AccumDotWidth_acc_2698_nl[21:0];
  assign AccumDotWidth_mux_154_nl = MUX_v_22_2_2((AccumDotWidth_acc_2698_nl), (z_out_1158_29_7[21:0]),
      fsm_output[8]);
  assign nl_z_out_801 = (AccumDotWidth_mux_153_nl) + (AccumDotWidth_mux_154_nl);
  assign z_out_801 = nl_z_out_801[21:0];
  assign nl_AccumDotWidth_acc_2699_nl = conv_s2s_21_22(z_out_868_29_7[22:2]) + conv_s2s_21_22(z_out_931_29_7[22:2]);
  assign AccumDotWidth_acc_2699_nl = nl_AccumDotWidth_acc_2699_nl[21:0];
  assign nl_AccumDotWidth_acc_2700_nl = conv_s2s_21_22(z_out_1164_29_7[22:2]) + conv_s2s_21_22(z_out_875_29_7[22:2]);
  assign AccumDotWidth_acc_2700_nl = nl_AccumDotWidth_acc_2700_nl[21:0];
  assign nl_AccumDotWidth_acc_2701_nl = conv_s2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm)
      + conv_s2s_21_22(z_out_990_29_7[22:2]);
  assign AccumDotWidth_acc_2701_nl = nl_AccumDotWidth_acc_2701_nl[21:0];
  assign AccumDotWidth_mux1h_1412_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2699_nl),
      z_out_354, (AccumDotWidth_acc_2700_nl), z_out_395, (AccumDotWidth_acc_2701_nl),
      z_out_747, (z_out_1011_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2702_nl = conv_s2s_21_22(z_out_924_29_7[22:2]) + conv_s2s_21_22(z_out_926_29_7[22:2]);
  assign AccumDotWidth_acc_2702_nl = nl_AccumDotWidth_acc_2702_nl[21:0];
  assign nl_AccumDotWidth_acc_2703_nl = conv_s2s_21_22(z_out_923_29_7[22:2]) + conv_s2s_21_22(z_out_967_29_7[22:2]);
  assign AccumDotWidth_acc_2703_nl = nl_AccumDotWidth_acc_2703_nl[21:0];
  assign nl_AccumDotWidth_acc_2704_nl = conv_s2s_21_22(z_out_1075_29_7[22:2]) + conv_s2s_21_22(z_out_1067_29_9);
  assign AccumDotWidth_acc_2704_nl = nl_AccumDotWidth_acc_2704_nl[21:0];
  assign AccumDotWidth_mux1h_1413_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2702_nl),
      z_out_357, (AccumDotWidth_acc_2703_nl), z_out_386, (AccumDotWidth_acc_2704_nl),
      z_out_741, (z_out_1013_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_802 = (AccumDotWidth_mux1h_1412_nl) + (AccumDotWidth_mux1h_1413_nl);
  assign z_out_802 = nl_z_out_802[21:0];
  assign MultLoop_mux_107_nl = MUX_v_22_2_2(z_out_294, z_out_135_28_7, fsm_output[3]);
  assign MultLoop_mux_108_nl = MUX_v_22_2_2(z_out_295, z_out_130_28_7, fsm_output[3]);
  assign nl_z_out_803 = (MultLoop_mux_107_nl) + (MultLoop_mux_108_nl);
  assign z_out_803 = nl_z_out_803[21:0];
  assign nl_AccumDotWidth_acc_2705_nl = conv_s2s_21_22(z_out_870_29_7[22:2]) + conv_s2s_21_22(z_out_869_29_7[22:2]);
  assign AccumDotWidth_acc_2705_nl = nl_AccumDotWidth_acc_2705_nl[21:0];
  assign AccumDotWidth_mux1h_1414_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2705_nl),
      z_out_716, z_out_356, z_out_732, z_out_372, (z_out_929_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2706_nl = conv_s2s_21_22(z_out_874_29_7[22:2]) + conv_s2s_21_22(z_out_878_29_7[22:2]);
  assign AccumDotWidth_acc_2706_nl = nl_AccumDotWidth_acc_2706_nl[21:0];
  assign AccumDotWidth_mux1h_1415_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2706_nl),
      z_out_717, z_out_361, z_out_737, z_out_371, (z_out_893_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_804 = (AccumDotWidth_mux1h_1414_nl) + (AccumDotWidth_mux1h_1415_nl);
  assign z_out_804 = nl_z_out_804[21:0];
  assign nl_AccumDotWidth_acc_2707_nl = conv_s2s_21_22(z_out_866_29_7[22:2]) + conv_s2s_21_22(z_out_873_29_7[22:2]);
  assign AccumDotWidth_acc_2707_nl = nl_AccumDotWidth_acc_2707_nl[21:0];
  assign nl_AccumDotWidth_acc_2708_nl = conv_s2s_21_22(z_out_953_29_7[22:2]) + conv_s2s_21_22(z_out_1168_29_7[22:2]);
  assign AccumDotWidth_acc_2708_nl = nl_AccumDotWidth_acc_2708_nl[21:0];
  assign nl_AccumDotWidth_acc_2709_nl = conv_s2s_21_22(z_out_1029_29_7[22:2]) + conv_s2s_21_22(z_out_1015_29_7[22:2]);
  assign AccumDotWidth_acc_2709_nl = nl_AccumDotWidth_acc_2709_nl[21:0];
  assign AccumDotWidth_mux1h_1416_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2707_nl),
      z_out_362, z_out_360, (AccumDotWidth_acc_2708_nl), (AccumDotWidth_acc_2709_nl),
      z_out_382, (z_out_1157_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2710_nl = conv_s2s_21_22(z_out_867_29_7[22:2]) + conv_s2s_21_22(z_out_871_29_7[22:2]);
  assign AccumDotWidth_acc_2710_nl = nl_AccumDotWidth_acc_2710_nl[21:0];
  assign nl_AccumDotWidth_acc_2711_nl = conv_s2s_21_22(z_out_919_29_7[22:2]) + conv_s2s_21_22(z_out_1085_29_7[22:2]);
  assign AccumDotWidth_acc_2711_nl = nl_AccumDotWidth_acc_2711_nl[21:0];
  assign nl_AccumDotWidth_acc_2712_nl = conv_s2s_21_22(z_out_1039_29_7[22:2]) + conv_s2s_21_22(z_out_962_29_9);
  assign AccumDotWidth_acc_2712_nl = nl_AccumDotWidth_acc_2712_nl[21:0];
  assign AccumDotWidth_mux1h_1417_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2710_nl),
      z_out_352, z_out_359, (AccumDotWidth_acc_2711_nl), (AccumDotWidth_acc_2712_nl),
      z_out_374, (z_out_1185_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_805 = (AccumDotWidth_mux1h_1416_nl) + (AccumDotWidth_mux1h_1417_nl);
  assign z_out_805 = nl_z_out_805[21:0];
  assign nl_MultLoop_acc_1642_nl = (MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[21:11])
      + conv_s2s_8_11(InitAccum_io_read_b4_rsc_cse_sva[79:72]);
  assign MultLoop_acc_1642_nl = nl_MultLoop_acc_1642_nl[10:0];
  assign AccumDotWidth_mux1h_1418_nl = MUX1HOT_v_22_7_2(z_out_710, z_out_718, z_out_379,
      z_out_700, z_out_380, z_out_377, ({(MultLoop_acc_1642_nl) , (MultLoop_1123_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[10:0])}),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1419_nl = MUX1HOT_v_22_7_2(z_out_398, z_out_719, z_out_377,
      z_out_705, z_out_385, AccumDotWidth_acc_1837_itm, AccumDotWidth_acc_1133_itm,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_806 = (AccumDotWidth_mux1h_1418_nl) + (AccumDotWidth_mux1h_1419_nl);
  assign z_out_806 = nl_z_out_806[21:0];
  assign nl_AccumDotWidth_acc_2713_nl = conv_s2s_21_22(z_out_933_29_7[22:2]) + conv_s2s_21_22(z_out_936_29_7[22:2]);
  assign AccumDotWidth_acc_2713_nl = nl_AccumDotWidth_acc_2713_nl[21:0];
  assign nl_AccumDotWidth_acc_2714_nl = conv_s2s_21_22(z_out_1106_29_7[22:2]) + conv_s2s_21_22(z_out_1013_29_7[22:2]);
  assign AccumDotWidth_acc_2714_nl = nl_AccumDotWidth_acc_2714_nl[21:0];
  assign nl_AccumDotWidth_acc_2715_nl = conv_s2s_21_22(z_out_961_29_7[22:2]) + conv_s2s_21_22(z_out_1068_29_7[22:2]);
  assign AccumDotWidth_acc_2715_nl = nl_AccumDotWidth_acc_2715_nl[21:0];
  assign AccumDotWidth_mux1h_1420_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2713_nl),
      z_out_358, (AccumDotWidth_acc_2714_nl), z_out_392, (AccumDotWidth_acc_2715_nl),
      z_out_742, (z_out_864_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_AccumDotWidth_acc_2716_nl = conv_s2s_21_22(z_out_935_29_7[22:2]) + conv_s2s_21_22(z_out_927_29_7[22:2]);
  assign AccumDotWidth_acc_2716_nl = nl_AccumDotWidth_acc_2716_nl[21:0];
  assign nl_AccumDotWidth_acc_2717_nl = conv_s2s_21_22(z_out_870_29_7[22:2]) + conv_s2s_21_22(z_out_1033_29_9);
  assign AccumDotWidth_acc_2717_nl = nl_AccumDotWidth_acc_2717_nl[21:0];
  assign nl_AccumDotWidth_acc_2718_nl = conv_s2s_21_22(z_out_605_29_7[22:2]) + conv_s2s_21_22(z_out_882_29_7[22:2]);
  assign AccumDotWidth_acc_2718_nl = nl_AccumDotWidth_acc_2718_nl[21:0];
  assign AccumDotWidth_mux1h_1421_nl = MUX1HOT_v_22_7_2((AccumDotWidth_acc_2716_nl),
      z_out_356, (AccumDotWidth_acc_2717_nl), z_out_389, (AccumDotWidth_acc_2718_nl),
      z_out_743, (z_out_863_29_7[21:0]), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_807 = (AccumDotWidth_mux1h_1420_nl) + (AccumDotWidth_mux1h_1421_nl);
  assign z_out_807 = nl_z_out_807[21:0];
  assign AccumDotWidth_mux1h_1422_nl = MUX1HOT_v_22_6_2(z_out_381, z_out_694, z_out_733,
      z_out_318, z_out_450, z_out_754, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1423_nl = MUX1HOT_v_22_6_2(z_out_383, z_out_697, z_out_739,
      z_out_508, z_out_244, z_out_469, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_808 = (AccumDotWidth_mux1h_1422_nl) + (AccumDotWidth_mux1h_1423_nl);
  assign z_out_808 = nl_z_out_808[21:0];
  assign AccumDotWidth_mux1h_1424_nl = MUX1HOT_v_22_8_2(z_out_732, AccumDotWidth_acc_1274_itm,
      z_out_467, z_out_816, z_out_319, z_out_454, z_out_541, AccumDotWidth_acc_1378_itm,
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1425_nl = MUX1HOT_v_22_8_2(z_out_735, MultLoop_acc_113_itm,
      z_out_842, z_out_536, z_out_509, z_out_549, z_out_317, z_out_285, {(fsm_output[1])
      , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_809 = (AccumDotWidth_mux1h_1424_nl) + (AccumDotWidth_mux1h_1425_nl);
  assign z_out_809 = nl_z_out_809[21:0];
  assign nl_MultLoop_acc_1643_nl = z_out_227 + z_out_529;
  assign MultLoop_acc_1643_nl = nl_MultLoop_acc_1643_nl[21:0];
  assign MultLoop_mux_109_nl = MUX_v_22_2_2(z_out_151_28_7, (MultLoop_acc_1643_nl),
      fsm_output[8]);
  assign MultLoop_mux_110_nl = MUX_v_22_2_2(z_out_152_28_7, z_out_470, fsm_output[8]);
  assign nl_z_out_810 = (MultLoop_mux_109_nl) + (MultLoop_mux_110_nl);
  assign z_out_810 = nl_z_out_810[21:0];
  assign nl_MultLoop_acc_1645_nl = MultLoop_acc_215_itm + z_out_328;
  assign MultLoop_acc_1645_nl = nl_MultLoop_acc_1645_nl[21:0];
  assign nl_MultLoop_acc_1644_nl = z_out_275 + (MultLoop_acc_1645_nl);
  assign MultLoop_acc_1644_nl = nl_MultLoop_acc_1644_nl[21:0];
  assign AccumDotWidth_mux1h_1426_nl = MUX1HOT_v_22_8_2(z_out_738, z_out_676_28_7,
      z_out_689, z_out_467, z_out_317, z_out_264, z_out_265, (MultLoop_acc_1644_nl),
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1427_nl = MUX1HOT_v_22_8_2(z_out_734, z_out_667_28_7,
      z_out_691, z_out_456, z_out_510, z_out_326, z_out_836, z_out_481, {(fsm_output[1])
      , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_811 = (AccumDotWidth_mux1h_1426_nl) + (AccumDotWidth_mux1h_1427_nl);
  assign z_out_811 = nl_z_out_811[21:0];
  assign AccumDotWidth_mux1h_1428_nl = MUX1HOT_v_22_8_2(z_out_725, z_out_844, z_out_267,
      z_out_466, z_out_816, z_out_471, z_out_835, z_out_758, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1429_nl = MUX1HOT_v_22_7_2(z_out_731, z_out_319, z_out_557,
      z_out_472, AccumDotWidth_acc_1186_itm, z_out_270, AccumDotWidth_acc_1181_itm,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , AccumDotWidth_or_145_cse
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_812 = (AccumDotWidth_mux1h_1428_nl) + (AccumDotWidth_mux1h_1429_nl);
  assign z_out_812 = nl_z_out_812[21:0];
  assign AccumDotWidth_mux1h_1430_nl = MUX1HOT_v_22_7_2(z_out_733, z_out_826, z_out_263,
      z_out_467, z_out_481, z_out_269, z_out_530, {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1431_nl = MUX1HOT_v_22_7_2(z_out_737, z_out_547, z_out_844,
      z_out_269, z_out_473, z_out_837, AccumDotWidth_acc_1186_itm, {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_813 = (AccumDotWidth_mux1h_1430_nl) + (AccumDotWidth_mux1h_1431_nl);
  assign z_out_813 = nl_z_out_813[21:0];
  assign MultLoop_mux_111_nl = MUX_v_22_2_2(z_out_668_28_7, MultLoop_acc_372_itm,
      fsm_output[8]);
  assign nl_MultLoop_acc_1646_nl = MultLoop_acc_54_itm + z_out_228;
  assign MultLoop_acc_1646_nl = nl_MultLoop_acc_1646_nl[21:0];
  assign MultLoop_mux_112_nl = MUX_v_22_2_2(z_out_669_28_7, (MultLoop_acc_1646_nl),
      fsm_output[8]);
  assign nl_z_out_814 = (MultLoop_mux_111_nl) + (MultLoop_mux_112_nl);
  assign z_out_814 = nl_z_out_814[21:0];
  assign nl_AccumDotWidth_acc_2719_nl = conv_s2s_21_22(z_out_890_29_7[22:2]) + conv_s2s_21_22(z_out_608_29_7[22:2]);
  assign AccumDotWidth_acc_2719_nl = nl_AccumDotWidth_acc_2719_nl[21:0];
  assign nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[9999:9992]));
  assign MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1649_nl = (readslicef_29_22_7((MultLoop_1250_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)))
      + MultLoop_1251_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1649_nl = nl_MultLoop_acc_1649_nl[21:0];
  assign nl_MultLoop_acc_1651_nl = MultLoop_1252_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + z_out_669_28_7;
  assign MultLoop_acc_1651_nl = nl_MultLoop_acc_1651_nl[21:0];
  assign nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = $signed(conv_u2s_21_22(nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm))
      * $signed((MultLoop_io_read_w4_rsc_cse_sva[10039:10032]));
  assign MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl
      = nl_MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl[28:0];
  assign nl_MultLoop_acc_1652_nl = z_out_676_28_7 + (readslicef_29_22_7((MultLoop_1255_nnet_product_layer3_t_config4_weight_t_config4_accum_t_mul_1_nl)));
  assign MultLoop_acc_1652_nl = nl_MultLoop_acc_1652_nl[21:0];
  assign nl_MultLoop_acc_1647_nl = z_out_504 + (MultLoop_acc_1649_nl) + (MultLoop_acc_1651_nl)
      + (MultLoop_acc_1652_nl);
  assign MultLoop_acc_1647_nl = nl_MultLoop_acc_1647_nl[21:0];
  assign AccumDotWidth_mux1h_1432_nl = MUX1HOT_v_22_6_2((AccumDotWidth_acc_2719_nl),
      z_out_731, z_out_387, z_out_471, z_out_271, (MultLoop_acc_1647_nl), {(fsm_output[2])
      , (fsm_output[3]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1433_nl = MUX1HOT_v_22_6_2(z_out_379, z_out_735, z_out_394,
      z_out_469, z_out_330, z_out_456, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_815 = (AccumDotWidth_mux1h_1432_nl) + (AccumDotWidth_mux1h_1433_nl);
  assign z_out_815 = nl_z_out_815[21:0];
  assign nl_MultLoop_acc_1654_nl = (z_out_931_29_7[21:0]) + MultLoop_995_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1654_nl = nl_MultLoop_acc_1654_nl[21:0];
  assign nl_MultLoop_acc_1653_nl = z_out_794 + (MultLoop_acc_1654_nl);
  assign MultLoop_acc_1653_nl = nl_MultLoop_acc_1653_nl[21:0];
  assign AccumDotWidth_mux1h_1434_nl = MUX1HOT_v_22_8_2(z_out_432, z_out_484, z_out_736,
      z_out_329, z_out_520, z_out_263, z_out_696, (MultLoop_acc_1653_nl), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1656_nl = (z_out_1012_29_7[21:0]) + (z_out_1014_29_7[21:0]);
  assign MultLoop_acc_1656_nl = nl_MultLoop_acc_1656_nl[21:0];
  assign nl_MultLoop_acc_1655_nl = z_out_257 + (MultLoop_acc_1656_nl);
  assign MultLoop_acc_1655_nl = nl_MultLoop_acc_1655_nl[21:0];
  assign AccumDotWidth_mux1h_1435_nl = MUX1HOT_v_22_8_2(z_out_435, z_out_483, z_out_739,
      z_out_320, AccumDotWidth_acc_1184_itm, AccumDotWidth_acc_1133_itm, z_out_689,
      (MultLoop_acc_1655_nl), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_816 = (AccumDotWidth_mux1h_1434_nl) + (AccumDotWidth_mux1h_1435_nl);
  assign z_out_816 = nl_z_out_816[21:0];
  assign MultLoop_mux_113_nl = MUX_v_22_2_2(z_out_670_28_7, z_out_471, fsm_output[8]);
  assign MultLoop_mux_114_nl = MUX_v_22_2_2(z_out_671_28_7, MultLoop_519_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      fsm_output[8]);
  assign nl_z_out_817 = (MultLoop_mux_113_nl) + (MultLoop_mux_114_nl);
  assign z_out_817 = nl_z_out_817[21:0];
  assign AccumDotWidth_mux1h_1436_nl = MUX1HOT_v_22_5_2(z_out_748, z_out_469, z_out_536,
      z_out_266, z_out_540, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1437_nl = MUX1HOT_v_22_4_2(z_out_742, z_out_450, AccumDotWidth_acc_1169_itm,
      z_out_285, {(fsm_output[2]) , (fsm_output[3]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_48_cse
      , (fsm_output[6])});
  assign nl_z_out_818 = (AccumDotWidth_mux1h_1436_nl) + (AccumDotWidth_mux1h_1437_nl);
  assign z_out_818 = nl_z_out_818[21:0];
  assign MultLoop_mux_115_nl = MUX_v_22_2_2(z_out_459, z_out_539, fsm_output[8]);
  assign MultLoop_mux_116_nl = MUX_v_22_2_2(z_out_453, z_out_847, fsm_output[8]);
  assign nl_z_out_819 = (MultLoop_mux_115_nl) + (MultLoop_mux_116_nl);
  assign z_out_819 = nl_z_out_819[21:0];
  assign MultLoop_mux1h_556_nl = MUX1HOT_v_22_4_2(z_out_169_28_7, z_out_749, z_out_162_28_7,
      z_out_812, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3])});
  assign MultLoop_mux1h_557_nl = MUX1HOT_v_22_4_2(z_out_664_28_7, z_out_743, z_out_149_28_7,
      z_out_542, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[3])});
  assign nl_z_out_820 = (MultLoop_mux1h_556_nl) + (MultLoop_mux1h_557_nl);
  assign z_out_820 = nl_z_out_820[21:0];
  assign MultLoop_mux1h_558_nl = MUX1HOT_v_22_5_2(z_out_165_28_7, z_out_349, z_out_676_28_7,
      z_out_265, z_out_467, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign MultLoop_mux1h_559_nl = MUX1HOT_v_22_5_2(z_out_179_28_7, z_out_356, z_out_665_28_7,
      z_out_275, MultLoop_acc_250_itm, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_821 = (MultLoop_mux1h_558_nl) + (MultLoop_mux1h_559_nl);
  assign z_out_821 = nl_z_out_821[21:0];
  assign AccumDotWidth_mux_155_nl = MUX_v_22_2_2(z_out_463, z_out_534, fsm_output[8]);
  assign nl_z_out_822 = (AccumDotWidth_mux_155_nl) + AccumDotWidth_acc_1184_itm;
  assign z_out_822 = nl_z_out_822[21:0];
  assign nl_MultLoop_acc_1659_nl = z_out_666_28_7 + (z_out_630_29_7[21:0]);
  assign MultLoop_acc_1659_nl = nl_MultLoop_acc_1659_nl[21:0];
  assign nl_MultLoop_acc_1660_nl = z_out_670_28_7 + z_out_671_28_7;
  assign MultLoop_acc_1660_nl = nl_MultLoop_acc_1660_nl[21:0];
  assign nl_MultLoop_acc_1658_nl = (MultLoop_acc_1659_nl) + (MultLoop_acc_1660_nl);
  assign MultLoop_acc_1658_nl = nl_MultLoop_acc_1658_nl[21:0];
  assign nl_MultLoop_acc_1657_nl = z_out_337 + (MultLoop_acc_1658_nl);
  assign MultLoop_acc_1657_nl = nl_MultLoop_acc_1657_nl[21:0];
  assign MultLoop_mux1h_560_nl = MUX1HOT_v_22_5_2(z_out_666_28_7, z_out_746, z_out_150_28_7,
      z_out_453, (MultLoop_acc_1657_nl), {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign MultLoop_mux1h_561_nl = MUX1HOT_v_22_5_2(z_out_149_28_7, z_out_745, z_out_679_28_7,
      z_out_558, z_out_464, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[8])});
  assign nl_z_out_823 = (MultLoop_mux1h_560_nl) + (MultLoop_mux1h_561_nl);
  assign z_out_823 = nl_z_out_823[21:0];
  assign nl_MultLoop_acc_1662_nl = (z_out_943_29_7[21:0]) + (z_out_941_29_7[21:0]);
  assign MultLoop_acc_1662_nl = nl_MultLoop_acc_1662_nl[21:0];
  assign nl_MultLoop_acc_1663_nl = (z_out_940_29_7[21:0]) + (z_out_883_29_7[21:0]);
  assign MultLoop_acc_1663_nl = nl_MultLoop_acc_1663_nl[21:0];
  assign nl_MultLoop_acc_1661_nl = (MultLoop_acc_1662_nl) + (MultLoop_acc_1663_nl);
  assign MultLoop_acc_1661_nl = nl_MultLoop_acc_1661_nl[21:0];
  assign MultLoop_mux1h_562_nl = MUX1HOT_v_22_4_2(z_out_501, z_out_456, z_out_510,
      (MultLoop_acc_1661_nl), {MultLoop_or_89_cse , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[8])});
  assign nl_MultLoop_acc_1665_nl = (z_out_882_29_7[21:0]) + (z_out_888_29_7[21:0]);
  assign MultLoop_acc_1665_nl = nl_MultLoop_acc_1665_nl[21:0];
  assign nl_MultLoop_acc_1666_nl = (z_out_875_29_7[21:0]) + (z_out_886_29_7[21:0]);
  assign MultLoop_acc_1666_nl = nl_MultLoop_acc_1666_nl[21:0];
  assign nl_MultLoop_acc_1664_nl = (MultLoop_acc_1665_nl) + (MultLoop_acc_1666_nl);
  assign MultLoop_acc_1664_nl = nl_MultLoop_acc_1664_nl[21:0];
  assign MultLoop_mux1h_563_nl = MUX1HOT_v_22_4_2(z_out_502, z_out_450, MultLoop_acc_1089_itm,
      (MultLoop_acc_1664_nl), {MultLoop_or_89_cse , (fsm_output[5]) , (fsm_output[3])
      , (fsm_output[8])});
  assign nl_z_out_824 = (MultLoop_mux1h_562_nl) + (MultLoop_mux1h_563_nl);
  assign z_out_824 = nl_z_out_824[21:0];
  assign AccumDotWidth_AccumDotWidth_mux_22_nl = MUX_v_22_2_2(z_out_325, MultLoop_acc_229_itm,
      AccumDotWidth_or_156_cse);
  assign AccumDotWidth_mux1h_1438_nl = MUX1HOT_v_22_4_2(z_out_237, AccumDotWidth_acc_1135_itm,
      z_out_512, z_out_241, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[8])});
  assign nl_z_out_825 = (AccumDotWidth_AccumDotWidth_mux_22_nl) + (AccumDotWidth_mux1h_1438_nl);
  assign z_out_825 = nl_z_out_825[21:0];
  assign MultLoop_mux1h_564_nl = MUX1HOT_v_22_8_2(z_out_171_28_7, z_out_166_28_7,
      z_out_712, z_out_258, z_out_379, z_out_517, z_out_718, z_out_562, {(fsm_output[5])
      , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign MultLoop_mux1h_565_nl = MUX1HOT_v_22_8_2(z_out_665_28_7, z_out_167_28_7,
      z_out_718, z_out_249, z_out_382, z_out_334, z_out_716, MultLoop_acc_994_itm,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_826 = (MultLoop_mux1h_564_nl) + (MultLoop_mux1h_565_nl);
  assign z_out_826 = nl_z_out_826[21:0];
  assign MultLoop_mux_117_nl = MUX_v_22_2_2(z_out_180_28_7, z_out_648_28_7, fsm_output[5]);
  assign MultLoop_mux_118_nl = MUX_v_22_2_2(z_out_178_28_7, z_out_656_28_7, fsm_output[5]);
  assign nl_z_out_827 = (MultLoop_mux_117_nl) + (MultLoop_mux_118_nl);
  assign z_out_827 = nl_z_out_827[21:0];
  assign nl_MultLoop_acc_1667_nl = z_out_806 + MultLoop_acc_1089_itm;
  assign MultLoop_acc_1667_nl = nl_MultLoop_acc_1667_nl[21:0];
  assign MultLoop_mux1h_566_nl = MUX1HOT_v_22_4_2(z_out_150_28_7, z_out_550, z_out_158_28_7,
      (MultLoop_acc_1667_nl), {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[8])});
  assign MultLoop_mux1h_567_nl = MUX1HOT_v_22_4_2(z_out_176_28_7, z_out_548, z_out_159_28_7,
      MultLoop_acc_1121_itm, {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[8])});
  assign nl_z_out_828 = (MultLoop_mux1h_566_nl) + (MultLoop_mux1h_567_nl);
  assign z_out_828 = nl_z_out_828[21:0];
  assign MultLoop_mux1h_568_nl = MUX1HOT_v_22_3_2(z_out_151_28_7, z_out_139_28_7,
      z_out_661_28_7, {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5])});
  assign MultLoop_mux1h_569_nl = MUX1HOT_v_22_3_2(z_out_152_28_7, z_out_193_28_7,
      z_out_632_28_7, {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5])});
  assign nl_z_out_829 = (MultLoop_mux1h_568_nl) + (MultLoop_mux1h_569_nl);
  assign z_out_829 = nl_z_out_829[21:0];
  assign MultLoop_mux1h_570_nl = MUX1HOT_v_22_3_2((z_out_620_29_7[21:0]), z_out_169_28_7,
      z_out_633_28_7, {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5])});
  assign MultLoop_mux1h_571_nl = MUX1HOT_v_22_3_2(z_out_667_28_7, z_out_114_28_7,
      z_out_173_28_7, {(fsm_output[4]) , (fsm_output[6]) , (fsm_output[5])});
  assign nl_z_out_830 = (MultLoop_mux1h_570_nl) + (MultLoop_mux1h_571_nl);
  assign z_out_830 = nl_z_out_830[21:0];
  assign MultLoop_mux1h_572_nl = MUX1HOT_v_22_6_2(z_out_668_28_7, z_out_128_28_7,
      z_out_491, z_out_178_28_7, MultLoop_acc_36_itm, z_out_828, {(fsm_output[4])
      , (fsm_output[5]) , (fsm_output[2]) , (fsm_output[6]) , (fsm_output[3]) , (fsm_output[8])});
  assign MultLoop_mux1h_573_nl = MUX1HOT_v_22_5_2(z_out_669_28_7, z_out_182_28_7,
      MultLoop_391_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      z_out_174_28_7, z_out_248, {(fsm_output[4]) , (fsm_output[5]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_56_cse
      , (fsm_output[6]) , (fsm_output[3])});
  assign nl_z_out_831 = (MultLoop_mux1h_572_nl) + (MultLoop_mux1h_573_nl);
  assign z_out_831 = nl_z_out_831[21:0];
  assign MultLoop_mux1h_574_nl = MUX1HOT_v_22_4_2(z_out_488, z_out_172_28_7, z_out_185_28_7,
      z_out_566, {MultLoop_or_89_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign MultLoop_mux1h_575_nl = MUX1HOT_v_22_5_2(z_out_491, z_out_170_28_7, z_out_164_28_7,
      z_out_504, MultLoop_acc_968_itm, {(fsm_output[6]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[8])});
  assign nl_z_out_832 = (MultLoop_mux1h_574_nl) + (MultLoop_mux1h_575_nl);
  assign z_out_832 = nl_z_out_832[21:0];
  assign nl_MultLoop_acc_1669_nl = (z_out_581_29_7[21:0]) + (z_out_578_29_7[21:0]);
  assign MultLoop_acc_1669_nl = nl_MultLoop_acc_1669_nl[21:0];
  assign nl_MultLoop_acc_1668_nl = z_out_312 + (MultLoop_acc_1669_nl);
  assign MultLoop_acc_1668_nl = nl_MultLoop_acc_1668_nl[21:0];
  assign MultLoop_mux1h_576_nl = MUX1HOT_v_22_5_2(z_out_498, z_out_188_28_7, z_out_494,
      z_out_168_28_7, (MultLoop_acc_1668_nl), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1670_nl = z_out_245 + z_out_308;
  assign MultLoop_acc_1670_nl = nl_MultLoop_acc_1670_nl[21:0];
  assign MultLoop_mux1h_577_nl = MUX1HOT_v_22_5_2(z_out_499, z_out_163_28_7, z_out_498,
      z_out_157_28_7, (MultLoop_acc_1670_nl), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_833 = (MultLoop_mux1h_576_nl) + (MultLoop_mux1h_577_nl);
  assign z_out_833 = nl_z_out_833[21:0];
  assign nl_MultLoop_acc_1672_nl = (z_out_907_29_7[21:0]) + (z_out_918_29_7[21:0]);
  assign MultLoop_acc_1672_nl = nl_MultLoop_acc_1672_nl[21:0];
  assign nl_MultLoop_acc_1673_nl = (z_out_917_29_7[21:0]) + (z_out_987_29_7[21:0]);
  assign MultLoop_acc_1673_nl = nl_MultLoop_acc_1673_nl[21:0];
  assign nl_MultLoop_acc_1671_nl = (MultLoop_acc_1672_nl) + (MultLoop_acc_1673_nl);
  assign MultLoop_acc_1671_nl = nl_MultLoop_acc_1671_nl[21:0];
  assign MultLoop_mux1h_578_nl = MUX1HOT_v_22_5_2(z_out_504, z_out_187_28_7, z_out_499,
      z_out_666_28_7, (MultLoop_acc_1671_nl), {(fsm_output[6]) , (fsm_output[5])
      , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_579_nl = MUX1HOT_v_22_4_2(z_out_490, z_out_186_28_7, (z_out_630_29_7[21:0]),
      MultLoop_acc_206_itm, {MultLoop_or_89_cse , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[8])});
  assign nl_z_out_834 = (MultLoop_mux1h_578_nl) + (MultLoop_mux1h_579_nl);
  assign z_out_834 = nl_z_out_834[21:0];
  assign nl_MultLoop_acc_1675_nl = (z_out_873_29_7[21:0]) + (z_out_872_29_7[21:0]);
  assign MultLoop_acc_1675_nl = nl_MultLoop_acc_1675_nl[21:0];
  assign nl_MultLoop_acc_1674_nl = z_out_258 + (MultLoop_acc_1675_nl);
  assign MultLoop_acc_1674_nl = nl_MultLoop_acc_1674_nl[21:0];
  assign AccumDotWidth_mux1h_1439_nl = MUX1HOT_v_22_7_2(z_out_420, z_out_566, z_out_520,
      z_out_717, z_out_353, z_out_563, (MultLoop_acc_1674_nl), {(fsm_output[2]) ,
      (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1440_nl = MUX1HOT_v_22_7_2(z_out_710, z_out_521, MultLoop_acc_1018_itm,
      z_out_718, z_out_363, z_out_523, MultLoop_acc_861_itm, {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_835 = (AccumDotWidth_mux1h_1439_nl) + (AccumDotWidth_mux1h_1440_nl);
  assign z_out_835 = nl_z_out_835[21:0];
  assign AccumDotWidth_mux1h_1441_nl = MUX1HOT_v_22_7_2(z_out_704, z_out_178_28_7,
      z_out_156_28_7, z_out_714, MultLoop_acc_308_itm, z_out_320, z_out_564, {(fsm_output[2])
      , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1442_nl = MUX1HOT_v_22_7_2(z_out_701, z_out_174_28_7,
      z_out_664_28_7, z_out_702, z_out_514, z_out_529, MultLoop_acc_740_itm, {(fsm_output[2])
      , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_836 = (AccumDotWidth_mux1h_1441_nl) + (AccumDotWidth_mux1h_1442_nl);
  assign z_out_836 = nl_z_out_836[21:0];
  assign AccumDotWidth_mux1h_1443_nl = MUX1HOT_v_22_4_2(z_out_700, MultLoop_acc_483_itm,
      z_out_323, z_out_320, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1444_nl = MUX1HOT_v_22_4_2(z_out_707, z_out_559, z_out_527,
      z_out_327, {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_837 = (AccumDotWidth_mux1h_1443_nl) + (AccumDotWidth_mux1h_1444_nl);
  assign z_out_837 = nl_z_out_837[21:0];
  assign AccumDotWidth_mux1h_1445_nl = MUX1HOT_v_22_3_2(z_out_708, z_out_519, MultLoop_acc_435_itm,
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_156_cse});
  assign AccumDotWidth_mux1h_1446_nl = MUX1HOT_v_22_4_2(z_out_711, z_out_523, z_out_560,
      z_out_824, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign nl_z_out_838 = (AccumDotWidth_mux1h_1445_nl) + (AccumDotWidth_mux1h_1446_nl);
  assign z_out_838 = nl_z_out_838[21:0];
  assign MultLoop_mux_119_nl = MUX_v_22_2_2(z_out_171_28_7, z_out_180_28_7, fsm_output[5]);
  assign MultLoop_mux_120_nl = MUX_v_22_2_2(z_out_173_28_7, z_out_631_28_7, fsm_output[5]);
  assign nl_z_out_839 = (MultLoop_mux_119_nl) + (MultLoop_mux_120_nl);
  assign z_out_839 = nl_z_out_839[21:0];
  assign MultLoop_mux1h_580_nl = MUX1HOT_v_22_3_2(z_out_637_28_7, z_out_138_28_7,
      z_out_192_28_7, {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[4])});
  assign MultLoop_mux1h_581_nl = MUX1HOT_v_22_3_2(z_out_175_28_7, z_out_141_28_7,
      z_out_191_28_7, {(fsm_output[5]) , (fsm_output[6]) , (fsm_output[4])});
  assign nl_z_out_840 = (MultLoop_mux1h_580_nl) + (MultLoop_mux1h_581_nl);
  assign z_out_840 = nl_z_out_840[21:0];
  assign MultLoop_mux_121_nl = MUX_v_22_2_2(z_out_156_28_7, z_out_559, fsm_output[8]);
  assign MultLoop_mux_122_nl = MUX_v_22_2_2(z_out_193_28_7, MultLoop_acc_105_itm,
      fsm_output[8]);
  assign nl_z_out_841 = (MultLoop_mux_121_nl) + (MultLoop_mux_122_nl);
  assign z_out_841 = nl_z_out_841[21:0];
  assign nl_MultLoop_acc_1677_nl = (z_out_975_29_7[21:0]) + (z_out_973_29_7[21:0]);
  assign MultLoop_acc_1677_nl = nl_MultLoop_acc_1677_nl[21:0];
  assign nl_MultLoop_acc_1676_nl = z_out_852 + (MultLoop_acc_1677_nl);
  assign MultLoop_acc_1676_nl = nl_MultLoop_acc_1676_nl[21:0];
  assign MultLoop_mux1h_582_nl = MUX1HOT_v_22_8_2(z_out_166_28_7, z_out_174_28_7,
      z_out_716, z_out_521, z_out_385, z_out_327, z_out_695, (MultLoop_acc_1676_nl),
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign MultLoop_mux1h_583_nl = MUX1HOT_v_22_8_2(z_out_167_28_7, z_out_175_28_7,
      z_out_715, z_out_236, z_out_387, z_out_338, z_out_691, MultLoop_acc_333_itm,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_842 = (MultLoop_mux1h_582_nl) + (MultLoop_mux1h_583_nl);
  assign z_out_842 = nl_z_out_842[21:0];
  assign nl_MultLoop_acc_1679_nl = (z_out_871_29_7[21:0]) + (z_out_870_29_7[21:0]);
  assign MultLoop_acc_1679_nl = nl_MultLoop_acc_1679_nl[21:0];
  assign nl_MultLoop_acc_1680_nl = (z_out_869_29_7[21:0]) + (z_out_868_29_7[21:0]);
  assign MultLoop_acc_1680_nl = nl_MultLoop_acc_1680_nl[21:0];
  assign nl_MultLoop_acc_1678_nl = (MultLoop_acc_1679_nl) + (MultLoop_acc_1680_nl);
  assign MultLoop_acc_1678_nl = nl_MultLoop_acc_1678_nl[21:0];
  assign MultLoop_mux_123_nl = MUX_v_22_2_2(z_out_158_28_7, (MultLoop_acc_1678_nl),
      fsm_output[8]);
  assign MultLoop_mux_124_nl = MUX_v_22_2_2(z_out_159_28_7, z_out_324, fsm_output[8]);
  assign nl_z_out_843 = (MultLoop_mux_123_nl) + (MultLoop_mux_124_nl);
  assign z_out_843 = nl_z_out_843[21:0];
  assign nl_AccumDotWidth_acc_2722_nl = conv_s2s_21_22(z_out_862_29_7[22:2]) + conv_s2s_21_22(z_out_864_29_7[22:2])
      + conv_s2s_21_22(z_out_1187_29_7[22:2]) + conv_s2s_21_22(z_out_615_29_7[22:2]);
  assign AccumDotWidth_acc_2722_nl = nl_AccumDotWidth_acc_2722_nl[21:0];
  assign nl_AccumDotWidth_acc_2720_nl = z_out_805 + (AccumDotWidth_acc_2722_nl) +
      z_out_344;
  assign AccumDotWidth_acc_2720_nl = nl_AccumDotWidth_acc_2720_nl[21:0];
  assign AccumDotWidth_mux1h_1447_nl = MUX1HOT_v_22_8_2((AccumDotWidth_acc_2720_nl),
      z_out_251, z_out_347, z_out_714, z_out_351, z_out_315, z_out_349, AccumDotWidth_acc_1274_itm,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1448_nl = MUX1HOT_v_22_8_2(z_out_242, z_out_256, z_out_704,
      z_out_716, z_out_339, z_out_346, z_out_681, MultLoop_775_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_844 = (AccumDotWidth_mux1h_1447_nl) + (AccumDotWidth_mux1h_1448_nl);
  assign z_out_844 = nl_z_out_844[21:0];
  assign nl_MultLoop_acc_1682_nl = (z_out_957_29_7[21:0]) + (z_out_958_29_7[21:0]);
  assign MultLoop_acc_1682_nl = nl_MultLoop_acc_1682_nl[21:0];
  assign nl_MultLoop_acc_1683_nl = (z_out_959_29_7[21:0]) + MultLoop_355_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm;
  assign MultLoop_acc_1683_nl = nl_MultLoop_acc_1683_nl[21:0];
  assign nl_MultLoop_acc_1681_nl = (MultLoop_acc_1682_nl) + (MultLoop_acc_1683_nl);
  assign MultLoop_acc_1681_nl = nl_MultLoop_acc_1681_nl[21:0];
  assign MultLoop_mux1h_584_nl = MUX1HOT_v_22_3_2(z_out_172_28_7, z_out_160_28_7,
      (MultLoop_acc_1681_nl), {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_MultLoop_acc_1685_nl = MultLoop_356_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm
      + (z_out_960_29_7[21:0]);
  assign MultLoop_acc_1685_nl = nl_MultLoop_acc_1685_nl[21:0];
  assign nl_MultLoop_acc_1686_nl = (z_out_961_29_7[21:0]) + (z_out_906_29_7[21:0]);
  assign MultLoop_acc_1686_nl = nl_MultLoop_acc_1686_nl[21:0];
  assign nl_MultLoop_acc_1684_nl = (MultLoop_acc_1685_nl) + (MultLoop_acc_1686_nl);
  assign MultLoop_acc_1684_nl = nl_MultLoop_acc_1684_nl[21:0];
  assign MultLoop_mux1h_585_nl = MUX1HOT_v_22_3_2(z_out_170_28_7, z_out_161_28_7,
      (MultLoop_acc_1684_nl), {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign nl_z_out_845 = (MultLoop_mux1h_584_nl) + (MultLoop_mux1h_585_nl);
  assign z_out_845 = nl_z_out_845[21:0];
  assign MultLoop_mux1h_586_nl = MUX1HOT_v_22_4_2(z_out_544, z_out_183_28_7, z_out_677_28_7,
      z_out_844, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[4]) , (fsm_output[8])});
  assign MultLoop_mux1h_587_nl = MUX1HOT_v_22_4_2(z_out_561, z_out_117_28_7, z_out_678_28_7,
      MultLoop_acc_1012_itm, {(fsm_output[2]) , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[8])});
  assign nl_z_out_846 = (MultLoop_mux1h_586_nl) + (MultLoop_mux1h_587_nl);
  assign z_out_846 = nl_z_out_846[21:0];
  assign AccumDotWidth_mux1h_1449_nl = MUX1HOT_v_22_4_2(z_out_706, z_out_541, z_out_237,
      z_out_832, {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1450_nl = MUX1HOT_v_22_3_2(z_out_703, z_out_522, MultLoop_acc_1000_itm,
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_156_cse});
  assign nl_z_out_847 = (AccumDotWidth_mux1h_1449_nl) + (AccumDotWidth_mux1h_1450_nl);
  assign z_out_847 = nl_z_out_847[21:0];
  assign nl_AccumDotWidth_acc_2725_nl = conv_s2s_21_22(z_out_932_29_7[22:2]) + conv_s2s_21_22(z_out_928_29_7[22:2]);
  assign AccumDotWidth_acc_2725_nl = nl_AccumDotWidth_acc_2725_nl[21:0];
  assign AccumDotWidth_mux1h_1451_nl = MUX1HOT_v_22_5_2((AccumDotWidth_acc_2725_nl),
      z_out_712, z_out_702, z_out_373, z_out_379, {(fsm_output[1]) , MultLoop_or_22_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1452_nl = MUX1HOT_v_22_5_2(z_out_701, z_out_713, z_out_369,
      z_out_376, z_out_702, {AccumDotWidth_or_132_cse_1 , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_848 = (AccumDotWidth_mux1h_1451_nl) + (AccumDotWidth_mux1h_1452_nl);
  assign z_out_848 = nl_z_out_848[21:0];
  assign AccumDotWidth_mux1h_1453_nl = MUX1HOT_v_22_8_2(z_out_706, AccumDotWidth_acc_1352_itm,
      z_out_384, z_out_365, z_out_693, z_out_721, z_out_357, (z_out_998_29_7[21:0]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1454_nl = MUX1HOT_v_22_8_2(z_out_711, z_out_425, z_out_386,
      z_out_352, z_out_357, z_out_713, z_out_354, (z_out_1001_29_7[21:0]), {(fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_849 = (AccumDotWidth_mux1h_1453_nl) + (AccumDotWidth_mux1h_1454_nl);
  assign z_out_849 = nl_z_out_849[21:0];
  assign AccumDotWidth_mux1h_1455_nl = MUX1HOT_v_22_5_2(z_out_719, z_out_381, z_out_363,
      z_out_361, z_out_375, {AccumDotWidth_or_149_cse , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6])});
  assign AccumDotWidth_mux1h_1456_nl = MUX1HOT_v_22_5_2(z_out_717, z_out_383, z_out_364,
      z_out_381, z_out_715, {(fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse
      , (fsm_output[6]) , (fsm_output[7])});
  assign nl_z_out_850 = (AccumDotWidth_mux1h_1455_nl) + (AccumDotWidth_mux1h_1456_nl);
  assign z_out_850 = nl_z_out_850[21:0];
  assign AccumDotWidth_mux1h_1457_nl = MUX1HOT_v_22_4_2(z_out_362, z_out_707, z_out_720,
      (z_out_1056_29_7[21:0]), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1458_nl = MUX1HOT_v_22_4_2(z_out_357, z_out_698, z_out_721,
      (z_out_573_29_7[21:0]), {(fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign nl_z_out_851 = (AccumDotWidth_mux1h_1457_nl) + (AccumDotWidth_mux1h_1458_nl);
  assign z_out_851 = nl_z_out_851[21:0];
  assign AccumDotWidth_mux1h_1459_nl = MUX1HOT_v_22_3_2(z_out_358, z_out_698, (z_out_977_29_7[21:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign AccumDotWidth_mux1h_1460_nl = MUX1HOT_v_22_3_2(z_out_356, z_out_699, (z_out_976_29_7[21:0]),
      {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign nl_z_out_852 = (AccumDotWidth_mux1h_1459_nl) + (AccumDotWidth_mux1h_1460_nl);
  assign z_out_852 = nl_z_out_852[21:0];
  assign ConvFiltWidth_else_mux1h_923_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]),
      (w2_rsci_idat_mxwt[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]), (MultLoop_io_read_w4_rsc_cse_sva[8615:8608]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_924_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_53_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_89_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_272_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_923_nl)) *
      $signed((ConvFiltWidth_else_mux1h_924_nl)));
  assign z_out_853_29_7 = readslicef_30_23_7((mul_272_nl));
  assign ConvFiltWidth_else_mux1h_925_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]), (w2_rsci_idat_mxwt[111:104]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]),
      (MultLoop_io_read_w4_rsc_cse_sva[8607:8600]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_926_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), (input_1_rsci_idat_mxwt[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_52_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , ConvFiltWidth_else_or_752_cse
      , (fsm_output[1]) , (fsm_output[8])});
  assign mul_273_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_925_nl)) *
      $signed((ConvFiltWidth_else_mux1h_926_nl)));
  assign z_out_854_29_7 = readslicef_30_23_7((mul_273_nl));
  assign ConvFiltWidth_else_mux1h_927_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]),
      (w2_rsci_idat_mxwt[119:112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (MultLoop_io_read_w4_rsc_cse_sva[8639:8632]), {ConvFiltWidth_else_or_752_cse
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_928_nl = MUX1HOT_v_22_7_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_274_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_927_nl)) *
      $signed((ConvFiltWidth_else_mux1h_928_nl)));
  assign z_out_855_29_7 = readslicef_30_23_7((mul_274_nl));
  assign ConvFiltWidth_else_mux1h_929_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (w2_rsci_idat_mxwt[823:816]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]), (MultLoop_io_read_w4_rsc_cse_sva[8623:8616]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_152_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_930_nl = MUX1HOT_v_22_7_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_54_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_275_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_929_nl)) *
      $signed((ConvFiltWidth_else_mux1h_930_nl)));
  assign z_out_856_29_7 = readslicef_30_23_7((mul_275_nl));
  assign ConvFiltWidth_else_mux1h_931_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]),
      (w2_rsci_idat_mxwt[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (MultLoop_io_read_w4_rsc_cse_sva[8215:8208]), {(fsm_output[2]) , (fsm_output[1])
      , MultLoop_or_22_cse , (fsm_output[4]) , AccumDotWidth_or_152_cse , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_932_nl = MUX1HOT_v_22_7_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_276_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_931_nl)) *
      $signed((ConvFiltWidth_else_mux1h_932_nl)));
  assign z_out_857_29_7 = readslicef_30_23_7((mul_276_nl));
  assign ConvFiltWidth_else_mux1h_933_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[759:752]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (MultLoop_io_read_w4_rsc_cse_sva[8647:8640]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_934_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_277_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_933_nl)) *
      $signed((ConvFiltWidth_else_mux1h_934_nl)));
  assign z_out_858_29_7 = readslicef_30_23_7((mul_277_nl));
  assign ConvFiltWidth_else_mux1h_935_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]),
      (w2_rsci_idat_mxwt[695:688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (MultLoop_io_read_w4_rsc_cse_sva[8655:8648]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_936_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_278_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_935_nl)) *
      $signed((ConvFiltWidth_else_mux1h_936_nl)));
  assign z_out_859_29_7 = readslicef_30_23_7((mul_278_nl));
  assign ConvFiltWidth_else_mux1h_937_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (w2_rsci_idat_mxwt[183:176]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (MultLoop_io_read_w4_rsc_cse_sva[8631:8624]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_938_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_55_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_279_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_937_nl)) *
      $signed((ConvFiltWidth_else_mux1h_938_nl)));
  assign z_out_860_29_7 = readslicef_30_23_7((mul_279_nl));
  assign ConvFiltWidth_else_mux1h_939_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[375:368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (MultLoop_io_read_w4_rsc_cse_sva[8207:8200]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_940_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_280_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_939_nl)) *
      $signed((ConvFiltWidth_else_mux1h_940_nl)));
  assign z_out_861_29_7 = readslicef_30_23_7((mul_280_nl));
  assign ConvFiltWidth_else_mux1h_941_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]),
      (w2_rsci_idat_mxwt[375:368]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]),
      (MultLoop_io_read_w4_rsc_cse_sva[8199:8192]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_942_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_281_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_941_nl)) *
      $signed((ConvFiltWidth_else_mux1h_942_nl)));
  assign z_out_862_29_7 = readslicef_30_23_7((mul_281_nl));
  assign ConvFiltWidth_else_mux1h_943_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]),
      (w2_rsci_idat_mxwt[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (MultLoop_io_read_w4_rsc_cse_sva[7191:7184]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_944_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_282_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_943_nl)) *
      $signed((ConvFiltWidth_else_mux1h_944_nl)));
  assign z_out_863_29_7 = readslicef_30_23_7((mul_282_nl));
  assign ConvFiltWidth_else_mux1h_945_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]), (w2_rsci_idat_mxwt[567:560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (MultLoop_io_read_w4_rsc_cse_sva[7183:7176]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_946_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), (input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_730_cse , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_283_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_945_nl)) *
      $signed((ConvFiltWidth_else_mux1h_946_nl)));
  assign z_out_864_29_7 = readslicef_30_23_7((mul_283_nl));
  assign ConvFiltWidth_else_mux1h_947_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]), (MultLoop_io_read_w4_rsc_cse_sva[3695:3688]),
      {(fsm_output[1]) , ConvFiltWidth_else_or_752_cse , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_948_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[6]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign mul_284_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_947_nl)) *
      $signed((ConvFiltWidth_else_mux1h_948_nl)));
  assign z_out_865_29_7 = readslicef_30_23_7((mul_284_nl));
  assign ConvFiltWidth_else_mux1h_949_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (w2_rsci_idat_mxwt[247:240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (MultLoop_io_read_w4_rsc_cse_sva[7655:7648]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_950_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign mul_285_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_949_nl)) *
      $signed((ConvFiltWidth_else_mux1h_950_nl)));
  assign z_out_866_29_7 = readslicef_30_23_7((mul_285_nl));
  assign ConvFiltWidth_else_mux1h_951_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[631:624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]),
      (MultLoop_io_read_w4_rsc_cse_sva[7647:7640]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_952_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_286_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_951_nl)) *
      $signed((ConvFiltWidth_else_mux1h_952_nl)));
  assign z_out_867_29_7 = readslicef_30_23_7((mul_286_nl));
  assign ConvFiltWidth_else_mux1h_953_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[695:688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (MultLoop_io_read_w4_rsc_cse_sva[7639:7632]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_954_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , AccumDotWidth_or_138_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_287_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_953_nl)) *
      $signed((ConvFiltWidth_else_mux1h_954_nl)));
  assign z_out_868_29_7 = readslicef_30_23_7((mul_287_nl));
  assign ConvFiltWidth_else_mux1h_955_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[119:112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), (MultLoop_io_read_w4_rsc_cse_sva[7631:7624]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_956_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , AccumDotWidth_or_138_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_288_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_955_nl)) *
      $signed((ConvFiltWidth_else_mux1h_956_nl)));
  assign z_out_869_29_7 = readslicef_30_23_7((mul_288_nl));
  assign ConvFiltWidth_else_mux1h_957_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (MultLoop_io_read_w4_rsc_cse_sva[7623:7616]),
      {(fsm_output[1]) , AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_958_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[1011:990]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_289_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_957_nl)) *
      $signed((ConvFiltWidth_else_mux1h_958_nl)));
  assign z_out_870_29_7 = readslicef_30_23_7((mul_289_nl));
  assign ConvFiltWidth_else_mux1h_959_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]),
      (w2_rsci_idat_mxwt[823:816]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]),
      (MultLoop_io_read_w4_rsc_cse_sva[7615:7608]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_960_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]),
      (input_1_rsci_idat_mxwt[945:924]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_730_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_290_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_959_nl)) *
      $signed((ConvFiltWidth_else_mux1h_960_nl)));
  assign z_out_871_29_7 = readslicef_30_23_7((mul_290_nl));
  assign ConvFiltWidth_else_mux1h_961_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (MultLoop_io_read_w4_rsc_cse_sva[7383:7376]), {(fsm_output[2]) , (fsm_output[3])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_962_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[8])});
  assign mul_291_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_961_nl)) *
      $signed((ConvFiltWidth_else_mux1h_962_nl)));
  assign z_out_872_29_7 = readslicef_30_23_7((mul_291_nl));
  assign ConvFiltWidth_else_mux1h_963_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (w2_rsci_idat_mxwt[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (MultLoop_io_read_w4_rsc_cse_sva[7375:7368]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_964_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_2_ConvChan_1_ConvFiltHeight_1_ConvFiltWidth_2_else_slc_29_9_itm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign mul_292_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_963_nl)) *
      $signed((ConvFiltWidth_else_mux1h_964_nl)));
  assign z_out_873_29_7 = readslicef_30_23_7((mul_292_nl));
  assign ConvFiltWidth_else_mux1h_965_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]),
      (w2_rsci_idat_mxwt[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]), (MultLoop_io_read_w4_rsc_cse_sva[7367:7360]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_966_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , ConvOutHeight_1_ConvOutWidth_3_ConvFilt_6_ConvChan_2_ConvFiltHeight_2_ConvFiltWidth_2_else_slc_29_9_itm}),
      {MultLoop_or_89_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_293_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_965_nl)) *
      $signed((ConvFiltWidth_else_mux1h_966_nl)));
  assign z_out_874_29_7 = readslicef_30_23_7((mul_293_nl));
  assign ConvFiltWidth_else_mux1h_967_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]), (MultLoop_io_read_w4_rsc_cse_sva[3567:3560]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_40_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_294_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_967_nl)) *
      $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_40_nl)));
  assign z_out_875_29_7 = readslicef_30_23_7((mul_294_nl));
  assign ConvFiltWidth_else_mux1h_968_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]), (MultLoop_io_read_w4_rsc_cse_sva[3687:3680]),
      {(fsm_output[2]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_969_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , AccumDotWidth_or_138_cse
      , (fsm_output[8])});
  assign mul_295_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_968_nl)) *
      $signed((ConvFiltWidth_else_mux1h_969_nl)));
  assign z_out_876_29_7 = readslicef_30_23_7((mul_295_nl));
  assign ConvFiltWidth_else_mux1h_970_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[1103:1096]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (MultLoop_io_read_w4_rsc_cse_sva[4871:4864]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_971_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[1055:1034]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_296_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_970_nl)) *
      $signed((ConvFiltWidth_else_mux1h_971_nl)));
  assign z_out_877_29_7 = readslicef_30_23_7((mul_296_nl));
  assign ConvFiltWidth_else_mux1h_972_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (w2_rsci_idat_mxwt[503:496]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]), (MultLoop_io_read_w4_rsc_cse_sva[4863:4856]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_973_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_89_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_297_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_972_nl)) *
      $signed((ConvFiltWidth_else_mux1h_973_nl)));
  assign z_out_878_29_7 = readslicef_30_23_7((mul_297_nl));
  assign ConvFiltWidth_else_mux1h_974_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (w2_rsci_idat_mxwt[55:48]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (MultLoop_io_read_w4_rsc_cse_sva[5775:5768]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , AccumDotWidth_or_152_cse , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_975_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_89_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign mul_298_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_974_nl)) *
      $signed((ConvFiltWidth_else_mux1h_975_nl)));
  assign z_out_879_29_7 = readslicef_30_23_7((mul_298_nl));
  assign ConvFiltWidth_else_or_844_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[6]);
  assign ConvFiltWidth_else_mux1h_976_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[367:360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]),
      (MultLoop_io_read_w4_rsc_cse_sva[3583:3576]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[5]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_977_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_844_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_299_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_976_nl)) *
      $signed((ConvFiltWidth_else_mux1h_977_nl)));
  assign z_out_880_29_7 = readslicef_30_23_7((mul_299_nl));
  assign ConvFiltWidth_else_mux1h_978_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[567:560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]), (MultLoop_io_read_w4_rsc_cse_sva[2687:2680]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_979_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_25_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_300_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_978_nl)) *
      $signed((ConvFiltWidth_else_mux1h_979_nl)));
  assign z_out_881_29_7 = readslicef_30_23_7((mul_300_nl));
  assign ConvFiltWidth_else_or_847_cse = (fsm_output[6:2]!=5'b00000);
  assign ConvFiltWidth_else_mux1h_980_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[375:368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]), (MultLoop_io_read_w4_rsc_cse_sva[3551:3544]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_981_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_301_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_980_nl)) *
      $signed((ConvFiltWidth_else_mux1h_981_nl)));
  assign z_out_882_29_7 = readslicef_30_23_7((mul_301_nl));
  assign ConvFiltWidth_else_mux1h_982_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (MultLoop_io_read_w4_rsc_cse_sva[3543:3536]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_983_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_87_cse , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign mul_302_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_982_nl)) *
      $signed((ConvFiltWidth_else_mux1h_983_nl)));
  assign z_out_883_29_7 = readslicef_30_23_7((mul_302_nl));
  assign ConvFiltWidth_else_or_849_cse = (fsm_output[7:2]!=6'b000000);
  assign ConvFiltWidth_else_mux1h_984_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[759:752]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]),
      (MultLoop_io_read_w4_rsc_cse_sva[3599:3592]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_985_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_303_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_984_nl)) *
      $signed((ConvFiltWidth_else_mux1h_985_nl)));
  assign z_out_884_29_7 = readslicef_30_23_7((mul_303_nl));
  assign ConvFiltWidth_else_mux1h_986_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[351:344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]), (MultLoop_io_read_w4_rsc_cse_sva[3607:3600]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_987_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_304_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_986_nl)) *
      $signed((ConvFiltWidth_else_mux1h_987_nl)));
  assign z_out_885_29_7 = readslicef_30_23_7((mul_304_nl));
  assign ConvFiltWidth_else_mux1h_988_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]),
      (w2_rsci_idat_mxwt[543:536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]),
      (MultLoop_io_read_w4_rsc_cse_sva[3575:3568]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_989_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (input_1_rsci_idat_mxwt[725:704]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_849_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_305_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_988_nl)) *
      $signed((ConvFiltWidth_else_mux1h_989_nl)));
  assign z_out_886_29_7 = readslicef_30_23_7((mul_305_nl));
  assign ConvFiltWidth_else_mux1h_990_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[751:744]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (MultLoop_io_read_w4_rsc_cse_sva[3679:3672]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_991_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_87_cse , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign mul_306_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_990_nl)) *
      $signed((ConvFiltWidth_else_mux1h_991_nl)));
  assign z_out_887_29_7 = readslicef_30_23_7((mul_306_nl));
  assign ConvFiltWidth_else_mux1h_992_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]),
      (w2_rsci_idat_mxwt[559:552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]), (MultLoop_io_read_w4_rsc_cse_sva[3559:3552]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_993_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_844_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_307_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_992_nl)) *
      $signed((ConvFiltWidth_else_mux1h_993_nl)));
  assign z_out_888_29_7 = readslicef_30_23_7((mul_307_nl));
  assign ConvFiltWidth_else_mux1h_994_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]),
      (MultLoop_io_read_w4_rsc_cse_sva[5759:5752]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_995_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_308_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_994_nl)) *
      $signed((ConvFiltWidth_else_mux1h_995_nl)));
  assign z_out_889_29_7 = readslicef_30_23_7((mul_308_nl));
  assign ConvFiltWidth_else_mux1h_996_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]),
      (MultLoop_io_read_w4_rsc_cse_sva[5767:5760]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_997_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_309_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_996_nl)) *
      $signed((ConvFiltWidth_else_mux1h_997_nl)));
  assign z_out_890_29_7 = readslicef_30_23_7((mul_309_nl));
  assign ConvFiltWidth_else_mux1h_998_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]),
      (w2_rsci_idat_mxwt[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (MultLoop_io_read_w4_rsc_cse_sva[1871:1864]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_999_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[6]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign mul_310_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_998_nl)) *
      $signed((ConvFiltWidth_else_mux1h_999_nl)));
  assign z_out_891_29_7 = readslicef_30_23_7((mul_310_nl));
  assign ConvFiltWidth_else_mux1h_1000_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]),
      (w2_rsci_idat_mxwt[1095:1088]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (MultLoop_io_read_w4_rsc_cse_sva[7671:7664]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1001_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_311_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1000_nl))
      * $signed((ConvFiltWidth_else_mux1h_1001_nl)));
  assign z_out_892_29_7 = readslicef_30_23_7((mul_311_nl));
  assign ConvFiltWidth_else_or_861_cse = (fsm_output[7:3]!=5'b00000);
  assign ConvFiltWidth_else_mux1h_1002_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[679:672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]), (MultLoop_io_read_w4_rsc_cse_sva[1863:1856]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1003_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_312_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1002_nl))
      * $signed((ConvFiltWidth_else_mux1h_1003_nl)));
  assign z_out_893_29_7 = readslicef_30_23_7((mul_312_nl));
  assign ConvFiltWidth_else_mux1h_1004_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]),
      (w2_rsci_idat_mxwt[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]), (MultLoop_io_read_w4_rsc_cse_sva[4951:4944]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1005_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_87_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_313_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1004_nl))
      * $signed((ConvFiltWidth_else_mux1h_1005_nl)));
  assign z_out_894_29_7 = readslicef_30_23_7((mul_313_nl));
  assign ConvFiltWidth_else_mux1h_1006_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[95:88]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (MultLoop_io_read_w4_rsc_cse_sva[4943:4936]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1007_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_314_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1006_nl))
      * $signed((ConvFiltWidth_else_mux1h_1007_nl)));
  assign z_out_895_29_7 = readslicef_30_23_7((mul_314_nl));
  assign ConvFiltWidth_else_mux1h_1008_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (w2_rsci_idat_mxwt[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (MultLoop_io_read_w4_rsc_cse_sva[4935:4928]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1009_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[8])});
  assign mul_315_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1008_nl))
      * $signed((ConvFiltWidth_else_mux1h_1009_nl)));
  assign z_out_896_29_7 = readslicef_30_23_7((mul_315_nl));
  assign ConvFiltWidth_else_mux1h_1010_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[671:664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]),
      (MultLoop_io_read_w4_rsc_cse_sva[4927:4920]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1011_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[8])});
  assign mul_316_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1010_nl))
      * $signed((ConvFiltWidth_else_mux1h_1011_nl)));
  assign z_out_897_29_7 = readslicef_30_23_7((mul_316_nl));
  assign ConvFiltWidth_else_mux1h_1012_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]), (MultLoop_io_read_w4_rsc_cse_sva[4919:4912]),
      {(fsm_output[1]) , AccumDotWidth_or_157_cse , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1013_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[989:968]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_317_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1012_nl))
      * $signed((ConvFiltWidth_else_mux1h_1013_nl)));
  assign z_out_898_29_7 = readslicef_30_23_7((mul_317_nl));
  assign ConvFiltWidth_else_or_871_cse = (fsm_output[2]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1014_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]),
      (w2_rsci_idat_mxwt[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]), (MultLoop_io_read_w4_rsc_cse_sva[4911:4904]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_157_cse , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1015_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_871_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_318_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1014_nl))
      * $signed((ConvFiltWidth_else_mux1h_1015_nl)));
  assign z_out_899_29_7 = readslicef_30_23_7((mul_318_nl));
  assign ConvFiltWidth_else_mux1h_1016_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]),
      (w2_rsci_idat_mxwt[159:152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]), (MultLoop_io_read_w4_rsc_cse_sva[4903:4896]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_157_cse , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1017_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_871_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[8])});
  assign mul_319_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1016_nl))
      * $signed((ConvFiltWidth_else_mux1h_1017_nl)));
  assign z_out_900_29_7 = readslicef_30_23_7((mul_319_nl));
  assign ConvFiltWidth_else_mux1h_1018_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (MultLoop_io_read_w4_rsc_cse_sva[4879:4872]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_41_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_320_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1018_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_41_nl)));
  assign z_out_901_29_7 = readslicef_30_23_7((mul_320_nl));
  assign ConvFiltWidth_else_mux1h_1019_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[1063:1056]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]),
      (MultLoop_io_read_w4_rsc_cse_sva[6999:6992]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1020_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_321_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1019_nl))
      * $signed((ConvFiltWidth_else_mux1h_1020_nl)));
  assign z_out_902_29_7 = readslicef_30_23_7((mul_321_nl));
  assign ConvFiltWidth_else_mux1h_1021_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[999:992]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]), (MultLoop_io_read_w4_rsc_cse_sva[6991:6984]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1022_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_322_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1021_nl))
      * $signed((ConvFiltWidth_else_mux1h_1022_nl)));
  assign z_out_903_29_7 = readslicef_30_23_7((mul_322_nl));
  assign ConvFiltWidth_else_mux1h_1023_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]), {(fsm_output[3]) , (fsm_output[2])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_42_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), AccumDotWidth_or_140_cse);
  assign mul_323_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1023_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_42_nl)));
  assign z_out_904_29_9 = readslicef_30_21_9((mul_323_nl));
  assign ConvFiltWidth_else_mux1h_1024_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (w2_rsci_idat_mxwt[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (MultLoop_io_read_w4_rsc_cse_sva[6983:6976]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1025_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_871_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[8])});
  assign mul_324_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1024_nl))
      * $signed((ConvFiltWidth_else_mux1h_1025_nl)));
  assign z_out_905_29_7 = readslicef_30_23_7((mul_324_nl));
  assign ConvFiltWidth_else_mux1h_1026_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]),
      (w2_rsci_idat_mxwt[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]), (MultLoop_io_read_w4_rsc_cse_sva[2871:2864]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1027_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_87_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_325_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1026_nl))
      * $signed((ConvFiltWidth_else_mux1h_1027_nl)));
  assign z_out_906_29_7 = readslicef_30_23_7((mul_325_nl));
  assign ConvFiltWidth_else_mux1h_1028_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (MultLoop_io_read_w4_rsc_cse_sva[2879:2872]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_43_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_326_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1028_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_43_nl)));
  assign z_out_907_29_7 = readslicef_30_23_7((mul_326_nl));
  assign ConvFiltWidth_else_mux1h_1029_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]),
      (w2_rsci_idat_mxwt[351:344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (MultLoop_io_read_w4_rsc_cse_sva[2799:2792]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_157_cse , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1030_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_871_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4])
      , (fsm_output[8])});
  assign mul_327_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1029_nl))
      * $signed((ConvFiltWidth_else_mux1h_1030_nl)));
  assign z_out_908_29_7 = readslicef_30_23_7((mul_327_nl));
  assign ConvFiltWidth_else_or_882_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[6]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1031_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[207:200]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]),
      (MultLoop_io_read_w4_rsc_cse_sva[5743:5736]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1032_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_328_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1031_nl))
      * $signed((ConvFiltWidth_else_mux1h_1032_nl)));
  assign z_out_909_29_7 = readslicef_30_23_7((mul_328_nl));
  assign ConvFiltWidth_else_mux1h_1033_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[199:192]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]),
      (MultLoop_io_read_w4_rsc_cse_sva[4103:4096]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1034_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_329_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1033_nl))
      * $signed((ConvFiltWidth_else_mux1h_1034_nl)));
  assign z_out_910_29_7 = readslicef_30_23_7((mul_329_nl));
  assign ConvFiltWidth_else_mux1h_1035_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (w2_rsci_idat_mxwt[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (MultLoop_io_read_w4_rsc_cse_sva[5783:5776]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1036_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_330_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1035_nl))
      * $signed((ConvFiltWidth_else_mux1h_1036_nl)));
  assign z_out_911_29_7 = readslicef_30_23_7((mul_330_nl));
  assign ConvFiltWidth_else_mux1h_1037_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]),
      (w2_rsci_idat_mxwt[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]), (MultLoop_io_read_w4_rsc_cse_sva[5967:5960]),
      {MultLoop_or_89_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1038_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign mul_331_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1037_nl))
      * $signed((ConvFiltWidth_else_mux1h_1038_nl)));
  assign z_out_912_29_7 = readslicef_30_23_7((mul_331_nl));
  assign ConvFiltWidth_else_mux1h_1039_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[191:184]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]),
      (MultLoop_io_read_w4_rsc_cse_sva[5975:5968]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1040_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_332_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1039_nl))
      * $signed((ConvFiltWidth_else_mux1h_1040_nl)));
  assign z_out_913_29_7 = readslicef_30_23_7((mul_332_nl));
  assign ConvFiltWidth_else_mux1h_1041_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (w2_rsci_idat_mxwt[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]),
      (MultLoop_io_read_w4_rsc_cse_sva[5791:5784]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1042_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_333_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1041_nl))
      * $signed((ConvFiltWidth_else_mux1h_1042_nl)));
  assign z_out_914_29_7 = readslicef_30_23_7((mul_333_nl));
  assign ConvFiltWidth_else_or_892_cse = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1043_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]),
      (w2_rsci_idat_mxwt[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]), (MultLoop_io_read_w4_rsc_cse_sva[5799:5792]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1044_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , ConvFiltWidth_else_or_892_cse , (fsm_output[6]) , (fsm_output[8])});
  assign mul_334_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1043_nl))
      * $signed((ConvFiltWidth_else_mux1h_1044_nl)));
  assign z_out_915_29_7 = readslicef_30_23_7((mul_334_nl));
  assign ConvFiltWidth_else_mux1h_1045_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[983:976]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]),
      (MultLoop_io_read_w4_rsc_cse_sva[5751:5744]), {(fsm_output[1]) , MultLoop_or_89_cse
      , AccumDotWidth_or_139_cse , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1046_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , ConvFiltWidth_else_or_892_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign mul_335_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1045_nl))
      * $signed((ConvFiltWidth_else_mux1h_1046_nl)));
  assign z_out_916_29_7 = readslicef_30_23_7((mul_335_nl));
  assign ConvFiltWidth_else_mux1h_1047_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]), (MultLoop_io_read_w4_rsc_cse_sva[2895:2888]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_44_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_336_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1047_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_44_nl)));
  assign z_out_917_29_7 = readslicef_30_23_7((mul_336_nl));
  assign ConvFiltWidth_else_mux1h_1048_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]), (MultLoop_io_read_w4_rsc_cse_sva[2887:2880]),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1049_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_337_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1048_nl))
      * $signed((ConvFiltWidth_else_mux1h_1049_nl)));
  assign z_out_918_29_7 = readslicef_30_23_7((mul_337_nl));
  assign ConvFiltWidth_else_mux1h_1050_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (w2_rsci_idat_mxwt[15:8]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]), (MultLoop_io_read_w4_rsc_cse_sva[7679:7672]),
      {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1051_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[681:660]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_338_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1050_nl))
      * $signed((ConvFiltWidth_else_mux1h_1051_nl)));
  assign z_out_919_29_7 = readslicef_30_23_7((mul_338_nl));
  assign ConvFiltWidth_else_mux1h_1052_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[295:288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]), (MultLoop_io_read_w4_rsc_cse_sva[1767:1760]),
      {(fsm_output[1]) , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1053_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_339_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1052_nl))
      * $signed((ConvFiltWidth_else_mux1h_1053_nl)));
  assign z_out_920_29_7 = readslicef_30_23_7((mul_339_nl));
  assign ConvFiltWidth_else_mux1h_1054_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (w2_rsci_idat_mxwt[583:576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]),
      (MultLoop_io_read_w4_rsc_cse_sva[1759:1752]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1055_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_340_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1054_nl))
      * $signed((ConvFiltWidth_else_mux1h_1055_nl)));
  assign z_out_921_29_7 = readslicef_30_23_7((mul_340_nl));
  assign ConvFiltWidth_else_mux1h_1056_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]),
      (w2_rsci_idat_mxwt[591:584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]),
      (MultLoop_io_read_w4_rsc_cse_sva[7943:7936]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1057_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_89_cse , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_892_cse
      , (fsm_output[8])});
  assign mul_341_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1056_nl))
      * $signed((ConvFiltWidth_else_mux1h_1057_nl)));
  assign z_out_922_29_7 = readslicef_30_23_7((mul_341_nl));
  assign ConvFiltWidth_else_mux1h_1058_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (MultLoop_io_read_w4_rsc_cse_sva[7175:7168]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1059_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[8])});
  assign mul_342_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1058_nl))
      * $signed((ConvFiltWidth_else_mux1h_1059_nl)));
  assign z_out_923_29_7 = readslicef_30_23_7((mul_342_nl));
  assign ConvFiltWidth_else_mux1h_1060_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]),
      (w2_rsci_idat_mxwt[1079:1072]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (MultLoop_io_read_w4_rsc_cse_sva[1799:1792]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1061_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      (input_1_rsci_idat_mxwt[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_343_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1060_nl))
      * $signed((ConvFiltWidth_else_mux1h_1061_nl)));
  assign z_out_924_29_7 = readslicef_30_23_7((mul_343_nl));
  assign ConvFiltWidth_else_mux1h_1062_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[47:40]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (MultLoop_io_read_w4_rsc_cse_sva[1807:1800]), {(fsm_output[1]) , MultLoop_or_22_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1063_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_344_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1062_nl))
      * $signed((ConvFiltWidth_else_mux1h_1063_nl)));
  assign z_out_925_29_7 = readslicef_30_23_7((mul_344_nl));
  assign ConvFiltWidth_else_mux1h_1064_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[183:176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]), (MultLoop_io_read_w4_rsc_cse_sva[1831:1824]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1065_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[3]) , AccumDotWidth_or_38_cse , (fsm_output[8])});
  assign mul_345_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1064_nl))
      * $signed((ConvFiltWidth_else_mux1h_1065_nl)));
  assign z_out_926_29_7 = readslicef_30_23_7((mul_345_nl));
  assign ConvFiltWidth_else_mux1h_1066_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (w2_rsci_idat_mxwt[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]), (MultLoop_io_read_w4_rsc_cse_sva[1839:1832]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1067_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign mul_346_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1066_nl))
      * $signed((ConvFiltWidth_else_mux1h_1067_nl)));
  assign z_out_927_29_7 = readslicef_30_23_7((mul_346_nl));
  assign ConvFiltWidth_else_mux1h_1068_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[111:104]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]),
      (MultLoop_io_read_w4_rsc_cse_sva[1847:1840]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1069_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_347_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1068_nl))
      * $signed((ConvFiltWidth_else_mux1h_1069_nl)));
  assign z_out_928_29_7 = readslicef_30_23_7((mul_347_nl));
  assign ConvFiltWidth_else_mux1h_1070_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (w2_rsci_idat_mxwt[303:296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (MultLoop_io_read_w4_rsc_cse_sva[1855:1848]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1071_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[8])});
  assign mul_348_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1070_nl))
      * $signed((ConvFiltWidth_else_mux1h_1071_nl)));
  assign z_out_929_29_7 = readslicef_30_23_7((mul_348_nl));
  assign ConvFiltWidth_else_mux1h_1072_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]), (MultLoop_io_read_w4_rsc_cse_sva[1791:1784]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_45_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_349_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1072_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_45_nl)));
  assign z_out_930_29_7 = readslicef_30_23_7((mul_349_nl));
  assign ConvFiltWidth_else_mux1h_1073_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (w2_rsci_idat_mxwt[887:880]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (MultLoop_io_read_w4_rsc_cse_sva[7951:7944]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1074_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[8])});
  assign mul_350_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1073_nl))
      * $signed((ConvFiltWidth_else_mux1h_1074_nl)));
  assign z_out_931_29_7 = readslicef_30_23_7((mul_350_nl));
  assign ConvFiltWidth_else_mux1h_1075_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (w2_rsci_idat_mxwt[1007:1000]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]), (MultLoop_io_read_w4_rsc_cse_sva[6791:6784]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1076_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_351_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1075_nl))
      * $signed((ConvFiltWidth_else_mux1h_1076_nl)));
  assign z_out_932_29_7 = readslicef_30_23_7((mul_351_nl));
  assign ConvFiltWidth_else_mux1h_1077_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (w2_rsci_idat_mxwt[239:232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]),
      (MultLoop_io_read_w4_rsc_cse_sva[6799:6792]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1078_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , AccumDotWidth_or_145_cse , (fsm_output[8])});
  assign mul_352_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1077_nl))
      * $signed((ConvFiltWidth_else_mux1h_1078_nl)));
  assign z_out_933_29_7 = readslicef_30_23_7((mul_352_nl));
  assign ConvFiltWidth_else_mux1h_1079_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]), (MultLoop_io_read_w4_rsc_cse_sva[3783:3776]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_46_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}), fsm_output[8]);
  assign mul_353_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1079_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_46_nl)));
  assign z_out_934_29_7 = readslicef_30_23_7((mul_353_nl));
  assign ConvFiltWidth_else_mux1h_1080_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]),
      (w2_rsci_idat_mxwt[623:616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]),
      (MultLoop_io_read_w4_rsc_cse_sva[3855:3848]), {MultLoop_or_93_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1081_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5])
      , (fsm_output[8])});
  assign mul_354_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1080_nl))
      * $signed((ConvFiltWidth_else_mux1h_1081_nl)));
  assign z_out_935_29_7 = readslicef_30_23_7((mul_354_nl));
  assign ConvFiltWidth_else_mux1h_1082_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (w2_rsci_idat_mxwt[431:424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]),
      (MultLoop_io_read_w4_rsc_cse_sva[8807:8800]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1083_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[923:902]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[241:220]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , AccumDotWidth_or_145_cse , (fsm_output[8])});
  assign mul_355_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1082_nl))
      * $signed((ConvFiltWidth_else_mux1h_1083_nl)));
  assign z_out_936_29_7 = readslicef_30_23_7((mul_355_nl));
  assign ConvFiltWidth_else_mux1h_1084_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[431:424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]), (MultLoop_io_read_w4_rsc_cse_sva[8815:8808]),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1085_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[681:660]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_356_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1084_nl))
      * $signed((ConvFiltWidth_else_mux1h_1085_nl)));
  assign z_out_937_29_7 = readslicef_30_23_7((mul_356_nl));
  assign ConvFiltWidth_else_mux1h_1086_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]), (MultLoop_io_read_w4_rsc_cse_sva[6871:6864]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_47_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      fsm_output[8]);
  assign mul_357_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1086_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_47_nl)));
  assign z_out_938_29_7 = readslicef_30_23_7((mul_357_nl));
  assign ConvFiltWidth_else_mux1h_1087_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[815:808]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]), (MultLoop_io_read_w4_rsc_cse_sva[6951:6944]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1088_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_751_cse , (fsm_output[8])});
  assign mul_358_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1087_nl))
      * $signed((ConvFiltWidth_else_mux1h_1088_nl)));
  assign z_out_939_29_7 = readslicef_30_23_7((mul_358_nl));
  assign ConvFiltWidth_else_mux1h_1089_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (MultLoop_io_read_w4_rsc_cse_sva[3535:3528]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_or_931_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[5]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1090_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (ConvFiltWidth_else_or_931_nl) , (fsm_output[8])});
  assign mul_359_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1089_nl))
      * $signed((ConvFiltWidth_else_mux1h_1090_nl)));
  assign z_out_940_29_7 = readslicef_30_23_7((mul_359_nl));
  assign ConvFiltWidth_else_mux1h_1091_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[799:792]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]),
      (MultLoop_io_read_w4_rsc_cse_sva[3527:3520]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1092_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_360_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1091_nl))
      * $signed((ConvFiltWidth_else_mux1h_1092_nl)));
  assign z_out_941_29_7 = readslicef_30_23_7((mul_360_nl));
  assign ConvFiltWidth_else_mux1h_1093_nl = MUX1HOT_v_8_3_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (w2_rsci_idat_mxwt[631:624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1094_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (input_1_rsci_idat_mxwt[813:792]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_145_cse});
  assign mul_361_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1093_nl))
      * $signed((ConvFiltWidth_else_mux1h_1094_nl)));
  assign z_out_942_29_9 = readslicef_30_21_9((mul_361_nl));
  assign ConvFiltWidth_else_mux1h_1095_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[743:736]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]),
      (MultLoop_io_read_w4_rsc_cse_sva[3519:3512]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1096_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_362_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1095_nl))
      * $signed((ConvFiltWidth_else_mux1h_1096_nl)));
  assign z_out_943_29_7 = readslicef_30_23_7((mul_362_nl));
  assign ConvFiltWidth_else_mux1h_1097_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[359:352]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]),
      (MultLoop_io_read_w4_rsc_cse_sva[3095:3088]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1098_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_363_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1097_nl))
      * $signed((ConvFiltWidth_else_mux1h_1098_nl)));
  assign z_out_944_29_7 = readslicef_30_23_7((mul_363_nl));
  assign ConvFiltWidth_else_mux1h_1099_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]),
      (MultLoop_io_read_w4_rsc_cse_sva[3087:3080]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1100_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_364_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1099_nl))
      * $signed((ConvFiltWidth_else_mux1h_1100_nl)));
  assign z_out_945_29_7 = readslicef_30_23_7((mul_364_nl));
  assign ConvFiltWidth_else_mux1h_1101_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (w2_rsci_idat_mxwt[415:408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (MultLoop_io_read_w4_rsc_cse_sva[3079:3072]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1102_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (input_1_rsci_idat_mxwt[681:660]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {ConvFiltWidth_else_or_849_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_365_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1101_nl))
      * $signed((ConvFiltWidth_else_mux1h_1102_nl)));
  assign z_out_946_29_7 = readslicef_30_23_7((mul_365_nl));
  assign ConvFiltWidth_else_mux1h_1103_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]),
      (MultLoop_io_read_w4_rsc_cse_sva[6959:6952]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1104_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_366_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1103_nl))
      * $signed((ConvFiltWidth_else_mux1h_1104_nl)));
  assign z_out_947_29_7 = readslicef_30_23_7((mul_366_nl));
  assign ConvFiltWidth_else_mux1h_1105_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (w2_rsci_idat_mxwt[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]), (MultLoop_io_read_w4_rsc_cse_sva[6967:6960]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1106_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_367_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1105_nl))
      * $signed((ConvFiltWidth_else_mux1h_1106_nl)));
  assign z_out_948_29_7 = readslicef_30_23_7((mul_367_nl));
  assign ConvFiltWidth_else_mux1h_1107_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]), (w2_rsci_idat_mxwt[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]), (MultLoop_io_read_w4_rsc_cse_sva[6975:6968]),
      {AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[1]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1108_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]), (input_1_rsci_idat_mxwt[879:858]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_368_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1107_nl))
      * $signed((ConvFiltWidth_else_mux1h_1108_nl)));
  assign z_out_949_29_7 = readslicef_30_23_7((mul_368_nl));
  assign ConvFiltWidth_else_mux1h_1109_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[487:480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]),
      (MultLoop_io_read_w4_rsc_cse_sva[6863:6856]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1110_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]), ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_369_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1109_nl))
      * $signed((ConvFiltWidth_else_mux1h_1110_nl)));
  assign z_out_950_29_7 = readslicef_30_23_7((mul_369_nl));
  assign ConvFiltWidth_else_mux1h_1111_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]),
      (w2_rsci_idat_mxwt[103:96]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]),
      (MultLoop_io_read_w4_rsc_cse_sva[6879:6872]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1112_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      (input_1_rsci_idat_mxwt[571:550]), ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {ConvFiltWidth_else_or_849_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_370_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1111_nl))
      * $signed((ConvFiltWidth_else_mux1h_1112_nl)));
  assign z_out_951_29_7 = readslicef_30_23_7((mul_370_nl));
  assign ConvFiltWidth_else_mux1h_1113_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[855:848]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]),
      (MultLoop_io_read_w4_rsc_cse_sva[6919:6912]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1114_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_371_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1113_nl))
      * $signed((ConvFiltWidth_else_mux1h_1114_nl)));
  assign z_out_952_29_7 = readslicef_30_23_7((mul_371_nl));
  assign ConvFiltWidth_else_mux1h_1115_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (w2_rsci_idat_mxwt[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), (MultLoop_io_read_w4_rsc_cse_sva[2655:2648]),
      {(fsm_output[3]) , (fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1116_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_861_cse , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[8])});
  assign mul_372_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1115_nl))
      * $signed((ConvFiltWidth_else_mux1h_1116_nl)));
  assign z_out_953_29_7 = readslicef_30_23_7((mul_372_nl));
  assign ConvFiltWidth_else_mux1h_1117_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]), (w2_rsci_idat_mxwt[583:576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]), (MultLoop_io_read_w4_rsc_cse_sva[2783:2776]),
      {(fsm_output[2]) , MultLoop_or_22_cse , (fsm_output[1]) , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1118_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), (input_1_rsci_idat_mxwt[879:858]),
      ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[1]) , (fsm_output[8])});
  assign mul_373_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1117_nl))
      * $signed((ConvFiltWidth_else_mux1h_1118_nl)));
  assign z_out_954_29_7 = readslicef_30_23_7((mul_373_nl));
  assign ConvFiltWidth_else_mux1h_1119_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]), (w2_rsci_idat_mxwt[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (MultLoop_io_read_w4_rsc_cse_sva[2791:2784]), {(fsm_output[2]) , (fsm_output[6])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1120_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_374_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1119_nl))
      * $signed((ConvFiltWidth_else_mux1h_1120_nl)));
  assign z_out_955_29_7 = readslicef_30_23_7((mul_374_nl));
  assign ConvFiltWidth_else_mux1h_1121_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (w2_rsci_idat_mxwt[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]), (MultLoop_io_read_w4_rsc_cse_sva[2807:2800]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1122_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_375_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1121_nl))
      * $signed((ConvFiltWidth_else_mux1h_1122_nl)));
  assign z_out_956_29_7 = readslicef_30_23_7((mul_375_nl));
  assign ConvFiltWidth_else_mux1h_1123_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (w2_rsci_idat_mxwt[463:456]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]), (MultLoop_io_read_w4_rsc_cse_sva[2815:2808]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1124_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_376_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1123_nl))
      * $signed((ConvFiltWidth_else_mux1h_1124_nl)));
  assign z_out_957_29_7 = readslicef_30_23_7((mul_376_nl));
  assign ConvFiltWidth_else_mux1h_1125_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]),
      (w2_rsci_idat_mxwt[391:384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (MultLoop_io_read_w4_rsc_cse_sva[2823:2816]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1126_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_377_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1125_nl))
      * $signed((ConvFiltWidth_else_mux1h_1126_nl)));
  assign z_out_958_29_7 = readslicef_30_23_7((mul_377_nl));
  assign ConvFiltWidth_else_mux1h_1127_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (w2_rsci_idat_mxwt[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]),
      (MultLoop_io_read_w4_rsc_cse_sva[2831:2824]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1128_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_378_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1127_nl))
      * $signed((ConvFiltWidth_else_mux1h_1128_nl)));
  assign z_out_959_29_7 = readslicef_30_23_7((mul_378_nl));
  assign ConvFiltWidth_else_mux1h_1129_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]),
      (MultLoop_io_read_w4_rsc_cse_sva[2855:2848]), {(fsm_output[1]) , AccumDotWidth_or_25_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1130_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign mul_379_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1129_nl))
      * $signed((ConvFiltWidth_else_mux1h_1130_nl)));
  assign z_out_960_29_7 = readslicef_30_23_7((mul_379_nl));
  assign ConvFiltWidth_else_mux1h_1131_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[143:136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]), (MultLoop_io_read_w4_rsc_cse_sva[2863:2856]),
      {(fsm_output[1]) , AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1132_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_380_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1131_nl))
      * $signed((ConvFiltWidth_else_mux1h_1132_nl)));
  assign z_out_961_29_7 = readslicef_30_23_7((mul_380_nl));
  assign ConvFiltWidth_else_mux1h_1133_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]),
      (w2_rsci_idat_mxwt[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), {(fsm_output[2]) ,
      (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) ,
      (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1134_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[6])});
  assign mul_381_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1133_nl))
      * $signed((ConvFiltWidth_else_mux1h_1134_nl)));
  assign z_out_962_29_9 = readslicef_30_21_9((mul_381_nl));
  assign ConvFiltWidth_else_mux1h_1135_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (w2_rsci_idat_mxwt[271:264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]), {(fsm_output[2]) ,
      (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) , (fsm_output[5]) ,
      (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1136_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse});
  assign mul_382_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1135_nl))
      * $signed((ConvFiltWidth_else_mux1h_1136_nl)));
  assign z_out_963_29_9 = readslicef_30_21_9((mul_382_nl));
  assign ConvFiltWidth_else_mux1h_1137_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[623:616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]), (MultLoop_io_read_w4_rsc_cse_sva[6887:6880]),
      {(fsm_output[1]) , (fsm_output[2]) , AccumDotWidth_or_139_cse , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1138_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_383_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1137_nl))
      * $signed((ConvFiltWidth_else_mux1h_1138_nl)));
  assign z_out_964_29_7 = readslicef_30_23_7((mul_383_nl));
  assign ConvFiltWidth_else_mux1h_1139_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]),
      (w2_rsci_idat_mxwt[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]), {AccumDotWidth_or_25_cse
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1140_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse});
  assign mul_384_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1139_nl))
      * $signed((ConvFiltWidth_else_mux1h_1140_nl)));
  assign z_out_965_29_9 = readslicef_30_21_9((mul_384_nl));
  assign ConvFiltWidth_else_mux1h_1141_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]), (MultLoop_io_read_w4_rsc_cse_sva[6927:6920]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_48_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_98_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_385_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1141_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_48_nl)));
  assign z_out_966_29_7 = readslicef_30_23_7((mul_385_nl));
  assign ConvFiltWidth_else_mux1h_1142_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]), (MultLoop_io_read_w4_rsc_cse_sva[5607:5600]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_49_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[439:418]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_386_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1142_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_49_nl)));
  assign z_out_967_29_7 = readslicef_30_23_7((mul_386_nl));
  assign ConvFiltWidth_else_mux1h_1143_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]),
      (w2_rsci_idat_mxwt[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (MultLoop_io_read_w4_rsc_cse_sva[3887:3880]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1144_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_387_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1143_nl))
      * $signed((ConvFiltWidth_else_mux1h_1144_nl)));
  assign z_out_968_29_7 = readslicef_30_23_7((mul_387_nl));
  assign ConvFiltWidth_else_mux1h_1145_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]),
      (w2_rsci_idat_mxwt[23:16]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]), (MultLoop_io_read_w4_rsc_cse_sva[5135:5128]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1146_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]),
      (input_1_rsci_idat_mxwt[549:528]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_388_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1145_nl))
      * $signed((ConvFiltWidth_else_mux1h_1146_nl)));
  assign z_out_969_29_7 = readslicef_30_23_7((mul_388_nl));
  assign ConvFiltWidth_else_mux1h_1147_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (w2_rsci_idat_mxwt[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]), (MultLoop_io_read_w4_rsc_cse_sva[5143:5136]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1148_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_389_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1147_nl))
      * $signed((ConvFiltWidth_else_mux1h_1148_nl)));
  assign z_out_970_29_7 = readslicef_30_23_7((mul_389_nl));
  assign ConvFiltWidth_else_mux1h_1149_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[47:40]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]),
      (MultLoop_io_read_w4_rsc_cse_sva[5127:5120]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1150_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_390_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1149_nl))
      * $signed((ConvFiltWidth_else_mux1h_1150_nl)));
  assign z_out_971_29_7 = readslicef_30_23_7((mul_390_nl));
  assign ConvFiltWidth_else_mux1h_1151_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[55:48]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]), (MultLoop_io_read_w4_rsc_cse_sva[5567:5560]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1152_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_391_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1151_nl))
      * $signed((ConvFiltWidth_else_mux1h_1152_nl)));
  assign z_out_972_29_7 = readslicef_30_23_7((mul_391_nl));
  assign ConvFiltWidth_else_mux1h_1153_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]),
      (w2_rsci_idat_mxwt[31:24]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (MultLoop_io_read_w4_rsc_cse_sva[3927:3920]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1154_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]),
      (input_1_rsci_idat_mxwt[549:528]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_392_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1153_nl))
      * $signed((ConvFiltWidth_else_mux1h_1154_nl)));
  assign z_out_973_29_7 = readslicef_30_23_7((mul_392_nl));
  assign ConvFiltWidth_else_mux1h_1155_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[39:32]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]), (MultLoop_io_read_w4_rsc_cse_sva[3895:3888]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1156_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_393_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1155_nl))
      * $signed((ConvFiltWidth_else_mux1h_1156_nl)));
  assign z_out_974_29_7 = readslicef_30_23_7((mul_393_nl));
  assign ConvFiltWidth_else_mux1h_1157_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]),
      (MultLoop_io_read_w4_rsc_cse_sva[3919:3912]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_50_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_106_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_394_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1157_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_50_nl)));
  assign z_out_975_29_7 = readslicef_30_23_7((mul_394_nl));
  assign ConvFiltWidth_else_or_987_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1158_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (w2_rsci_idat_mxwt[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]),
      (MultLoop_io_read_w4_rsc_cse_sva[3911:3904]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1159_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (input_1_rsci_idat_mxwt[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_987_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_395_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1158_nl))
      * $signed((ConvFiltWidth_else_mux1h_1159_nl)));
  assign z_out_976_29_7 = readslicef_30_23_7((mul_395_nl));
  assign ConvFiltWidth_else_mux1h_1160_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]),
      (MultLoop_io_read_w4_rsc_cse_sva[3903:3896]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_51_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_396_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1160_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_51_nl)));
  assign z_out_977_29_7 = readslicef_30_23_7((mul_396_nl));
  assign ConvFiltWidth_else_mux1h_1161_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]),
      (w2_rsci_idat_mxwt[79:72]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_or_989_nl = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1162_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (input_1_rsci_idat_mxwt[571:550]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (ConvFiltWidth_else_or_989_nl)});
  assign mul_397_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1161_nl))
      * $signed((ConvFiltWidth_else_mux1h_1162_nl)));
  assign z_out_978_29_9 = readslicef_30_21_9((mul_397_nl));
  assign ConvFiltWidth_else_mux1h_1163_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]),
      (w2_rsci_idat_mxwt[1119:1112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1164_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse});
  assign mul_398_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1163_nl))
      * $signed((ConvFiltWidth_else_mux1h_1164_nl)));
  assign z_out_979_29_9 = readslicef_30_21_9((mul_398_nl));
  assign ConvFiltWidth_else_mux1h_1165_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (w2_rsci_idat_mxwt[1047:1040]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]), (MultLoop_io_read_w4_rsc_cse_sva[6615:6608]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1166_nl = MUX1HOT_v_22_7_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse , (fsm_output[4])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_399_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1165_nl))
      * $signed((ConvFiltWidth_else_mux1h_1166_nl)));
  assign z_out_980_29_7 = readslicef_30_23_7((mul_399_nl));
  assign ConvFiltWidth_else_mux1h_1167_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]),
      (w2_rsci_idat_mxwt[79:72]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (MultLoop_io_read_w4_rsc_cse_sva[6607:6600]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1168_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (input_1_rsci_idat_mxwt[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_400_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1167_nl))
      * $signed((ConvFiltWidth_else_mux1h_1168_nl)));
  assign z_out_981_29_7 = readslicef_30_23_7((mul_400_nl));
  assign ConvFiltWidth_else_mux1h_1169_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (w2_rsci_idat_mxwt[975:968]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]),
      (MultLoop_io_read_w4_rsc_cse_sva[6599:6592]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1170_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_401_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1169_nl))
      * $signed((ConvFiltWidth_else_mux1h_1170_nl)));
  assign z_out_982_29_7 = readslicef_30_23_7((mul_401_nl));
  assign ConvFiltWidth_else_mux1h_1171_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (w2_rsci_idat_mxwt[15:8]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (MultLoop_io_read_w4_rsc_cse_sva[6591:6584]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1172_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_402_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1171_nl))
      * $signed((ConvFiltWidth_else_mux1h_1172_nl)));
  assign z_out_983_29_7 = readslicef_30_23_7((mul_402_nl));
  assign ConvFiltWidth_else_mux1h_1173_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]), (w2_rsci_idat_mxwt[207:200]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (MultLoop_io_read_w4_rsc_cse_sva[6167:6160]),
      {(fsm_output[2]) , (fsm_output[6]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1174_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , AccumDotWidth_or_38_cse
      , (fsm_output[8])});
  assign mul_403_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1173_nl))
      * $signed((ConvFiltWidth_else_mux1h_1174_nl)));
  assign z_out_984_29_7 = readslicef_30_23_7((mul_403_nl));
  assign ConvFiltWidth_else_mux1h_1175_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[151:144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]),
      (MultLoop_io_read_w4_rsc_cse_sva[6159:6152]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1176_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_404_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1175_nl))
      * $signed((ConvFiltWidth_else_mux1h_1176_nl)));
  assign z_out_985_29_7 = readslicef_30_23_7((mul_404_nl));
  assign ConvFiltWidth_else_mux1h_1177_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]),
      (MultLoop_io_read_w4_rsc_cse_sva[6151:6144]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1178_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]), ({1'b0 , ConvOutHeight_3_ConvOutWidth_1_ConvFilt_6_ConvChan_3_ConvFiltHeight_3_ConvFiltWidth_3_else_slc_29_9_itm}),
      {ConvFiltWidth_else_or_752_cse , AccumDotWidth_or_38_cse , (fsm_output[8])});
  assign mul_405_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1177_nl))
      * $signed((ConvFiltWidth_else_mux1h_1178_nl)));
  assign z_out_986_29_7 = readslicef_30_23_7((mul_405_nl));
  assign ConvFiltWidth_else_mux1h_1179_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (w2_rsci_idat_mxwt[591:584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (MultLoop_io_read_w4_rsc_cse_sva[2903:2896]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1180_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (input_1_rsci_idat_mxwt[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_107_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_38_cse
      , (fsm_output[8])});
  assign mul_406_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1179_nl))
      * $signed((ConvFiltWidth_else_mux1h_1180_nl)));
  assign z_out_987_29_7 = readslicef_30_23_7((mul_406_nl));
  assign ConvFiltWidth_else_mux1h_1181_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1182_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]), {(fsm_output[1])
      , (fsm_output[3]) , AccumDotWidth_or_38_cse , (fsm_output[7])});
  assign mul_407_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1181_nl))
      * $signed((ConvFiltWidth_else_mux1h_1182_nl)));
  assign z_out_988_29_9 = readslicef_30_21_9((mul_407_nl));
  assign ConvFiltWidth_else_mux1h_1183_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]), (w2_rsci_idat_mxwt[855:848]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]), {(fsm_output[4]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1184_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]), (input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), {(fsm_output[4])
      , (fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])});
  assign mul_408_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1183_nl))
      * $signed((ConvFiltWidth_else_mux1h_1184_nl)));
  assign z_out_989_29_9 = readslicef_30_21_9((mul_408_nl));
  assign ConvFiltWidth_else_mux1h_1185_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1047:1040]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]), (MultLoop_io_read_w4_rsc_cse_sva[6895:6888]),
      {(fsm_output[1]) , (fsm_output[2]) , AccumDotWidth_or_157_cse , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1186_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_409_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1185_nl))
      * $signed((ConvFiltWidth_else_mux1h_1186_nl)));
  assign z_out_990_29_7 = readslicef_30_23_7((mul_409_nl));
  assign ConvFiltWidth_else_mux1h_1187_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (w2_rsci_idat_mxwt[239:232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]), (MultLoop_io_read_w4_rsc_cse_sva[5599:5592]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1188_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      (input_1_rsci_idat_mxwt[615:594]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_410_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1187_nl))
      * $signed((ConvFiltWidth_else_mux1h_1188_nl)));
  assign z_out_991_29_7 = readslicef_30_23_7((mul_410_nl));
  assign ConvFiltWidth_else_mux1h_1189_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]),
      (w2_rsci_idat_mxwt[399:392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1190_nl = MUX1HOT_v_22_7_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[879:858]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign mul_411_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1189_nl))
      * $signed((ConvFiltWidth_else_mux1h_1190_nl)));
  assign z_out_992_29_9 = readslicef_30_21_9((mul_411_nl));
  assign ConvFiltWidth_else_mux1h_1191_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      {(fsm_output[2]) , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_11_cse
      , (fsm_output[5]) , (fsm_output[6])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_52_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse);
  assign mul_412_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1191_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_52_nl)));
  assign z_out_993_29_9 = readslicef_30_21_9((mul_412_nl));
  assign ConvFiltWidth_else_mux1h_1192_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]),
      (w2_rsci_idat_mxwt[671:664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]), (MultLoop_io_read_w4_rsc_cse_sva[1703:1696]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_22_cse , (fsm_output[4]) ,
      (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1193_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_413_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1192_nl))
      * $signed((ConvFiltWidth_else_mux1h_1193_nl)));
  assign z_out_994_29_7 = readslicef_30_23_7((mul_413_nl));
  assign ConvFiltWidth_else_mux1h_1194_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]), (w2_rsci_idat_mxwt[991:984]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[119:112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (MultLoop_io_read_w4_rsc_cse_sva[1783:1776]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1195_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), (input_1_rsci_idat_mxwt[1011:990]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[1]) , (fsm_output[8])});
  assign mul_414_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1194_nl))
      * $signed((ConvFiltWidth_else_mux1h_1195_nl)));
  assign z_out_995_29_7 = readslicef_30_23_7((mul_414_nl));
  assign ConvFiltWidth_else_mux1h_1196_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]),
      (w2_rsci_idat_mxwt[479:472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (MultLoop_io_read_w4_rsc_cse_sva[1775:1768]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1197_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_415_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1196_nl))
      * $signed((ConvFiltWidth_else_mux1h_1197_nl)));
  assign z_out_996_29_7 = readslicef_30_23_7((mul_415_nl));
  assign ConvFiltWidth_else_mux1h_1198_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]),
      (w2_rsci_idat_mxwt[223:216]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[111:104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]),
      (MultLoop_io_read_w4_rsc_cse_sva[1711:1704]), {MultLoop_or_22_cse , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1199_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_416_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1198_nl))
      * $signed((ConvFiltWidth_else_mux1h_1199_nl)));
  assign z_out_997_29_7 = readslicef_30_23_7((mul_416_nl));
  assign ConvFiltWidth_else_or_1020_cse = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1200_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[863:856]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[103:96]), (MultLoop_io_read_w4_rsc_cse_sva[1727:1720]),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1020_cse , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1201_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_417_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1200_nl))
      * $signed((ConvFiltWidth_else_mux1h_1201_nl)));
  assign z_out_998_29_7 = readslicef_30_23_7((mul_417_nl));
  assign ConvFiltWidth_else_mux1h_1202_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]),
      (MultLoop_io_read_w4_rsc_cse_sva[1751:1744]), {(fsm_output[2]) , AccumDotWidth_or_157_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1203_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {ConvFiltWidth_else_or_752_cse , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_418_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1202_nl))
      * $signed((ConvFiltWidth_else_mux1h_1203_nl)));
  assign z_out_999_29_7 = readslicef_30_23_7((mul_418_nl));
  assign ConvFiltWidth_else_mux1h_1204_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]),
      (w2_rsci_idat_mxwt[95:88]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]), (MultLoop_io_read_w4_rsc_cse_sva[1719:1712]),
      {ConvFiltWidth_else_or_1020_cse , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1205_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_419_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1204_nl))
      * $signed((ConvFiltWidth_else_mux1h_1205_nl)));
  assign z_out_1000_29_7 = readslicef_30_23_7((mul_419_nl));
  assign ConvFiltWidth_else_mux1h_1206_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (MultLoop_io_read_w4_rsc_cse_sva[1735:1728]), {(fsm_output[1]) , MultLoop_or_22_cse
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1207_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}), {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_420_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1206_nl))
      * $signed((ConvFiltWidth_else_mux1h_1207_nl)));
  assign z_out_1001_29_7 = readslicef_30_23_7((mul_420_nl));
  assign ConvFiltWidth_else_mux1h_1208_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]),
      (w2_rsci_idat_mxwt[415:408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (MultLoop_io_read_w4_rsc_cse_sva[1743:1736]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1209_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}), {ConvFiltWidth_else_or_752_cse
      , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_421_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1208_nl))
      * $signed((ConvFiltWidth_else_mux1h_1209_nl)));
  assign z_out_1002_29_7 = readslicef_30_23_7((mul_421_nl));
  assign ConvFiltWidth_else_mux1h_1210_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]),
      (w2_rsci_idat_mxwt[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1211_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse});
  assign mul_422_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1210_nl))
      * $signed((ConvFiltWidth_else_mux1h_1211_nl)));
  assign z_out_1003_29_9 = readslicef_30_21_9((mul_422_nl));
  assign ConvFiltWidth_else_mux1h_1212_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]),
      (w2_rsci_idat_mxwt[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1213_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[1]) , (fsm_output[2]) , (fsm_output[6])});
  assign mul_423_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1212_nl))
      * $signed((ConvFiltWidth_else_mux1h_1213_nl)));
  assign z_out_1004_29_9 = readslicef_30_21_9((mul_423_nl));
  assign ConvFiltWidth_else_mux1h_1214_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[991:984]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]),
      (MultLoop_io_read_w4_rsc_cse_sva[5591:5584]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1215_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign mul_424_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1214_nl))
      * $signed((ConvFiltWidth_else_mux1h_1215_nl)));
  assign z_out_1005_29_7 = readslicef_30_23_7((mul_424_nl));
  assign ConvFiltWidth_else_mux1h_1216_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[87:80]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_53_nl = MUX_v_22_2_2((input_1_rsci_idat_mxwt[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]), nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse);
  assign mul_425_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1216_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_53_nl)));
  assign z_out_1006_29_9 = readslicef_30_21_9((mul_425_nl));
  assign ConvFiltWidth_else_mux1h_1217_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (MultLoop_io_read_w4_rsc_cse_sva[5615:5608]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_54_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_426_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1217_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_54_nl)));
  assign z_out_1007_29_7 = readslicef_30_23_7((mul_426_nl));
  assign ConvFiltWidth_else_mux1h_1218_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]), (w2_rsci_idat_mxwt[335:328]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (MultLoop_io_read_w4_rsc_cse_sva[7911:7904]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[3]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1219_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]), (input_1_rsci_idat_mxwt[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[1]) , (fsm_output[8])});
  assign mul_427_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1218_nl))
      * $signed((ConvFiltWidth_else_mux1h_1219_nl)));
  assign z_out_1008_29_7 = readslicef_30_23_7((mul_427_nl));
  assign ConvFiltWidth_else_mux1h_1220_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]),
      (w2_rsci_idat_mxwt[727:720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]), (MultLoop_io_read_w4_rsc_cse_sva[7935:7928]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1221_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (input_1_rsci_idat_mxwt[923:902]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_847_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_428_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1220_nl))
      * $signed((ConvFiltWidth_else_mux1h_1221_nl)));
  assign z_out_1009_29_7 = readslicef_30_23_7((mul_428_nl));
  assign ConvFiltWidth_else_mux1h_1222_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]),
      (w2_rsci_idat_mxwt[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (MultLoop_io_read_w4_rsc_cse_sva[7999:7992]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1223_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_104_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_429_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1222_nl))
      * $signed((ConvFiltWidth_else_mux1h_1223_nl)));
  assign z_out_1010_29_7 = readslicef_30_23_7((mul_429_nl));
  assign ConvFiltWidth_else_mux1h_1224_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]), (MultLoop_io_read_w4_rsc_cse_sva[7919:7912]),
      {(fsm_output[2]) , (fsm_output[3]) , AccumDotWidth_or_145_cse , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1225_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_430_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1224_nl))
      * $signed((ConvFiltWidth_else_mux1h_1225_nl)));
  assign z_out_1011_29_7 = readslicef_30_23_7((mul_430_nl));
  assign ConvFiltWidth_else_mux1h_1226_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[575:568]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]),
      (MultLoop_io_read_w4_rsc_cse_sva[7983:7976]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1227_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_102_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_431_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1226_nl))
      * $signed((ConvFiltWidth_else_mux1h_1227_nl)));
  assign z_out_1012_29_7 = readslicef_30_23_7((mul_431_nl));
  assign ConvFiltWidth_else_mux1h_1228_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (w2_rsci_idat_mxwt[767:760]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]), (MultLoop_io_read_w4_rsc_cse_sva[7927:7920]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1229_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_432_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1228_nl))
      * $signed((ConvFiltWidth_else_mux1h_1229_nl)));
  assign z_out_1013_29_7 = readslicef_30_23_7((mul_432_nl));
  assign ConvFiltWidth_else_mux1h_1230_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[343:336]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]), (MultLoop_io_read_w4_rsc_cse_sva[7991:7984]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , AccumDotWidth_or_145_cse
      , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1231_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_103_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_752_cse , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_433_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1230_nl))
      * $signed((ConvFiltWidth_else_mux1h_1231_nl)));
  assign z_out_1014_29_7 = readslicef_30_23_7((mul_433_nl));
  assign ConvFiltWidth_else_mux1h_1232_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (w2_rsci_idat_mxwt[735:728]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]), (MultLoop_io_read_w4_rsc_cse_sva[8007:8000]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1233_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_105_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_434_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1232_nl))
      * $signed((ConvFiltWidth_else_mux1h_1233_nl)));
  assign z_out_1015_29_7 = readslicef_30_23_7((mul_434_nl));
  assign ConvFiltWidth_else_mux1h_1234_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (w2_rsci_idat_mxwt[383:376]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (MultLoop_io_read_w4_rsc_cse_sva[7975:7968]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1235_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_435_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1234_nl))
      * $signed((ConvFiltWidth_else_mux1h_1235_nl)));
  assign z_out_1016_29_7 = readslicef_30_23_7((mul_435_nl));
  assign ConvFiltWidth_else_mux1h_1236_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[535:528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1237_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , ConvFiltWidth_else_or_730_cse});
  assign mul_436_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1236_nl))
      * $signed((ConvFiltWidth_else_mux1h_1237_nl)));
  assign z_out_1017_29_9 = readslicef_30_21_9((mul_436_nl));
  assign ConvFiltWidth_else_mux1h_1238_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (w2_rsci_idat_mxwt[959:952]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]), {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1239_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[989:968]), {(fsm_output[2])
      , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])});
  assign mul_437_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1238_nl))
      * $signed((ConvFiltWidth_else_mux1h_1239_nl)));
  assign z_out_1018_29_9 = readslicef_30_21_9((mul_437_nl));
  assign ConvFiltWidth_else_mux1h_1240_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[151:144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]), (MultLoop_io_read_w4_rsc_cse_sva[5583:5576]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1241_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_438_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1240_nl))
      * $signed((ConvFiltWidth_else_mux1h_1241_nl)));
  assign z_out_1019_29_7 = readslicef_30_23_7((mul_438_nl));
  assign ConvFiltWidth_else_mux1h_1242_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (w2_rsci_idat_mxwt[919:912]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]), {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1243_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[197:176]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), {(fsm_output[2])
      , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])});
  assign mul_439_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1242_nl))
      * $signed((ConvFiltWidth_else_mux1h_1243_nl)));
  assign z_out_1020_29_9 = readslicef_30_21_9((mul_439_nl));
  assign ConvFiltWidth_else_mux1h_1244_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[95:88]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]),
      (MultLoop_io_read_w4_rsc_cse_sva[5623:5616]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1245_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign mul_440_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1244_nl))
      * $signed((ConvFiltWidth_else_mux1h_1245_nl)));
  assign z_out_1021_29_7 = readslicef_30_23_7((mul_440_nl));
  assign ConvFiltWidth_else_mux1h_1246_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]),
      (MultLoop_io_read_w4_rsc_cse_sva[6855:6848]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1247_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]), ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_441_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1246_nl))
      * $signed((ConvFiltWidth_else_mux1h_1247_nl)));
  assign z_out_1022_29_7 = readslicef_30_23_7((mul_441_nl));
  assign ConvFiltWidth_else_mux1h_1248_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[1071:1064]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]),
      (MultLoop_io_read_w4_rsc_cse_sva[6847:6840]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1249_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}), {(fsm_output[1]) , (fsm_output[2])
      , ConvFiltWidth_else_or_751_cse , (fsm_output[8])});
  assign mul_442_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1248_nl))
      * $signed((ConvFiltWidth_else_mux1h_1249_nl)));
  assign z_out_1023_29_7 = readslicef_30_23_7((mul_442_nl));
  assign ConvFiltWidth_else_mux1h_1250_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]),
      (w2_rsci_idat_mxwt[311:304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]),
      (MultLoop_io_read_w4_rsc_cse_sva[6839:6832]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1251_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (input_1_rsci_idat_mxwt[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_443_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1250_nl))
      * $signed((ConvFiltWidth_else_mux1h_1251_nl)));
  assign z_out_1024_29_7 = readslicef_30_23_7((mul_443_nl));
  assign ConvFiltWidth_else_mux1h_1252_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (w2_rsci_idat_mxwt[1015:1008]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]),
      (MultLoop_io_read_w4_rsc_cse_sva[6831:6824]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1253_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_444_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1252_nl))
      * $signed((ConvFiltWidth_else_mux1h_1253_nl)));
  assign z_out_1025_29_7 = readslicef_30_23_7((mul_444_nl));
  assign ConvFiltWidth_else_mux1h_1254_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[1079:1072]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]),
      (MultLoop_io_read_w4_rsc_cse_sva[6823:6816]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1255_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]), ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_445_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1254_nl))
      * $signed((ConvFiltWidth_else_mux1h_1255_nl)));
  assign z_out_1026_29_7 = readslicef_30_23_7((mul_445_nl));
  assign ConvFiltWidth_else_mux1h_1256_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (w2_rsci_idat_mxwt[695:688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]),
      (MultLoop_io_read_w4_rsc_cse_sva[6775:6768]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1257_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (input_1_rsci_idat_mxwt[835:814]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_446_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1256_nl))
      * $signed((ConvFiltWidth_else_mux1h_1257_nl)));
  assign z_out_1027_29_7 = readslicef_30_23_7((mul_446_nl));
  assign ConvFiltWidth_else_mux1h_1258_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]), (MultLoop_io_read_w4_rsc_cse_sva[6815:6808]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_55_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_447_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1258_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_55_nl)));
  assign z_out_1028_29_7 = readslicef_30_23_7((mul_447_nl));
  assign ConvFiltWidth_else_mux1h_1259_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[175:168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (MultLoop_io_read_w4_rsc_cse_sva[6783:6776]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1260_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_448_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1259_nl))
      * $signed((ConvFiltWidth_else_mux1h_1260_nl)));
  assign z_out_1029_29_7 = readslicef_30_23_7((mul_448_nl));
  assign ConvFiltWidth_else_mux1h_1261_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (w2_rsci_idat_mxwt[119:112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]),
      (MultLoop_io_read_w4_rsc_cse_sva[6807:6800]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1262_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[571:550]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_449_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1261_nl))
      * $signed((ConvFiltWidth_else_mux1h_1262_nl)));
  assign z_out_1030_29_7 = readslicef_30_23_7((mul_449_nl));
  assign ConvFiltWidth_else_mux1h_1263_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign mul_450_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1263_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440])));
  assign z_out_1031_29_9 = readslicef_30_21_9((mul_450_nl));
  assign ConvFiltWidth_else_mux1h_1264_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[183:176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_56_nl = MUX_v_22_2_2((input_1_rsci_idat_mxwt[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]), ConvFiltWidth_else_or_861_cse);
  assign mul_451_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1264_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_56_nl)));
  assign z_out_1032_29_9 = readslicef_30_21_9((mul_451_nl));
  assign ConvFiltWidth_else_mux1h_1265_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[503:496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[527:520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_57_nl = MUX_v_22_2_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]), ConvFiltWidth_else_or_849_cse);
  assign mul_452_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1265_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_57_nl)));
  assign z_out_1033_29_9 = readslicef_30_21_9((mul_452_nl));
  assign ConvFiltWidth_else_mux1h_1266_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[279:272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]),
      (MultLoop_io_read_w4_rsc_cse_sva[5655:5648]), {(fsm_output[1]) , AccumDotWidth_or_157_cse
      , (fsm_output[2]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1267_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[3]) , MultLoop_or_93_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_453_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1266_nl))
      * $signed((ConvFiltWidth_else_mux1h_1267_nl)));
  assign z_out_1034_29_7 = readslicef_30_23_7((mul_453_nl));
  assign ConvFiltWidth_else_or_1081_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5])
      | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1268_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[663:656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (MultLoop_io_read_w4_rsc_cse_sva[5631:5624]), {(fsm_output[1]) , (fsm_output[2])
      , AccumDotWidth_or_139_cse , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1269_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1081_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_454_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1268_nl))
      * $signed((ConvFiltWidth_else_mux1h_1269_nl)));
  assign z_out_1035_29_7 = readslicef_30_23_7((mul_454_nl));
  assign ConvFiltWidth_else_mux1h_1270_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1343:1336]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[567:560]), (MultLoop_io_read_w4_rsc_cse_sva[3815:3808]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1271_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_455_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1270_nl))
      * $signed((ConvFiltWidth_else_mux1h_1271_nl)));
  assign z_out_1036_29_7 = readslicef_30_23_7((mul_455_nl));
  assign ConvFiltWidth_else_mux1h_1272_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[271:264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]), (MultLoop_io_read_w4_rsc_cse_sva[3879:3872]),
      {(fsm_output[1]) , (fsm_output[2]) , AccumDotWidth_or_157_cse , (fsm_output[5])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1273_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_101_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[8])});
  assign mul_456_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1272_nl))
      * $signed((ConvFiltWidth_else_mux1h_1273_nl)));
  assign z_out_1037_29_7 = readslicef_30_23_7((mul_456_nl));
  assign ConvFiltWidth_else_mux1h_1274_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[463:456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[535:528]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (MultLoop_io_read_w4_rsc_cse_sva[3847:3840]), {(fsm_output[1]) , (fsm_output[2])
      , AccumDotWidth_or_157_cse , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1275_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_97_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_457_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1274_nl))
      * $signed((ConvFiltWidth_else_mux1h_1275_nl)));
  assign z_out_1038_29_7 = readslicef_30_23_7((mul_457_nl));
  assign ConvFiltWidth_else_mux1h_1276_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1119:1112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[559:552]), (MultLoop_io_read_w4_rsc_cse_sva[3831:3824]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1277_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_458_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1276_nl))
      * $signed((ConvFiltWidth_else_mux1h_1277_nl)));
  assign z_out_1039_29_7 = readslicef_30_23_7((mul_458_nl));
  assign ConvFiltWidth_else_mux1h_1278_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[727:720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[551:544]), (MultLoop_io_read_w4_rsc_cse_sva[3791:3784]),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1279_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[857:836]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}), {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse
      , (fsm_output[3]) , (fsm_output[8])});
  assign mul_459_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1278_nl))
      * $signed((ConvFiltWidth_else_mux1h_1279_nl)));
  assign z_out_1040_29_7 = readslicef_30_23_7((mul_459_nl));
  assign ConvFiltWidth_else_mux1h_1280_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1151:1144]),
      (w2_rsci_idat_mxwt[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]),
      (MultLoop_io_read_w4_rsc_cse_sva[3799:3792]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1281_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign mul_460_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1280_nl))
      * $signed((ConvFiltWidth_else_mux1h_1281_nl)));
  assign z_out_1041_29_7 = readslicef_30_23_7((mul_460_nl));
  assign ConvFiltWidth_else_mux1h_1282_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[407:400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1143:1136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]),
      (MultLoop_io_read_w4_rsc_cse_sva[3839:3832]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1283_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[681:660]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_461_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1282_nl))
      * $signed((ConvFiltWidth_else_mux1h_1283_nl)));
  assign z_out_1042_29_7 = readslicef_30_23_7((mul_461_nl));
  assign ConvFiltWidth_else_mux1h_1284_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[599:592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1703:1696]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]),
      (MultLoop_io_read_w4_rsc_cse_sva[3807:3800]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1285_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_462_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1284_nl))
      * $signed((ConvFiltWidth_else_mux1h_1285_nl)));
  assign z_out_1043_29_7 = readslicef_30_23_7((mul_462_nl));
  assign ConvFiltWidth_else_mux1h_1286_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[343:336]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1711:1704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]), (MultLoop_io_read_w4_rsc_cse_sva[3823:3816]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1287_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[659:638]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[8])});
  assign mul_463_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1286_nl))
      * $signed((ConvFiltWidth_else_mux1h_1287_nl)));
  assign z_out_1044_29_7 = readslicef_30_23_7((mul_463_nl));
  assign ConvFiltWidth_else_mux1h_1288_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]),
      (w2_rsci_idat_mxwt[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]), (MultLoop_io_read_w4_rsc_cse_sva[5735:5728]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1289_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]),
      (input_1_rsci_idat_mxwt[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_464_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1288_nl))
      * $signed((ConvFiltWidth_else_mux1h_1289_nl)));
  assign z_out_1045_29_7 = readslicef_30_23_7((mul_464_nl));
  assign ConvFiltWidth_else_mux1h_1290_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1719:1712]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]),
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign mul_465_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1290_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638])));
  assign z_out_1046_29_9 = readslicef_30_21_9((mul_465_nl));
  assign ConvFiltWidth_else_mux1h_1291_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[535:528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1727:1720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]), {(fsm_output[1]) , (fsm_output[2])
      , AccumDotWidth_or_139_cse , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1292_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      {(fsm_output[1]) , ConvFiltWidth_else_or_882_cse , (fsm_output[3])});
  assign mul_466_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1291_nl))
      * $signed((ConvFiltWidth_else_mux1h_1292_nl)));
  assign z_out_1047_29_9 = readslicef_30_21_9((mul_466_nl));
  assign ConvFiltWidth_else_mux1h_1293_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[543:536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1294_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1081_cse , (fsm_output[3])});
  assign mul_467_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1293_nl))
      * $signed((ConvFiltWidth_else_mux1h_1294_nl)));
  assign z_out_1048_29_9 = readslicef_30_21_9((mul_467_nl));
  assign ConvFiltWidth_else_mux1h_1295_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[479:472]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]), (MultLoop_io_read_w4_rsc_cse_sva[5647:5640]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1296_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1081_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_468_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1295_nl))
      * $signed((ConvFiltWidth_else_mux1h_1296_nl)));
  assign z_out_1049_29_7 = readslicef_30_23_7((mul_468_nl));
  assign ConvFiltWidth_else_mux1h_1297_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (MultLoop_io_read_w4_rsc_cse_sva[8783:8776]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1298_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_74_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , ConvFiltWidth_else_or_730_cse
      , (fsm_output[8])});
  assign mul_469_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1297_nl))
      * $signed((ConvFiltWidth_else_mux1h_1298_nl)));
  assign z_out_1050_29_7 = readslicef_30_23_7((mul_469_nl));
  assign ConvFiltWidth_else_mux1h_1299_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[679:672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (MultLoop_io_read_w4_rsc_cse_sva[8799:8792]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1300_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[3]) , AccumDotWidth_or_145_cse , (fsm_output[5]) , (fsm_output[8])});
  assign mul_470_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1299_nl))
      * $signed((ConvFiltWidth_else_mux1h_1300_nl)));
  assign z_out_1051_29_7 = readslicef_30_23_7((mul_470_nl));
  assign ConvFiltWidth_else_mux1h_1301_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (w2_rsci_idat_mxwt[31:24]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (MultLoop_io_read_w4_rsc_cse_sva[8775:8768]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1302_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_73_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , AccumDotWidth_or_139_cse , AccumDotWidth_or_145_cse , (fsm_output[8])});
  assign mul_471_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1301_nl))
      * $signed((ConvFiltWidth_else_mux1h_1302_nl)));
  assign z_out_1052_29_7 = readslicef_30_23_7((mul_471_nl));
  assign ConvFiltWidth_else_mux1h_1303_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]), (MultLoop_io_read_w4_rsc_cse_sva[8823:8816]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_58_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_472_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1303_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_58_nl)));
  assign z_out_1053_29_7 = readslicef_30_23_7((mul_472_nl));
  assign ConvFiltWidth_else_mux1h_1304_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1063:1056]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]), (MultLoop_io_read_w4_rsc_cse_sva[8751:8744]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1305_nl = MUX1HOT_v_22_7_2((input_1_rsci_idat_mxwt[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[263:242]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_70_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_473_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1304_nl))
      * $signed((ConvFiltWidth_else_mux1h_1305_nl)));
  assign z_out_1054_29_7 = readslicef_30_23_7((mul_473_nl));
  assign ConvFiltWidth_else_mux1h_1306_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (w2_rsci_idat_mxwt[167:160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]), (MultLoop_io_read_w4_rsc_cse_sva[8767:8760]),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1307_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_72_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_474_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1306_nl))
      * $signed((ConvFiltWidth_else_mux1h_1307_nl)));
  assign z_out_1055_29_7 = readslicef_30_23_7((mul_474_nl));
  assign ConvFiltWidth_else_mux1h_1308_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[487:480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]),
      (MultLoop_io_read_w4_rsc_cse_sva[8831:8824]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1309_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_475_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1308_nl))
      * $signed((ConvFiltWidth_else_mux1h_1309_nl)));
  assign z_out_1056_29_7 = readslicef_30_23_7((mul_475_nl));
  assign ConvFiltWidth_else_mux1h_1310_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]), (MultLoop_io_read_w4_rsc_cse_sva[8791:8784]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_59_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_75_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_476_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1310_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_59_nl)));
  assign z_out_1057_29_7 = readslicef_30_23_7((mul_476_nl));
  assign ConvFiltWidth_else_mux1h_1311_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]),
      (w2_rsci_idat_mxwt[871:864]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]), (MultLoop_io_read_w4_rsc_cse_sva[8759:8752]),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1312_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[21:0]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_71_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_477_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1311_nl))
      * $signed((ConvFiltWidth_else_mux1h_1312_nl)));
  assign z_out_1058_29_7 = readslicef_30_23_7((mul_477_nl));
  assign ConvFiltWidth_else_mux1h_1313_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]),
      (w2_rsci_idat_mxwt[103:96]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_60_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[637:616]), fsm_output[1]);
  assign mul_478_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1313_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_60_nl)));
  assign z_out_1059_29_9 = readslicef_30_21_9((mul_478_nl));
  assign ConvFiltWidth_else_mux1h_1314_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6])});
  assign mul_479_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1314_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198])));
  assign z_out_1060_29_9 = readslicef_30_21_9((mul_479_nl));
  assign ConvFiltWidth_else_mux1h_1315_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6])});
  assign mul_480_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1315_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198])));
  assign z_out_1061_29_9 = readslicef_30_21_9((mul_480_nl));
  assign ConvFiltWidth_else_mux1h_1316_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (w2_rsci_idat_mxwt[359:352]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1317_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), {(fsm_output[2])
      , (fsm_output[1]) , AccumDotWidth_or_38_cse , (fsm_output[7])});
  assign mul_481_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1316_nl))
      * $signed((ConvFiltWidth_else_mux1h_1317_nl)));
  assign z_out_1062_29_9 = readslicef_30_21_9((mul_481_nl));
  assign ConvFiltWidth_else_mux1h_1318_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[167:160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1319_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[725:704]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[219:198]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[747:726]), {(fsm_output[1])
      , (fsm_output[2]) , AccumDotWidth_or_38_cse , (fsm_output[7])});
  assign mul_482_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1318_nl))
      * $signed((ConvFiltWidth_else_mux1h_1319_nl)));
  assign z_out_1063_29_9 = readslicef_30_21_9((mul_482_nl));
  assign ConvFiltWidth_else_mux1h_1320_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[471:464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]), (MultLoop_io_read_w4_rsc_cse_sva[5727:5720]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1321_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1081_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_483_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1320_nl))
      * $signed((ConvFiltWidth_else_mux1h_1321_nl)));
  assign z_out_1064_29_7 = readslicef_30_23_7((mul_483_nl));
  assign ConvFiltWidth_else_mux1h_1322_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]),
      (w2_rsci_idat_mxwt[1135:1128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1323_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]), {(fsm_output[2])
      , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , AccumDotWidth_or_140_cse});
  assign mul_484_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1322_nl))
      * $signed((ConvFiltWidth_else_mux1h_1323_nl)));
  assign z_out_1065_29_9 = readslicef_30_21_9((mul_484_nl));
  assign ConvFiltWidth_else_mux1h_1324_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (w2_rsci_idat_mxwt[295:288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_61_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[703:682]), fsm_output[1]);
  assign mul_485_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1324_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_61_nl)));
  assign z_out_1066_29_9 = readslicef_30_21_9((mul_485_nl));
  assign ConvFiltWidth_else_mux1h_1325_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (w2_rsci_idat_mxwt[999:992]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_62_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[835:814]),
      (input_1_rsci_idat_mxwt[1011:990]), fsm_output[1]);
  assign mul_486_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1325_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_62_nl)));
  assign z_out_1067_29_9 = readslicef_30_21_9((mul_486_nl));
  assign ConvFiltWidth_else_mux1h_1326_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]),
      (w2_rsci_idat_mxwt[175:168]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[743:736]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]), (MultLoop_io_read_w4_rsc_cse_sva[8743:8736]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1327_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_69_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5])
      , (fsm_output[8])});
  assign mul_487_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1326_nl))
      * $signed((ConvFiltWidth_else_mux1h_1327_nl)));
  assign z_out_1068_29_7 = readslicef_30_23_7((mul_487_nl));
  assign ConvFiltWidth_else_mux1h_1328_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (w2_rsci_idat_mxwt[879:872]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (MultLoop_io_read_w4_rsc_cse_sva[8735:8728]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1329_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_68_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_488_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1328_nl))
      * $signed((ConvFiltWidth_else_mux1h_1329_nl)));
  assign z_out_1069_29_7 = readslicef_30_23_7((mul_488_nl));
  assign ConvFiltWidth_else_mux1h_1330_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (w2_rsci_idat_mxwt[751:744]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]), (MultLoop_io_read_w4_rsc_cse_sva[8727:8720]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1331_nl = MUX1HOT_v_22_6_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_152_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_489_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1330_nl))
      * $signed((ConvFiltWidth_else_mux1h_1331_nl)));
  assign z_out_1070_29_7 = readslicef_30_23_7((mul_489_nl));
  assign ConvFiltWidth_else_mux1h_1332_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[367:360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (MultLoop_io_read_w4_rsc_cse_sva[8719:8712]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , AccumDotWidth_or_152_cse , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1333_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[5]) , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_490_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1332_nl))
      * $signed((ConvFiltWidth_else_mux1h_1333_nl)));
  assign z_out_1071_29_7 = readslicef_30_23_7((mul_490_nl));
  assign ConvFiltWidth_else_mux1h_1334_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]),
      (w2_rsci_idat_mxwt[687:680]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (MultLoop_io_read_w4_rsc_cse_sva[8711:8704]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1335_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_65_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_491_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1334_nl))
      * $signed((ConvFiltWidth_else_mux1h_1335_nl)));
  assign z_out_1072_29_7 = readslicef_30_23_7((mul_491_nl));
  assign ConvFiltWidth_else_mux1h_1336_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[103:96]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]), (MultLoop_io_read_w4_rsc_cse_sva[8663:8656]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1337_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , MultLoop_or_46_cse , (fsm_output[5]) ,
      (fsm_output[7]) , (fsm_output[8])});
  assign mul_492_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1336_nl))
      * $signed((ConvFiltWidth_else_mux1h_1337_nl)));
  assign z_out_1073_29_7 = readslicef_30_23_7((mul_492_nl));
  assign ConvFiltWidth_else_mux1h_1338_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[807:800]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1479:1472]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[135:128]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]),
      (MultLoop_io_read_w4_rsc_cse_sva[8671:8664]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1339_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[1011:990]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_493_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1338_nl))
      * $signed((ConvFiltWidth_else_mux1h_1339_nl)));
  assign z_out_1074_29_7 = readslicef_30_23_7((mul_493_nl));
  assign ConvFiltWidth_else_mux1h_1340_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]), (MultLoop_io_read_w4_rsc_cse_sva[8679:8672]),
      {(fsm_output[1]) , AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1341_nl = MUX1HOT_v_22_7_2((input_1_rsci_idat_mxwt[1033:1012]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[857:836]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[43:22]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_152_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_494_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1340_nl))
      * $signed((ConvFiltWidth_else_mux1h_1341_nl)));
  assign z_out_1075_29_7 = readslicef_30_23_7((mul_494_nl));
  assign ConvFiltWidth_else_mux1h_1342_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]),
      (w2_rsci_idat_mxwt[295:288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]),
      (MultLoop_io_read_w4_rsc_cse_sva[8703:8696]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1343_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_495_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1342_nl))
      * $signed((ConvFiltWidth_else_mux1h_1343_nl)));
  assign z_out_1076_29_7 = readslicef_30_23_7((mul_495_nl));
  assign ConvFiltWidth_else_mux1h_1344_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]),
      (w2_rsci_idat_mxwt[711:704]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1031:1024]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[471:464]),
      (MultLoop_io_read_w4_rsc_cse_sva[8695:8688]), {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1345_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_787_cse , (fsm_output[8])});
  assign mul_496_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1344_nl))
      * $signed((ConvFiltWidth_else_mux1h_1345_nl)));
  assign z_out_1077_29_7 = readslicef_30_23_7((mul_496_nl));
  assign ConvFiltWidth_else_mux1h_1346_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (w2_rsci_idat_mxwt[303:296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[351:344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (MultLoop_io_read_w4_rsc_cse_sva[4567:4560]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1347_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_59_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_497_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1346_nl))
      * $signed((ConvFiltWidth_else_mux1h_1347_nl)));
  assign z_out_1078_29_7 = readslicef_30_23_7((mul_497_nl));
  assign ConvFiltWidth_else_mux1h_1348_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (w2_rsci_idat_mxwt[679:672]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[735:728]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (MultLoop_io_read_w4_rsc_cse_sva[4607:4600]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1349_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[967:946]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[65:44]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_752_cse , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_498_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1348_nl))
      * $signed((ConvFiltWidth_else_mux1h_1349_nl)));
  assign z_out_1079_29_7 = readslicef_30_23_7((mul_498_nl));
  assign ConvFiltWidth_else_mux1h_1350_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[367:360]),
      (w2_rsci_idat_mxwt[767:760]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]), (MultLoop_io_read_w4_rsc_cse_sva[4591:4584]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1351_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[857:836]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_499_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1350_nl))
      * $signed((ConvFiltWidth_else_mux1h_1351_nl)));
  assign z_out_1080_29_7 = readslicef_30_23_7((mul_499_nl));
  assign ConvFiltWidth_else_mux1h_1352_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]),
      (w2_rsci_idat_mxwt[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1327:1320]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]),
      (MultLoop_io_read_w4_rsc_cse_sva[8687:8680]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1353_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_871_cse , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_500_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1352_nl))
      * $signed((ConvFiltWidth_else_mux1h_1353_nl)));
  assign z_out_1081_29_7 = readslicef_30_23_7((mul_500_nl));
  assign ConvFiltWidth_else_mux1h_1354_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]),
      (w2_rsci_idat_mxwt[711:704]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (MultLoop_io_read_w4_rsc_cse_sva[7879:7872]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1355_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}), {ConvFiltWidth_else_or_871_cse
      , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_501_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1354_nl))
      * $signed((ConvFiltWidth_else_mux1h_1355_nl)));
  assign z_out_1082_29_7 = readslicef_30_23_7((mul_501_nl));
  assign ConvFiltWidth_else_mux1h_1356_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[527:520]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1311:1304]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (MultLoop_io_read_w4_rsc_cse_sva[7871:7864]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1357_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]), ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}),
      {(fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_502_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1356_nl))
      * $signed((ConvFiltWidth_else_mux1h_1357_nl)));
  assign z_out_1083_29_7 = readslicef_30_23_7((mul_502_nl));
  assign ConvFiltWidth_else_mux1h_1358_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]), (w2_rsci_idat_mxwt[911:904]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]),
      (MultLoop_io_read_w4_rsc_cse_sva[7831:7824]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1359_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_503_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1358_nl))
      * $signed((ConvFiltWidth_else_mux1h_1359_nl)));
  assign z_out_1084_29_7 = readslicef_30_23_7((mul_503_nl));
  assign ConvFiltWidth_else_mux1h_1360_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]),
      (MultLoop_io_read_w4_rsc_cse_sva[7823:7816]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_63_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_504_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1360_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_63_nl)));
  assign z_out_1085_29_7 = readslicef_30_23_7((mul_504_nl));
  assign ConvFiltWidth_else_mux1h_1361_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]), (w2_rsci_idat_mxwt[719:712]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1303:1296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (MultLoop_io_read_w4_rsc_cse_sva[7887:7880]), {(fsm_output[6]) , (fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1362_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}), {ConvFiltWidth_else_or_871_cse
      , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_505_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1361_nl))
      * $signed((ConvFiltWidth_else_mux1h_1362_nl)));
  assign z_out_1086_29_7 = readslicef_30_23_7((mul_505_nl));
  assign ConvFiltWidth_else_mux1h_1363_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]),
      (MultLoop_io_read_w4_rsc_cse_sva[7847:7840]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_64_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}), fsm_output[8]);
  assign mul_506_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1363_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_64_nl)));
  assign z_out_1087_29_7 = readslicef_30_23_7((mul_506_nl));
  assign ConvFiltWidth_else_mux1h_1364_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[383:376]),
      (w2_rsci_idat_mxwt[383:376]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1295:1288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (MultLoop_io_read_w4_rsc_cse_sva[7839:7832]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1365_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_29_cse , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_507_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1364_nl))
      * $signed((ConvFiltWidth_else_mux1h_1365_nl)));
  assign z_out_1088_29_7 = readslicef_30_23_7((mul_507_nl));
  assign ConvFiltWidth_else_mux1h_1366_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[375:368]),
      (w2_rsci_idat_mxwt[575:568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1335:1328]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]),
      (MultLoop_io_read_w4_rsc_cse_sva[7895:7888]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1367_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {AccumDotWidth_or_29_cse , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_508_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1366_nl))
      * $signed((ConvFiltWidth_else_mux1h_1367_nl)));
  assign z_out_1089_29_7 = readslicef_30_23_7((mul_508_nl));
  assign ConvFiltWidth_else_mux1h_1368_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (w2_rsci_idat_mxwt[519:512]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1319:1312]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]),
      (MultLoop_io_read_w4_rsc_cse_sva[7863:7856]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1369_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}), {ConvFiltWidth_else_or_871_cse
      , (fsm_output[1]) , MultLoop_or_46_cse , (fsm_output[8])});
  assign mul_509_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1368_nl))
      * $signed((ConvFiltWidth_else_mux1h_1369_nl)));
  assign z_out_1090_29_7 = readslicef_30_23_7((mul_509_nl));
  assign ConvFiltWidth_else_mux1h_1370_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[359:352]),
      (w2_rsci_idat_mxwt[327:320]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1287:1280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]), (MultLoop_io_read_w4_rsc_cse_sva[4559:4552]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1371_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_58_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_510_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1370_nl))
      * $signed((ConvFiltWidth_else_mux1h_1371_nl)));
  assign z_out_1091_29_7 = readslicef_30_23_7((mul_510_nl));
  assign ConvFiltWidth_else_mux1h_1372_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[671:664]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[727:720]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]), (MultLoop_io_read_w4_rsc_cse_sva[4583:4576]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1373_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_87_cse , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_511_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1372_nl))
      * $signed((ConvFiltWidth_else_mux1h_1373_nl)));
  assign z_out_1092_29_7 = readslicef_30_23_7((mul_511_nl));
  assign ConvFiltWidth_else_mux1h_1374_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]),
      (w2_rsci_idat_mxwt[111:104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]),
      (MultLoop_io_read_w4_rsc_cse_sva[7855:7848]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1375_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (input_1_rsci_idat_mxwt[571:550]), ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_512_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1374_nl))
      * $signed((ConvFiltWidth_else_mux1h_1375_nl)));
  assign z_out_1093_29_7 = readslicef_30_23_7((mul_512_nl));
  assign ConvFiltWidth_else_mux1h_1376_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1055:1048]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (MultLoop_io_read_w4_rsc_cse_sva[7903:7896]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1377_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[1]) , MultLoop_or_87_cse , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_513_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1376_nl))
      * $signed((ConvFiltWidth_else_mux1h_1377_nl)));
  assign z_out_1094_29_7 = readslicef_30_23_7((mul_513_nl));
  assign ConvFiltWidth_else_mux1h_1378_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]),
      (w2_rsci_idat_mxwt[1023:1016]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1623:1616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      (MultLoop_io_read_w4_rsc_cse_sva[4575:4568]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_or_1166_nl = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1379_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , (ConvFiltWidth_else_or_1166_nl) , (fsm_output[8])});
  assign mul_514_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1378_nl))
      * $signed((ConvFiltWidth_else_mux1h_1379_nl)));
  assign z_out_1095_29_7 = readslicef_30_23_7((mul_514_nl));
  assign ConvFiltWidth_else_mux1h_1380_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[687:680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (MultLoop_io_read_w4_rsc_cse_sva[5575:5568]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1381_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_515_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1380_nl))
      * $signed((ConvFiltWidth_else_mux1h_1381_nl)));
  assign z_out_1096_29_7 = readslicef_30_23_7((mul_515_nl));
  assign ConvFiltWidth_else_mux1h_1382_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[879:872]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[719:712]),
      (MultLoop_io_read_w4_rsc_cse_sva[6679:6672]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse , (fsm_output[6])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1383_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_87_cse , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_516_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1382_nl))
      * $signed((ConvFiltWidth_else_mux1h_1383_nl)));
  assign z_out_1097_29_7 = readslicef_30_23_7((mul_516_nl));
  assign ConvFiltWidth_else_or_1171_cse = (fsm_output[3]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1384_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      (w2_rsci_idat_mxwt[495:488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[959:952]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]), (MultLoop_io_read_w4_rsc_cse_sva[6639:6632]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1385_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_1171_cse , (fsm_output[8])});
  assign mul_517_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1384_nl))
      * $signed((ConvFiltWidth_else_mux1h_1385_nl)));
  assign z_out_1098_29_7 = readslicef_30_23_7((mul_517_nl));
  assign ConvFiltWidth_else_mux1h_1386_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[159:152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (MultLoop_io_read_w4_rsc_cse_sva[6767:6760]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1387_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_17_cse , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_518_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1386_nl))
      * $signed((ConvFiltWidth_else_mux1h_1387_nl)));
  assign z_out_1099_29_7 = readslicef_30_23_7((mul_518_nl));
  assign ConvFiltWidth_else_mux1h_1388_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[303:296]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[711:704]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]), (MultLoop_io_read_w4_rsc_cse_sva[6671:6664]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1389_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[461:440]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_519_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1388_nl))
      * $signed((ConvFiltWidth_else_mux1h_1389_nl)));
  assign z_out_1100_29_7 = readslicef_30_23_7((mul_519_nl));
  assign ConvFiltWidth_else_mux1h_1390_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1007:1000]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (MultLoop_io_read_w4_rsc_cse_sva[6759:6752]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1391_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , ConvFiltWidth_else_or_1171_cse , (fsm_output[8])});
  assign mul_520_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1390_nl))
      * $signed((ConvFiltWidth_else_mux1h_1391_nl)));
  assign z_out_1101_29_7 = readslicef_30_23_7((mul_520_nl));
  assign ConvFiltWidth_else_mux1h_1392_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]),
      (MultLoop_io_read_w4_rsc_cse_sva[6631:6624]), {(fsm_output[3]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_65_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_521_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1392_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_65_nl)));
  assign z_out_1102_29_7 = readslicef_30_23_7((mul_521_nl));
  assign ConvFiltWidth_else_mux1h_1393_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[863:856]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (MultLoop_io_read_w4_rsc_cse_sva[6751:6744]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1394_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[417:396]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_6_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_522_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1393_nl))
      * $signed((ConvFiltWidth_else_mux1h_1394_nl)));
  assign z_out_1103_29_7 = readslicef_30_23_7((mul_522_nl));
  assign ConvFiltWidth_else_mux1h_1395_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[167:160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]),
      (MultLoop_io_read_w4_rsc_cse_sva[6655:6648]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1396_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[593:572]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[373:352]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_17_cse , (fsm_output[8])});
  assign mul_523_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1395_nl))
      * $signed((ConvFiltWidth_else_mux1h_1396_nl)));
  assign z_out_1104_29_7 = readslicef_30_23_7((mul_523_nl));
  assign ConvFiltWidth_else_mux1h_1397_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]),
      (w2_rsci_idat_mxwt[319:312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (MultLoop_io_read_w4_rsc_cse_sva[6623:6616]),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1398_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_60_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_524_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1397_nl))
      * $signed((ConvFiltWidth_else_mux1h_1398_nl)));
  assign z_out_1105_29_7 = readslicef_30_23_7((mul_524_nl));
  assign ConvFiltWidth_else_mux1h_1399_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      (w2_rsci_idat_mxwt[831:824]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[503:496]),
      (MultLoop_io_read_w4_rsc_cse_sva[6647:6640]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1400_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_987_cse , (fsm_output[1]) , AccumDotWidth_or_139_cse
      , (fsm_output[8])});
  assign mul_525_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1399_nl))
      * $signed((ConvFiltWidth_else_mux1h_1400_nl)));
  assign z_out_1106_29_7 = readslicef_30_23_7((mul_525_nl));
  assign ConvFiltWidth_else_mux1h_1401_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[511:504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1487:1480]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[463:456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]), (MultLoop_io_read_w4_rsc_cse_sva[4543:4536]),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1402_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_56_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_526_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1401_nl))
      * $signed((ConvFiltWidth_else_mux1h_1402_nl)));
  assign z_out_1107_29_7 = readslicef_30_23_7((mul_526_nl));
  assign ConvFiltWidth_else_or_1183_cse = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[7]);
  assign ConvFiltWidth_else_mux1h_1403_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]),
      (w2_rsci_idat_mxwt[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1687:1680]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (MultLoop_io_read_w4_rsc_cse_sva[4119:4112]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1404_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_3_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1183_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign mul_527_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1403_nl))
      * $signed((ConvFiltWidth_else_mux1h_1404_nl)));
  assign z_out_1108_29_7 = readslicef_30_23_7((mul_527_nl));
  assign ConvFiltWidth_else_mux1h_1405_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]),
      (w2_rsci_idat_mxwt[1023:1016]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]),
      (MultLoop_io_read_w4_rsc_cse_sva[4551:4544]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1406_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[945:924]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_57_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_528_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1405_nl))
      * $signed((ConvFiltWidth_else_mux1h_1406_nl)));
  assign z_out_1109_29_7 = readslicef_30_23_7((mul_528_nl));
  assign ConvFiltWidth_else_mux1h_1407_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (w2_rsci_idat_mxwt[79:72]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]), (MultLoop_io_read_w4_rsc_cse_sva[4855:4848]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1408_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_26_cse , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_529_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1407_nl))
      * $signed((ConvFiltWidth_else_mux1h_1408_nl)));
  assign z_out_1110_29_7 = readslicef_30_23_7((mul_529_nl));
  assign ConvFiltWidth_else_mux1h_1409_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[279:272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]),
      (MultLoop_io_read_w4_rsc_cse_sva[4847:4840]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1410_nl = MUX1HOT_v_22_6_2((input_1_rsci_idat_mxwt[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_94_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_29_cse , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_530_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1409_nl))
      * $signed((ConvFiltWidth_else_mux1h_1410_nl)));
  assign z_out_1111_29_7 = readslicef_30_23_7((mul_530_nl));
  assign ConvFiltWidth_else_mux1h_1411_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]),
      (w2_rsci_idat_mxwt[343:336]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (MultLoop_io_read_w4_rsc_cse_sva[4839:4832]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1412_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[791:770]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {AccumDotWidth_or_26_cse , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[8])});
  assign mul_531_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1411_nl))
      * $signed((ConvFiltWidth_else_mux1h_1412_nl)));
  assign z_out_1112_29_7 = readslicef_30_23_7((mul_531_nl));
  assign ConvFiltWidth_else_mux1h_1413_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]),
      (w2_rsci_idat_mxwt[783:776]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]),
      (MultLoop_io_read_w4_rsc_cse_sva[4775:4768]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1414_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[1011:990]), ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}),
      {AccumDotWidth_or_26_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_532_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1413_nl))
      * $signed((ConvFiltWidth_else_mux1h_1414_nl)));
  assign z_out_1113_29_7 = readslicef_30_23_7((mul_532_nl));
  assign ConvFiltWidth_else_mux1h_1415_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]),
      (w2_rsci_idat_mxwt[271:264]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (MultLoop_io_read_w4_rsc_cse_sva[4783:4776]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1416_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[769:748]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_533_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1415_nl))
      * $signed((ConvFiltWidth_else_mux1h_1416_nl)));
  assign z_out_1114_29_7 = readslicef_30_23_7((mul_533_nl));
  assign ConvFiltWidth_else_mux1h_1417_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]),
      (w2_rsci_idat_mxwt[663:656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (MultLoop_io_read_w4_rsc_cse_sva[4791:4784]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1418_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1011:990]), ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_534_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1417_nl))
      * $signed((ConvFiltWidth_else_mux1h_1418_nl)));
  assign z_out_1115_29_7 = readslicef_30_23_7((mul_534_nl));
  assign ConvFiltWidth_else_mux1h_1419_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]),
      (w2_rsci_idat_mxwt[151:144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[575:568]),
      (MultLoop_io_read_w4_rsc_cse_sva[4799:4792]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1420_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[725:704]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[527:506]), ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[6]) , (fsm_output[7]) ,
      (fsm_output[8])});
  assign mul_535_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1419_nl))
      * $signed((ConvFiltWidth_else_mux1h_1420_nl)));
  assign z_out_1116_29_7 = readslicef_30_23_7((mul_535_nl));
  assign ConvFiltWidth_else_mux1h_1421_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]),
      (w2_rsci_idat_mxwt[655:648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[519:512]),
      (MultLoop_io_read_w4_rsc_cse_sva[4807:4800]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1422_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[967:946]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}), {MultLoop_or_17_cse , (fsm_output[1])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_536_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1421_nl))
      * $signed((ConvFiltWidth_else_mux1h_1422_nl)));
  assign z_out_1117_29_7 = readslicef_30_23_7((mul_536_nl));
  assign ConvFiltWidth_else_mux1h_1423_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (w2_rsci_idat_mxwt[87:80]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1175:1168]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]), (MultLoop_io_read_w4_rsc_cse_sva[4815:4808]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , operator_22_4_true_AC_TRN_AC_WRAP_or_8_cse
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1424_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[703:682]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1033:1012]), ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_537_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1423_nl))
      * $signed((ConvFiltWidth_else_mux1h_1424_nl)));
  assign z_out_1118_29_7 = readslicef_30_23_7((mul_537_nl));
  assign ConvFiltWidth_else_mux1h_1425_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]),
      (w2_rsci_idat_mxwt[727:720]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]),
      (MultLoop_io_read_w4_rsc_cse_sva[4823:4816]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1426_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[989:968]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {MultLoop_or_17_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_538_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1425_nl))
      * $signed((ConvFiltWidth_else_mux1h_1426_nl)));
  assign z_out_1119_29_7 = readslicef_30_23_7((mul_538_nl));
  assign ConvFiltWidth_else_mux1h_1427_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1183:1176]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]), (MultLoop_io_read_w4_rsc_cse_sva[2583:2576]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1428_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_539_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1427_nl))
      * $signed((ConvFiltWidth_else_mux1h_1428_nl)));
  assign z_out_1120_29_7 = readslicef_30_23_7((mul_539_nl));
  assign ConvFiltWidth_else_mux1h_1429_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]),
      (w2_rsci_idat_mxwt[855:848]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[919:912]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]),
      (MultLoop_io_read_w4_rsc_cse_sva[2535:2528]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1430_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[285:264]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[725:704]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_540_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1429_nl))
      * $signed((ConvFiltWidth_else_mux1h_1430_nl)));
  assign z_out_1121_29_7 = readslicef_30_23_7((mul_540_nl));
  assign ConvFiltWidth_else_mux1h_1431_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[127:120]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[751:744]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[167:160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[191:184]),
      (MultLoop_io_read_w4_rsc_cse_sva[2543:2536]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1432_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_541_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1431_nl))
      * $signed((ConvFiltWidth_else_mux1h_1432_nl)));
  assign z_out_1122_29_7 = readslicef_30_23_7((mul_541_nl));
  assign ConvFiltWidth_else_mux1h_1433_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[759:752]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[183:176]), (MultLoop_io_read_w4_rsc_cse_sva[4831:4824]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1434_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_542_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1433_nl))
      * $signed((ConvFiltWidth_else_mux1h_1434_nl)));
  assign z_out_1123_29_7 = readslicef_30_23_7((mul_542_nl));
  assign ConvFiltWidth_else_mux1h_1435_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]),
      (MultLoop_io_read_w4_rsc_cse_sva[2575:2568]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_66_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_543_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1435_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_66_nl)));
  assign z_out_1124_29_7 = readslicef_30_23_7((mul_543_nl));
  assign ConvFiltWidth_else_mux1h_1436_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]),
      (MultLoop_io_read_w4_rsc_cse_sva[2663:2656]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_67_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_544_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1436_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_67_nl)));
  assign z_out_1125_29_7 = readslicef_30_23_7((mul_544_nl));
  assign ConvFiltWidth_else_mux1h_1437_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (w2_rsci_idat_mxwt[447:440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1095:1088]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[159:152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]),
      (MultLoop_io_read_w4_rsc_cse_sva[2551:2544]), {(fsm_output[2]) , (fsm_output[1])
      , AccumDotWidth_or_157_cse , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1438_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse
      , (fsm_output[8])});
  assign mul_545_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1437_nl))
      * $signed((ConvFiltWidth_else_mux1h_1438_nl)));
  assign z_out_1126_29_7 = readslicef_30_23_7((mul_545_nl));
  assign ConvFiltWidth_else_mux1h_1439_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1191:1184]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (MultLoop_io_read_w4_rsc_cse_sva[2559:2552]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1440_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_1081_cse , (fsm_output[8])});
  assign mul_546_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1439_nl))
      * $signed((ConvFiltWidth_else_mux1h_1440_nl)));
  assign z_out_1127_29_7 = readslicef_30_23_7((mul_546_nl));
  assign ConvFiltWidth_else_mux1h_1441_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]),
      (w2_rsci_idat_mxwt[895:888]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[935:928]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1695:1688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]), (MultLoop_io_read_w4_rsc_cse_sva[2679:2672]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1442_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1183_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])
      , (fsm_output[8])});
  assign mul_547_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1441_nl))
      * $signed((ConvFiltWidth_else_mux1h_1442_nl)));
  assign z_out_1128_29_7 = readslicef_30_23_7((mul_547_nl));
  assign ConvFiltWidth_else_mux1h_1443_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[511:504]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[943:936]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[767:760]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[175:168]), (MultLoop_io_read_w4_rsc_cse_sva[2671:2664]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1444_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse
      , (fsm_output[8])});
  assign mul_548_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1443_nl))
      * $signed((ConvFiltWidth_else_mux1h_1444_nl)));
  assign z_out_1129_29_7 = readslicef_30_23_7((mul_548_nl));
  assign ConvFiltWidth_else_mux1h_1445_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]), (w2_rsci_idat_mxwt[447:440]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1071:1064]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]),
      (MultLoop_io_read_w4_rsc_cse_sva[4111:4104]), {(fsm_output[2]) , (fsm_output[3])
      , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1446_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[87:66]), (input_1_rsci_idat_mxwt[747:726]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_2_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[1]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_549_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1445_nl))
      * $signed((ConvFiltWidth_else_mux1h_1446_nl)));
  assign z_out_1130_29_7 = readslicef_30_23_7((mul_549_nl));
  assign ConvFiltWidth_else_mux1h_1447_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[327:320]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1047:1040]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1495:1488]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[839:832]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]), (MultLoop_io_read_w4_rsc_cse_sva[4599:4592]),
      {(fsm_output[1]) , MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1448_nl = MUX1HOT_v_22_5_2((input_1_rsci_idat_mxwt[791:770]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[395:374]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_550_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1447_nl))
      * $signed((ConvFiltWidth_else_mux1h_1448_nl)));
  assign z_out_1131_29_7 = readslicef_30_23_7((mul_550_nl));
  assign ConvFiltWidth_else_mux1h_1449_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (w2_rsci_idat_mxwt[639:632]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[5])});
  assign ConvFiltWidth_else_mux1h_1450_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[813:792]),
      (input_1_rsci_idat_mxwt[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      {(fsm_output[2]) , (fsm_output[1]) , AccumDotWidth_or_139_cse});
  assign mul_551_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1449_nl))
      * $signed((ConvFiltWidth_else_mux1h_1450_nl)));
  assign z_out_1132_29_9 = readslicef_30_21_9((mul_551_nl));
  assign ConvFiltWidth_else_mux1h_1451_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[319:312]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[903:896]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[151:144]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1671:1664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1519:1512]),
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1452_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse});
  assign mul_552_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1451_nl))
      * $signed((ConvFiltWidth_else_mux1h_1452_nl)));
  assign z_out_1133_29_9 = readslicef_30_21_9((mul_552_nl));
  assign ConvFiltWidth_else_mux1h_1453_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[639:632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1103:1096]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[143:136]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[951:944]), {(fsm_output[1]) , AccumDotWidth_or_157_cse
      , (fsm_output[5]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1454_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse});
  assign mul_553_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1453_nl))
      * $signed((ConvFiltWidth_else_mux1h_1454_nl)));
  assign z_out_1134_29_9 = readslicef_30_21_9((mul_553_nl));
  assign ConvFiltWidth_else_mux1h_1455_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]),
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign mul_554_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1455_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528])));
  assign z_out_1135_29_9 = readslicef_30_21_9((mul_554_nl));
  assign ConvFiltWidth_else_mux1h_1456_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[295:288]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])});
  assign mul_555_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1456_nl))
      * $signed((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550])));
  assign z_out_1136_29_9 = readslicef_30_21_9((mul_555_nl));
  assign ConvFiltWidth_else_mux1h_1457_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[967:960]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1679:1672]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1527:1520]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1458_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[1011:990]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[153:132]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), {(fsm_output[1])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse});
  assign mul_556_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1457_nl))
      * $signed((ConvFiltWidth_else_mux1h_1458_nl)));
  assign z_out_1137_29_9 = readslicef_30_21_9((mul_556_nl));
  assign ConvFiltWidth_else_mux1h_1459_nl = MUX1HOT_v_8_4_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      (w2_rsci_idat_mxwt[663:656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), {AccumDotWidth_or_25_cse
      , (fsm_output[1]) , (fsm_output[5]) , (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1460_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , AccumDotWidth_or_152_cse});
  assign mul_557_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1459_nl))
      * $signed((ConvFiltWidth_else_mux1h_1460_nl)));
  assign z_out_1138_29_9 = readslicef_30_21_9((mul_557_nl));
  assign ConvFiltWidth_else_mux1h_1461_nl = MUX1HOT_v_8_3_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      {(fsm_output[2]) , AccumDotWidth_or_157_cse , (fsm_output[4])});
  assign ConvFiltWidth_else_mux1h_1462_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[791:770]),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[3]) , (fsm_output[6])});
  assign mul_558_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1461_nl))
      * $signed((ConvFiltWidth_else_mux1h_1462_nl)));
  assign z_out_1139_29_9 = readslicef_30_21_9((mul_558_nl));
  assign ConvFiltWidth_else_mux1h_1463_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      (w2_rsci_idat_mxwt[191:184]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[927:920]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1464_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[549:528]),
      (input_1_rsci_idat_mxwt[593:572]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[131:110]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]), {(fsm_output[2])
      , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse});
  assign mul_559_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1463_nl))
      * $signed((ConvFiltWidth_else_mux1h_1464_nl)));
  assign z_out_1140_29_9 = readslicef_30_21_9((mul_559_nl));
  assign ConvFiltWidth_else_mux1h_1465_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[63:56]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1607:1600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]),
      {(fsm_output[1]) , AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1466_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      {(fsm_output[1]) , (fsm_output[2]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse});
  assign mul_560_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1465_nl))
      * $signed((ConvFiltWidth_else_mux1h_1466_nl)));
  assign z_out_1141_29_9 = readslicef_30_21_9((mul_560_nl));
  assign ConvFiltWidth_else_mux1h_1467_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]),
      (w2_rsci_idat_mxwt[703:696]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1631:1624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[479:472]),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_1_cse , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])});
  assign ConvFiltWidth_else_mux1h_1468_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (input_1_rsci_idat_mxwt[901:880]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      {(fsm_output[2]) , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse});
  assign mul_561_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1467_nl))
      * $signed((ConvFiltWidth_else_mux1h_1468_nl)));
  assign z_out_1142_29_9 = readslicef_30_21_9((mul_561_nl));
  assign ConvFiltWidth_else_mux1h_1469_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]),
      (w2_rsci_idat_mxwt[127:120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1615:1608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1423:1416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1079:1072]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[495:488]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1470_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[637:616]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_861_cse});
  assign mul_562_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1469_nl))
      * $signed((ConvFiltWidth_else_mux1h_1470_nl)));
  assign z_out_1143_29_9 = readslicef_30_21_9((mul_562_nl));
  assign ConvFiltWidth_else_mux1h_1471_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]),
      (w2_rsci_idat_mxwt[255:248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[511:504]),
      {MultLoop_or_87_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[6]) ,
      (fsm_output[7])});
  assign ConvFiltWidth_else_mux1h_1472_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[901:880]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[505:484]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]), {(fsm_output[2])
      , (fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse
      , (fsm_output[5])});
  assign mul_563_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1471_nl))
      * $signed((ConvFiltWidth_else_mux1h_1472_nl)));
  assign z_out_1144_29_9 = readslicef_30_21_9((mul_563_nl));
  assign ConvFiltWidth_else_mux1h_1473_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[807:800]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[631:624]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[639:632]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[63:56]),
      (MultLoop_io_read_w4_rsc_cse_sva[3743:3736]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1474_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[879:858]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_849_cse , (fsm_output[8])});
  assign mul_564_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1473_nl))
      * $signed((ConvFiltWidth_else_mux1h_1474_nl)));
  assign z_out_1145_29_7 = readslicef_30_23_7((mul_564_nl));
  assign ConvFiltWidth_else_mux1h_1475_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]),
      (w2_rsci_idat_mxwt[143:136]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1167:1160]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[591:584]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[127:120]),
      (MultLoop_io_read_w4_rsc_cse_sva[3703:3696]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1476_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (input_1_rsci_idat_mxwt[593:572]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_565_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1475_nl))
      * $signed((ConvFiltWidth_else_mux1h_1476_nl)));
  assign z_out_1146_29_7 = readslicef_30_23_7((mul_565_nl));
  assign ConvFiltWidth_else_mux1h_1477_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (MultLoop_io_read_w4_rsc_cse_sva[3751:3744]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1478_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[901:880]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , (AccumDotWidth_acc_1871_itm[20:0])}), {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse
      , (fsm_output[7]) , (fsm_output[8])});
  assign mul_566_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1477_nl))
      * $signed((ConvFiltWidth_else_mux1h_1478_nl)));
  assign z_out_1147_29_7 = readslicef_30_23_7((mul_566_nl));
  assign ConvFiltWidth_else_mux1h_1479_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[623:616]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[47:40]), (MultLoop_io_read_w4_rsc_cse_sva[3759:3752]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_68_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}), fsm_output[8]);
  assign mul_567_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1479_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_68_nl)));
  assign z_out_1148_29_7 = readslicef_30_23_7((mul_567_nl));
  assign ConvFiltWidth_else_mux1h_1480_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[55:48]), (MultLoop_io_read_w4_rsc_cse_sva[3767:3760]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_69_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}), fsm_output[8]);
  assign mul_568_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1480_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_69_nl)));
  assign z_out_1149_29_7 = readslicef_30_23_7((mul_568_nl));
  assign ConvFiltWidth_else_mux1h_1481_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1199:1192]),
      (w2_rsci_idat_mxwt[247:240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (MultLoop_io_read_w4_rsc_cse_sva[3775:3768]), {(fsm_output[3]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1482_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}), {MultLoop_or_46_cse , (fsm_output[1])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_569_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1481_nl))
      * $signed((ConvFiltWidth_else_mux1h_1482_nl)));
  assign z_out_1150_29_7 = readslicef_30_23_7((mul_569_nl));
  assign ConvFiltWidth_else_mux1h_1483_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[423:416]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1215:1208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[23:16]), (MultLoop_io_read_w4_rsc_cse_sva[3735:3728]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1484_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[681:660]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse , (fsm_output[8])});
  assign mul_570_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1483_nl))
      * $signed((ConvFiltWidth_else_mux1h_1484_nl)));
  assign z_out_1151_29_7 = readslicef_30_23_7((mul_570_nl));
  assign ConvFiltWidth_else_mux1h_1485_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[231:224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1159:1152]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[615:608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[455:448]),
      (MultLoop_io_read_w4_rsc_cse_sva[3711:3704]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1486_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_17_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_571_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1485_nl))
      * $signed((ConvFiltWidth_else_mux1h_1486_nl)));
  assign z_out_1152_29_7 = readslicef_30_23_7((mul_571_nl));
  assign ConvFiltWidth_else_mux1h_1487_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[655:648]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[15:8]), (MultLoop_io_read_w4_rsc_cse_sva[3727:3720]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1488_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[835:814]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse , (fsm_output[8])});
  assign mul_572_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1487_nl))
      * $signed((ConvFiltWidth_else_mux1h_1488_nl)));
  assign z_out_1153_29_7 = readslicef_30_23_7((mul_572_nl));
  assign ConvFiltWidth_else_mux1h_1489_nl = MUX1HOT_v_8_7_2((w2_rsci_idat_mxwt[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[655:648]), (MultLoop_io_read_w4_rsc_cse_sva[3719:3712]),
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1490_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[967:946]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_17_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_573_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1489_nl))
      * $signed((ConvFiltWidth_else_mux1h_1490_nl)));
  assign z_out_1154_29_7 = readslicef_30_23_7((mul_573_nl));
  assign ConvFiltWidth_else_mux1h_1491_nl = MUX1HOT_v_8_8_2((w2_rsci_idat_mxwt[615:608]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1207:1200]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[7:0]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]),
      (MultLoop_io_read_w4_rsc_cse_sva[5863:5856]), {(fsm_output[1]) , (fsm_output[2])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1492_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[813:792]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_93_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_847_cse , (fsm_output[7]) , (fsm_output[8])});
  assign mul_574_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1491_nl))
      * $signed((ConvFiltWidth_else_mux1h_1492_nl)));
  assign z_out_1155_29_7 = readslicef_30_23_7((mul_574_nl));
  assign ConvFiltWidth_else_mux1h_1493_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[335:328]),
      (w2_rsci_idat_mxwt[1119:1112]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[847:840]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[87:80]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1535:1528]),
      (MultLoop_io_read_w4_rsc_cse_sva[7783:7776]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1494_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_77_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_575_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1493_nl))
      * $signed((ConvFiltWidth_else_mux1h_1494_nl)));
  assign z_out_1156_29_7 = readslicef_30_23_7((mul_575_nl));
  assign ConvFiltWidth_else_mux1h_1495_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[583:576]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[31:24]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[39:32]), (MultLoop_io_read_w4_rsc_cse_sva[7807:7800]),
      {(fsm_output[4]) , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_70_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_576_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1495_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_70_nl)));
  assign z_out_1157_29_7 = readslicef_30_23_7((mul_576_nl));
  assign ConvFiltWidth_else_mux1h_1496_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]),
      (w2_rsci_idat_mxwt[951:944]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[607:600]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]), (MultLoop_io_read_w4_rsc_cse_sva[7799:7792]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1497_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[351:330]),
      (input_1_rsci_idat_mxwt[923:902]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[703:682]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_79_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_17_cse , (fsm_output[1]) , (fsm_output[7]) , (fsm_output[8])});
  assign mul_577_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1496_nl))
      * $signed((ConvFiltWidth_else_mux1h_1497_nl)));
  assign z_out_1158_29_7 = readslicef_30_23_7((mul_577_nl));
  assign ConvFiltWidth_else_mux1h_1498_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[343:336]),
      (w2_rsci_idat_mxwt[1127:1120]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1063:1056]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[279:272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[79:72]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1503:1496]),
      (MultLoop_io_read_w4_rsc_cse_sva[5847:5840]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1499_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[329:308]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , (MultLoop_1124_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_578_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1498_nl))
      * $signed((ConvFiltWidth_else_mux1h_1499_nl)));
  assign z_out_1159_29_7 = readslicef_30_23_7((mul_578_nl));
  assign ConvFiltWidth_else_mux1h_1500_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1583:1576]), (w2_rsci_idat_mxwt[31:24]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1591:1584]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[439:432]), (MultLoop_io_read_w4_rsc_cse_sva[7167:7160]),
      {MultLoop_or_93_cse , (fsm_output[3]) , (fsm_output[1]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1501_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), (input_1_rsci_idat_mxwt[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_579_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1500_nl))
      * $signed((ConvFiltWidth_else_mux1h_1501_nl)));
  assign z_out_1160_29_7 = readslicef_30_23_7((mul_579_nl));
  assign ConvFiltWidth_else_mux1h_1502_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1007:1000]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1543:1536]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1599:1592]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[775:768]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[431:424]),
      (MultLoop_io_read_w4_rsc_cse_sva[8191:8184]), {MultLoop_or_93_cse , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1503_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , ConvFiltWidth_else_or_861_cse , (fsm_output[8])});
  assign mul_580_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1502_nl))
      * $signed((ConvFiltWidth_else_mux1h_1503_nl)));
  assign z_out_1161_29_7 = readslicef_30_23_7((mul_580_nl));
  assign ConvFiltWidth_else_mux1h_1504_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1575:1568]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1383:1376]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[967:960]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[823:816]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[207:200]), (MultLoop_io_read_w4_rsc_cse_sva[9215:9208]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_ConvFiltWidth_else_mux_71_nl = MUX_v_22_2_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_121_if_exu_pmx_20_0_lpi_1_dfm}),
      fsm_output[8]);
  assign mul_581_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1504_nl))
      * $signed((ConvFiltWidth_else_ConvFiltWidth_else_mux_71_nl)));
  assign z_out_1162_29_7 = readslicef_30_23_7((mul_581_nl));
  assign ConvFiltWidth_else_mux1h_1505_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[623:616]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1551:1544]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[815:808]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[215:208]),
      (MultLoop_io_read_w4_rsc_cse_sva[5831:5824]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1506_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , (AccumDotWidth_acc_1937_itm[20:0])}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse
      , (fsm_output[8])});
  assign mul_582_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1505_nl))
      * $signed((ConvFiltWidth_else_mux1h_1506_nl)));
  assign z_out_1163_29_7 = readslicef_30_23_7((mul_582_nl));
  assign ConvFiltWidth_else_mux1h_1507_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[999:992]),
      (w2_rsci_idat_mxwt[223:216]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1271:1264]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1351:1344]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[783:776]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[255:248]), (MultLoop_io_read_w4_rsc_cse_sva[5815:5808]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1508_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , (AccumDotWidth_acc_1916_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_583_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1507_nl))
      * $signed((ConvFiltWidth_else_mux1h_1508_nl)));
  assign z_out_1164_29_7 = readslicef_30_23_7((mul_583_nl));
  assign ConvFiltWidth_else_mux1h_1509_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (w2_rsci_idat_mxwt[239:232]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (MultLoop_io_read_w4_rsc_cse_sva[5823:5816]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1510_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      ({1'b0 , (AccumDotWidth_acc_1932_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , (fsm_output[8])});
  assign mul_584_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1509_nl))
      * $signed((ConvFiltWidth_else_mux1h_1510_nl)));
  assign z_out_1165_29_7 = readslicef_30_23_7((mul_584_nl));
  assign ConvFiltWidth_else_mux1h_1511_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]),
      (w2_rsci_idat_mxwt[607:600]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1567:1560]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1391:1384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[415:408]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[423:416]), (MultLoop_io_read_w4_rsc_cse_sva[5807:5800]),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1512_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]),
      ({1'b0 , (AccumDotWidth_acc_1877_itm[20:0])}), {(fsm_output[2]) , (fsm_output[1])
      , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse , (fsm_output[8])});
  assign mul_585_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1511_nl))
      * $signed((ConvFiltWidth_else_mux1h_1512_nl)));
  assign z_out_1166_29_7 = readslicef_30_23_7((mul_585_nl));
  assign ConvFiltWidth_else_mux1h_1513_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]),
      (w2_rsci_idat_mxwt[47:40]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1359:1352]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[991:984]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[791:784]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[247:240]),
      (MultLoop_io_read_w4_rsc_cse_sva[5839:5832]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1514_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , (AccumDotWidth_acc_1945_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_586_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1513_nl))
      * $signed((ConvFiltWidth_else_mux1h_1514_nl)));
  assign z_out_1167_29_7 = readslicef_30_23_7((mul_586_nl));
  assign ConvFiltWidth_else_mux1h_1515_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[975:968]),
      (w2_rsci_idat_mxwt[215:208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1375:1368]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[799:792]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[231:224]), (MultLoop_io_read_w4_rsc_cse_sva[5855:5848]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1516_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , (MultLoop_1131_nnet_product_layer3_t_config4_weight_t_config4_accum_t_slc_28_7_itm[20:0])}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_587_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1515_nl))
      * $signed((ConvFiltWidth_else_mux1h_1516_nl)));
  assign z_out_1168_29_7 = readslicef_30_23_7((mul_587_nl));
  assign ConvFiltWidth_else_mux1h_1517_nl = MUX1HOT_v_8_8_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[911:904]),
      (w2_rsci_idat_mxwt[1111:1104]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1039:1032]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[687:680]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[263:256]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1511:1504]),
      (MultLoop_io_read_w4_rsc_cse_sva[1511:1504]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1518_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[593:572]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[1055:1034]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_61_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign mul_588_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1517_nl))
      * $signed((ConvFiltWidth_else_mux1h_1518_nl)));
  assign z_out_1169_29_7 = readslicef_30_23_7((mul_588_nl));
  assign ConvFiltWidth_else_mux1h_1519_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]),
      (w2_rsci_idat_mxwt[615:608]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[391:384]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[199:192]),
      (MultLoop_io_read_w4_rsc_cse_sva[7791:7784]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1520_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[945:924]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_78_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_93_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_589_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1519_nl))
      * $signed((ConvFiltWidth_else_mux1h_1520_nl)));
  assign z_out_1170_29_7 = readslicef_30_23_7((mul_589_nl));
  assign ConvFiltWidth_else_mux1h_1521_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[983:976]),
      (w2_rsci_idat_mxwt[231:224]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1367:1360]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[407:400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[239:232]), (MultLoop_io_read_w4_rsc_cse_sva[1559:1552]),
      {MultLoop_or_93_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) ,
      (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1522_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[747:726]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[307:286]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , (fsm_output[3]) , ConvFiltWidth_else_or_787_cse
      , (fsm_output[8])});
  assign mul_590_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1521_nl))
      * $signed((ConvFiltWidth_else_mux1h_1522_nl)));
  assign z_out_1171_29_7 = readslicef_30_23_7((mul_590_nl));
  assign ConvFiltWidth_else_mux1h_1523_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[39:32]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1559:1552]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1399:1392]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[807:800]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[223:216]),
      (MultLoop_io_read_w4_rsc_cse_sva[7775:7768]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1524_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[681:660]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_76_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_55_cse
      , (fsm_output[8])});
  assign mul_591_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1523_nl))
      * $signed((ConvFiltWidth_else_mux1h_1524_nl)));
  assign z_out_1172_29_7 = readslicef_30_23_7((mul_591_nl));
  assign ConvFiltWidth_else_mux1h_1525_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1023:1016]),
      (w2_rsci_idat_mxwt[23:16]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1407:1400]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[399:392]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[447:440]),
      (MultLoop_io_read_w4_rsc_cse_sva[7703:7696]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1526_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[615:594]),
      (input_1_rsci_idat_mxwt[681:660]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[483:462]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_67_if_exu_pmx_20_0_lpi_1_dfm}),
      {MultLoop_or_93_cse , (fsm_output[1]) , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_592_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1525_nl))
      * $signed((ConvFiltWidth_else_mux1h_1526_nl)));
  assign z_out_1173_29_7 = readslicef_30_23_7((mul_592_nl));
  assign ConvFiltWidth_else_mux1h_1527_nl = MUX1HOT_v_8_7_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (w2_rsci_idat_mxwt[1151:1144]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1015:1008]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[831:824]), (MultLoop_io_read_w4_rsc_cse_sva[6903:6896]),
      {(fsm_output[3]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6])
      , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1528_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]),
      (input_1_rsci_idat_mxwt[1055:1034]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[681:660]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_95_if_exu_pmx_20_0_lpi_1_dfm}),
      {nnet_product_layer3_t_config4_weight_t_config4_accum_t_or_4_cse , (fsm_output[1])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_593_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1527_nl))
      * $signed((ConvFiltWidth_else_mux1h_1528_nl)));
  assign z_out_1174_29_7 = readslicef_30_23_7((mul_593_nl));
  assign ConvFiltWidth_else_mux1h_1529_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[471:464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1655:1648]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1663:1656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]), (MultLoop_io_read_w4_rsc_cse_sva[1671:1664]),
      {(fsm_output[1]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1530_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[769:748]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_142_cse , (fsm_output[8])});
  assign mul_594_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1529_nl))
      * $signed((ConvFiltWidth_else_mux1h_1530_nl)));
  assign z_out_1175_29_7 = readslicef_30_23_7((mul_594_nl));
  assign ConvFiltWidth_else_mux1h_1531_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[279:272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (MultLoop_io_read_w4_rsc_cse_sva[1663:1656]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1532_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[703:682]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_80_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , AccumDotWidth_or_139_cse , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_595_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1531_nl))
      * $signed((ConvFiltWidth_else_mux1h_1532_nl)));
  assign z_out_1176_29_7 = readslicef_30_23_7((mul_595_nl));
  assign ConvFiltWidth_else_mux1h_1533_nl = MUX1HOT_v_8_5_2((w2_rsci_idat_mxwt[87:80]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1639:1632]), (MultLoop_io_read_w4_rsc_cse_sva[1527:1520]),
      {(fsm_output[1]) , AccumDotWidth_or_157_cse , (fsm_output[4]) , (fsm_output[5])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1534_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[637:616]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_63_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_152_cse , (fsm_output[8])});
  assign mul_596_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1533_nl))
      * $signed((ConvFiltWidth_else_mux1h_1534_nl)));
  assign z_out_1177_29_7 = readslicef_30_23_7((mul_596_nl));
  assign ConvFiltWidth_else_mux1h_1535_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[671:664]),
      (w2_rsci_idat_mxwt[1055:1048]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[703:696]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1647:1640]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]),
      (MultLoop_io_read_w4_rsc_cse_sva[1679:1672]), {AccumDotWidth_or_25_cse , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1536_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[1033:1012]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_82_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_46_cse , AccumDotWidth_or_152_cse
      , (fsm_output[8])});
  assign mul_597_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1535_nl))
      * $signed((ConvFiltWidth_else_mux1h_1536_nl)));
  assign z_out_1178_29_7 = readslicef_30_23_7((mul_597_nl));
  assign ConvFiltWidth_else_mux1h_1537_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (w2_rsci_idat_mxwt[215:208]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1223:1216]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1255:1248]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[311:304]),
      (MultLoop_io_read_w4_rsc_cse_sva[1687:1680]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1538_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[681:660]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_83_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_598_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1537_nl))
      * $signed((ConvFiltWidth_else_mux1h_1538_nl)));
  assign z_out_1179_29_7 = readslicef_30_23_7((mul_598_nl));
  assign ConvFiltWidth_else_mux1h_1539_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[663:656]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1415:1408]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1279:1272]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[695:688]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[271:264]),
      (MultLoop_io_read_w4_rsc_cse_sva[1695:1688]), {AccumDotWidth_or_25_cse , (fsm_output[4])
      , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1540_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_84_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_882_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_599_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1539_nl))
      * $signed((ConvFiltWidth_else_mux1h_1540_nl)));
  assign z_out_1180_29_7 = readslicef_30_23_7((mul_599_nl));
  assign ConvFiltWidth_else_mux1h_1541_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]),
      (w2_rsci_idat_mxwt[159:152]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1463:1456]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[895:888]), (MultLoop_io_read_w4_rsc_cse_sva[1551:1544]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , AccumDotWidth_or_145_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1542_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[659:638]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_600_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1541_nl))
      * $signed((ConvFiltWidth_else_mux1h_1542_nl)));
  assign z_out_1181_29_7 = readslicef_30_23_7((mul_600_nl));
  assign ConvFiltWidth_else_mux1h_1543_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (w2_rsci_idat_mxwt[599:592]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1447:1440]), (MultLoop_io_read_w4_rsc_cse_sva[1519:1512]),
      {(fsm_output[2]) , (fsm_output[1]) , MultLoop_or_22_cse , AccumDotWidth_or_145_cse
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1544_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[879:858]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_601_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1543_nl))
      * $signed((ConvFiltWidth_else_mux1h_1544_nl)));
  assign z_out_1182_29_7 = readslicef_30_23_7((mul_601_nl));
  assign ConvFiltWidth_else_mux1h_1545_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[871:864]),
      (w2_rsci_idat_mxwt[407:400]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1231:1224]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1263:1256]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[71:64]),
      (MultLoop_io_read_w4_rsc_cse_sva[1535:1528]), {(fsm_output[2]) , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1546_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[747:726]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_64_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[1]) , (fsm_output[8])});
  assign mul_602_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1545_nl))
      * $signed((ConvFiltWidth_else_mux1h_1546_nl)));
  assign z_out_1183_29_7 = readslicef_30_23_7((mul_602_nl));
  assign ConvFiltWidth_else_mux1h_1547_nl = MUX1HOT_v_8_6_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[879:872]),
      (w2_rsci_idat_mxwt[23:16]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1471:1464]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1247:1240]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[319:312]),
      (MultLoop_io_read_w4_rsc_cse_sva[7695:7688]), {AccumDotWidth_or_25_cse , (fsm_output[1])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1548_nl = MUX1HOT_v_22_4_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[615:594]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_66_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[1]) , (fsm_output[3]) , (fsm_output[8])});
  assign mul_603_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1547_nl))
      * $signed((ConvFiltWidth_else_mux1h_1548_nl)));
  assign z_out_1184_29_7 = readslicef_30_23_7((mul_603_nl));
  assign ConvFiltWidth_else_mux1h_1549_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[647:640]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1439:1432]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1239:1232]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[303:296]), (MultLoop_io_read_w4_rsc_cse_sva[7815:7808]),
      {AccumDotWidth_or_25_cse , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1550_nl = MUX1HOT_v_22_3_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_81_if_exu_pmx_20_0_lpi_1_dfm}),
      {ConvFiltWidth_else_or_1081_cse , (fsm_output[3]) , (fsm_output[8])});
  assign mul_604_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1549_nl))
      * $signed((ConvFiltWidth_else_mux1h_1550_nl)));
  assign z_out_1185_29_7 = readslicef_30_23_7((mul_604_nl));
  assign ConvFiltWidth_else_mux1h_1551_nl = MUX1HOT_v_8_5_2((ConvFiltWidth_else_io_read_w2_rsc_cse_sva[855:848]),
      (w2_rsci_idat_mxwt[983:976]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1455:1448]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[863:856]), (MultLoop_io_read_w4_rsc_cse_sva[6911:6904]),
      {AccumDotWidth_or_25_cse , (fsm_output[1]) , AccumDotWidth_or_145_cse , (fsm_output[7])
      , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1552_nl = MUX1HOT_v_22_5_2((ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]),
      (input_1_rsci_idat_mxwt[1011:990]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_96_if_exu_pmx_20_0_lpi_1_dfm}),
      {operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[1]) , (fsm_output[3])
      , AccumDotWidth_or_140_cse , (fsm_output[8])});
  assign mul_605_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1551_nl))
      * $signed((ConvFiltWidth_else_mux1h_1552_nl)));
  assign z_out_1186_29_7 = readslicef_30_23_7((mul_605_nl));
  assign ConvFiltWidth_else_mux1h_1553_nl = MUX1HOT_v_8_6_2((w2_rsci_idat_mxwt[759:752]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1087:1080]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[679:672]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[487:480]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[95:88]),
      (MultLoop_io_read_w4_rsc_cse_sva[7663:7656]), {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[5]) , (fsm_output[6]) , (fsm_output[8])});
  assign ConvFiltWidth_else_mux1h_1554_nl = MUX1HOT_v_22_3_2((input_1_rsci_idat_mxwt[923:902]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[175:154]), ({1'b0 , nnet_relu_layer2_t_layer3_t_relu_config3_for_62_if_exu_pmx_20_0_lpi_1_dfm}),
      {(fsm_output[1]) , ConvFiltWidth_else_or_730_cse , (fsm_output[8])});
  assign mul_606_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1553_nl))
      * $signed((ConvFiltWidth_else_mux1h_1554_nl)));
  assign z_out_1187_29_7 = readslicef_30_23_7((mul_606_nl));
  assign ConvFiltWidth_else_mux1h_1555_nl = MUX1HOT_v_8_4_2((w2_rsci_idat_mxwt[791:784]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[287:280]), (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[887:880]),
      (ConvFiltWidth_else_io_read_w2_rsc_cse_sva[1431:1424]), {(fsm_output[1]) ,
      (fsm_output[2]) , MultLoop_or_22_cse , AccumDotWidth_or_145_cse});
  assign ConvFiltWidth_else_mux1h_1556_nl = MUX1HOT_v_22_4_2((input_1_rsci_idat_mxwt[945:924]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[571:550]), (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[109:88]),
      (ConvFiltWidth_else_io_read_input_1_rsc_cse_sva[769:748]), {(fsm_output[1])
      , operator_22_4_true_AC_TRN_AC_WRAP_or_7_cse , (fsm_output[3]) , AccumDotWidth_or_140_cse});
  assign mul_607_nl = conv_u2u_30_30($signed((ConvFiltWidth_else_mux1h_1555_nl))
      * $signed((ConvFiltWidth_else_mux1h_1556_nl)));
  assign z_out_1188_29_9 = readslicef_30_21_9((mul_607_nl));

  function automatic [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_6_2;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [5:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    MUX1HOT_v_10_6_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_7_2;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [6:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    MUX1HOT_v_10_7_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_4_2;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [3:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    MUX1HOT_v_11_4_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_5_2;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [4:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    MUX1HOT_v_11_5_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_6_2;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [5:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    result = result | ( input_5 & {11{sel[5]}});
    MUX1HOT_v_11_6_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_7_2;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [6:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    result = result | ( input_5 & {11{sel[5]}});
    result = result | ( input_6 & {11{sel[6]}});
    MUX1HOT_v_11_7_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_8_2;
    input [10:0] input_7;
    input [10:0] input_6;
    input [10:0] input_5;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [7:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | ( input_1 & {11{sel[1]}});
    result = result | ( input_2 & {11{sel[2]}});
    result = result | ( input_3 & {11{sel[3]}});
    result = result | ( input_4 & {11{sel[4]}});
    result = result | ( input_5 & {11{sel[5]}});
    result = result | ( input_6 & {11{sel[6]}});
    result = result | ( input_7 & {11{sel[7]}});
    MUX1HOT_v_11_8_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_3_2;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [2:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | ( input_1 & {21{sel[1]}});
    result = result | ( input_2 & {21{sel[2]}});
    MUX1HOT_v_21_3_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_4_2;
    input [20:0] input_3;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [3:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | ( input_1 & {21{sel[1]}});
    result = result | ( input_2 & {21{sel[2]}});
    result = result | ( input_3 & {21{sel[3]}});
    MUX1HOT_v_21_4_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_5_2;
    input [20:0] input_4;
    input [20:0] input_3;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [4:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | ( input_1 & {21{sel[1]}});
    result = result | ( input_2 & {21{sel[2]}});
    result = result | ( input_3 & {21{sel[3]}});
    result = result | ( input_4 & {21{sel[4]}});
    MUX1HOT_v_21_5_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_6_2;
    input [20:0] input_5;
    input [20:0] input_4;
    input [20:0] input_3;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [5:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | ( input_1 & {21{sel[1]}});
    result = result | ( input_2 & {21{sel[2]}});
    result = result | ( input_3 & {21{sel[3]}});
    result = result | ( input_4 & {21{sel[4]}});
    result = result | ( input_5 & {21{sel[5]}});
    MUX1HOT_v_21_6_2 = result;
  end
  endfunction


  function automatic [20:0] MUX1HOT_v_21_7_2;
    input [20:0] input_6;
    input [20:0] input_5;
    input [20:0] input_4;
    input [20:0] input_3;
    input [20:0] input_2;
    input [20:0] input_1;
    input [20:0] input_0;
    input [6:0] sel;
    reg [20:0] result;
  begin
    result = input_0 & {21{sel[0]}};
    result = result | ( input_1 & {21{sel[1]}});
    result = result | ( input_2 & {21{sel[2]}});
    result = result | ( input_3 & {21{sel[3]}});
    result = result | ( input_4 & {21{sel[4]}});
    result = result | ( input_5 & {21{sel[5]}});
    result = result | ( input_6 & {21{sel[6]}});
    MUX1HOT_v_21_7_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_3_2;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [2:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    MUX1HOT_v_22_3_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_4_2;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [3:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    MUX1HOT_v_22_4_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_5_2;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [4:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    result = result | ( input_4 & {22{sel[4]}});
    MUX1HOT_v_22_5_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_6_2;
    input [21:0] input_5;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [5:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    result = result | ( input_4 & {22{sel[4]}});
    result = result | ( input_5 & {22{sel[5]}});
    MUX1HOT_v_22_6_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_7_2;
    input [21:0] input_6;
    input [21:0] input_5;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [6:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    result = result | ( input_4 & {22{sel[4]}});
    result = result | ( input_5 & {22{sel[5]}});
    result = result | ( input_6 & {22{sel[6]}});
    MUX1HOT_v_22_7_2 = result;
  end
  endfunction


  function automatic [21:0] MUX1HOT_v_22_8_2;
    input [21:0] input_7;
    input [21:0] input_6;
    input [21:0] input_5;
    input [21:0] input_4;
    input [21:0] input_3;
    input [21:0] input_2;
    input [21:0] input_1;
    input [21:0] input_0;
    input [7:0] sel;
    reg [21:0] result;
  begin
    result = input_0 & {22{sel[0]}};
    result = result | ( input_1 & {22{sel[1]}});
    result = result | ( input_2 & {22{sel[2]}});
    result = result | ( input_3 & {22{sel[3]}});
    result = result | ( input_4 & {22{sel[4]}});
    result = result | ( input_5 & {22{sel[5]}});
    result = result | ( input_6 & {22{sel[6]}});
    result = result | ( input_7 & {22{sel[7]}});
    MUX1HOT_v_22_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_7_2;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [6:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    MUX1HOT_v_8_7_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_8_2;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [7:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    MUX1HOT_v_8_8_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_23_1_22;
    input [22:0] vector;
    reg [22:0] tmp;
  begin
    tmp = vector >> 22;
    readslicef_23_1_22 = tmp[0:0];
  end
  endfunction


  function automatic [21:0] readslicef_29_22_7;
    input [28:0] vector;
    reg [28:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_29_22_7 = tmp[21:0];
  end
  endfunction


  function automatic [20:0] readslicef_30_21_9;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_30_21_9 = tmp[20:0];
  end
  endfunction


  function automatic [22:0] readslicef_30_23_7;
    input [29:0] vector;
    reg [29:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_30_23_7 = tmp[22:0];
  end
  endfunction


  function automatic [10:0] signext_11_10;
    input [9:0] vector;
  begin
    signext_11_10= {{1{vector[9]}}, vector};
  end
  endfunction


  function automatic [21:0] signext_22_21;
    input [20:0] vector;
  begin
    signext_22_21= {{1{vector[20]}}, vector};
  end
  endfunction


  function automatic [9:0] conv_s2s_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2s_8_11 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_11 = {{3{vector[7]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2s_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2s_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2s_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [9:0] conv_s2u_8_10 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_10 = {{2{vector[7]}}, vector};
  end
  endfunction


  function automatic [10:0] conv_s2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_s2u_8_11 = {{3{vector[7]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_22_23 ;
    input [21:0]  vector ;
  begin
    conv_s2u_22_23 = {vector[21], vector};
  end
  endfunction


  function automatic [21:0] conv_u2s_21_22 ;
    input [20:0]  vector ;
  begin
    conv_u2s_21_22 =  {1'b0, vector};
  end
  endfunction


  function automatic [29:0] conv_u2u_30_30 ;
    input [29:0]  vector ;
  begin
    conv_u2u_30_30 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    econ_4x4_d10
// ------------------------------------------------------------------


module econ_4x4_d10 (
  clk, rst, input_1_rsc_dat, input_1_rsc_vld, input_1_rsc_triosy_lz, layer5_out_rsc_dat,
      layer5_out_rsc_vld, layer5_out_rsc_triosy_lz, const_size_in_1_rsc_dat, const_size_in_1_rsc_vld,
      const_size_in_1_rsc_triosy_lz, const_size_out_1_rsc_dat, const_size_out_1_rsc_vld,
      const_size_out_1_rsc_triosy_lz, w2_rsc_dat, w2_rsc_vld, w2_rsc_triosy_lz, b2_rsc_dat,
      b2_rsc_vld, b2_rsc_triosy_lz, w4_rsc_dat, w4_rsc_vld, w4_rsc_triosy_lz, b4_rsc_dat,
      b4_rsc_vld, b4_rsc_triosy_lz
);
  input clk;
  input rst;
  input [1055:0] input_1_rsc_dat;
  input input_1_rsc_vld;
  output input_1_rsc_triosy_lz;
  output [219:0] layer5_out_rsc_dat;
  output layer5_out_rsc_vld;
  output layer5_out_rsc_triosy_lz;
  output [15:0] const_size_in_1_rsc_dat;
  output const_size_in_1_rsc_vld;
  output const_size_in_1_rsc_triosy_lz;
  output [15:0] const_size_out_1_rsc_dat;
  output const_size_out_1_rsc_vld;
  output const_size_out_1_rsc_triosy_lz;
  input [1727:0] w2_rsc_dat;
  input w2_rsc_vld;
  output w2_rsc_triosy_lz;
  input [63:0] b2_rsc_dat;
  input b2_rsc_vld;
  output b2_rsc_triosy_lz;
  input [10239:0] w4_rsc_dat;
  input w4_rsc_vld;
  output w4_rsc_triosy_lz;
  input [79:0] b4_rsc_dat;
  input b4_rsc_vld;
  output b4_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  econ_4x4_d10_core econ_4x4_d10_core_inst (
      .clk(clk),
      .rst(rst),
      .input_1_rsc_dat(input_1_rsc_dat),
      .input_1_rsc_vld(input_1_rsc_vld),
      .input_1_rsc_triosy_lz(input_1_rsc_triosy_lz),
      .layer5_out_rsc_dat(layer5_out_rsc_dat),
      .layer5_out_rsc_vld(layer5_out_rsc_vld),
      .layer5_out_rsc_triosy_lz(layer5_out_rsc_triosy_lz),
      .const_size_in_1_rsc_dat(const_size_in_1_rsc_dat),
      .const_size_in_1_rsc_vld(const_size_in_1_rsc_vld),
      .const_size_in_1_rsc_triosy_lz(const_size_in_1_rsc_triosy_lz),
      .const_size_out_1_rsc_dat(const_size_out_1_rsc_dat),
      .const_size_out_1_rsc_vld(const_size_out_1_rsc_vld),
      .const_size_out_1_rsc_triosy_lz(const_size_out_1_rsc_triosy_lz),
      .w2_rsc_dat(w2_rsc_dat),
      .w2_rsc_vld(w2_rsc_vld),
      .w2_rsc_triosy_lz(w2_rsc_triosy_lz),
      .b2_rsc_dat(b2_rsc_dat),
      .b2_rsc_vld(b2_rsc_vld),
      .b2_rsc_triosy_lz(b2_rsc_triosy_lz),
      .w4_rsc_dat(w4_rsc_dat),
      .w4_rsc_vld(w4_rsc_vld),
      .w4_rsc_triosy_lz(w4_rsc_triosy_lz),
      .b4_rsc_dat(b4_rsc_dat),
      .b4_rsc_vld(b4_rsc_vld),
      .b4_rsc_triosy_lz(b4_rsc_triosy_lz)
    );
endmodule



